// This is the unpowered netlist.
module ExperiarCore (clk0,
    clk1,
    core_wb_ack_i,
    core_wb_cyc_o,
    core_wb_error_i,
    core_wb_stall_i,
    core_wb_stb_o,
    core_wb_we_o,
    jtag_tck,
    jtag_tdi,
    jtag_tdo,
    jtag_tms,
    localMemory_wb_ack_o,
    localMemory_wb_cyc_i,
    localMemory_wb_error_o,
    localMemory_wb_stall_o,
    localMemory_wb_stb_i,
    localMemory_wb_we_i,
    probe_state,
    wb_clk_i,
    wb_rst_i,
    web0,
    addr0,
    addr1,
    coreIndex,
    core_wb_adr_o,
    core_wb_data_i,
    core_wb_data_o,
    core_wb_sel_o,
    csb0,
    csb1,
    din0,
    dout0,
    dout1,
    irq,
    localMemory_wb_adr_i,
    localMemory_wb_data_i,
    localMemory_wb_data_o,
    localMemory_wb_sel_i,
    manufacturerID,
    partID,
    probe_env,
    probe_jtagInstruction,
    probe_programCounter,
    versionID,
    wmask0);
 output clk0;
 output clk1;
 input core_wb_ack_i;
 output core_wb_cyc_o;
 input core_wb_error_i;
 input core_wb_stall_i;
 output core_wb_stb_o;
 output core_wb_we_o;
 input jtag_tck;
 input jtag_tdi;
 output jtag_tdo;
 input jtag_tms;
 output localMemory_wb_ack_o;
 input localMemory_wb_cyc_i;
 output localMemory_wb_error_o;
 output localMemory_wb_stall_o;
 input localMemory_wb_stb_i;
 input localMemory_wb_we_i;
 output probe_state;
 input wb_clk_i;
 input wb_rst_i;
 output web0;
 output [8:0] addr0;
 output [8:0] addr1;
 input [7:0] coreIndex;
 output [27:0] core_wb_adr_o;
 input [31:0] core_wb_data_i;
 output [31:0] core_wb_data_o;
 output [3:0] core_wb_sel_o;
 output [1:0] csb0;
 output [1:0] csb1;
 output [31:0] din0;
 input [63:0] dout0;
 input [63:0] dout1;
 input [15:0] irq;
 input [23:0] localMemory_wb_adr_i;
 input [31:0] localMemory_wb_data_i;
 output [31:0] localMemory_wb_data_o;
 input [3:0] localMemory_wb_sel_i;
 input [10:0] manufacturerID;
 input [15:0] partID;
 output [1:0] probe_env;
 output [4:0] probe_jtagInstruction;
 output [31:0] probe_programCounter;
 input [3:0] versionID;
 output [3:0] wmask0;

 wire net2007;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_131_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_133_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_140_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_144_wb_clk_i;
 wire clknet_leaf_145_wb_clk_i;
 wire clknet_leaf_146_wb_clk_i;
 wire clknet_leaf_147_wb_clk_i;
 wire clknet_leaf_148_wb_clk_i;
 wire clknet_leaf_149_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_150_wb_clk_i;
 wire clknet_leaf_151_wb_clk_i;
 wire clknet_leaf_152_wb_clk_i;
 wire clknet_leaf_153_wb_clk_i;
 wire clknet_leaf_154_wb_clk_i;
 wire clknet_leaf_155_wb_clk_i;
 wire clknet_leaf_156_wb_clk_i;
 wire clknet_leaf_157_wb_clk_i;
 wire clknet_leaf_158_wb_clk_i;
 wire clknet_leaf_159_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_160_wb_clk_i;
 wire clknet_leaf_161_wb_clk_i;
 wire clknet_leaf_162_wb_clk_i;
 wire clknet_leaf_163_wb_clk_i;
 wire clknet_leaf_164_wb_clk_i;
 wire clknet_leaf_165_wb_clk_i;
 wire clknet_leaf_166_wb_clk_i;
 wire clknet_leaf_167_wb_clk_i;
 wire clknet_leaf_168_wb_clk_i;
 wire clknet_leaf_169_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_170_wb_clk_i;
 wire clknet_leaf_171_wb_clk_i;
 wire clknet_leaf_172_wb_clk_i;
 wire clknet_leaf_173_wb_clk_i;
 wire clknet_leaf_174_wb_clk_i;
 wire clknet_leaf_175_wb_clk_i;
 wire clknet_leaf_176_wb_clk_i;
 wire clknet_leaf_177_wb_clk_i;
 wire clknet_leaf_178_wb_clk_i;
 wire clknet_leaf_179_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_180_wb_clk_i;
 wire clknet_leaf_181_wb_clk_i;
 wire clknet_leaf_182_wb_clk_i;
 wire clknet_leaf_183_wb_clk_i;
 wire clknet_leaf_184_wb_clk_i;
 wire clknet_leaf_185_wb_clk_i;
 wire clknet_leaf_186_wb_clk_i;
 wire clknet_leaf_188_wb_clk_i;
 wire clknet_leaf_189_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_190_wb_clk_i;
 wire clknet_leaf_191_wb_clk_i;
 wire clknet_leaf_192_wb_clk_i;
 wire clknet_leaf_193_wb_clk_i;
 wire clknet_leaf_194_wb_clk_i;
 wire clknet_leaf_195_wb_clk_i;
 wire clknet_leaf_196_wb_clk_i;
 wire clknet_leaf_197_wb_clk_i;
 wire clknet_leaf_198_wb_clk_i;
 wire clknet_leaf_199_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_200_wb_clk_i;
 wire clknet_leaf_201_wb_clk_i;
 wire clknet_leaf_202_wb_clk_i;
 wire clknet_leaf_203_wb_clk_i;
 wire clknet_leaf_204_wb_clk_i;
 wire clknet_leaf_205_wb_clk_i;
 wire clknet_leaf_206_wb_clk_i;
 wire clknet_leaf_207_wb_clk_i;
 wire clknet_leaf_208_wb_clk_i;
 wire clknet_leaf_209_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_210_wb_clk_i;
 wire clknet_leaf_211_wb_clk_i;
 wire clknet_leaf_212_wb_clk_i;
 wire clknet_leaf_213_wb_clk_i;
 wire clknet_leaf_214_wb_clk_i;
 wire clknet_leaf_215_wb_clk_i;
 wire clknet_leaf_216_wb_clk_i;
 wire clknet_leaf_217_wb_clk_i;
 wire clknet_leaf_218_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \core.cancelStall ;
 wire \core.csr.currentInstruction[0] ;
 wire \core.csr.currentInstruction[10] ;
 wire \core.csr.currentInstruction[11] ;
 wire \core.csr.currentInstruction[12] ;
 wire \core.csr.currentInstruction[13] ;
 wire \core.csr.currentInstruction[14] ;
 wire \core.csr.currentInstruction[15] ;
 wire \core.csr.currentInstruction[16] ;
 wire \core.csr.currentInstruction[17] ;
 wire \core.csr.currentInstruction[18] ;
 wire \core.csr.currentInstruction[19] ;
 wire \core.csr.currentInstruction[1] ;
 wire \core.csr.currentInstruction[20] ;
 wire \core.csr.currentInstruction[21] ;
 wire \core.csr.currentInstruction[22] ;
 wire \core.csr.currentInstruction[23] ;
 wire \core.csr.currentInstruction[24] ;
 wire \core.csr.currentInstruction[25] ;
 wire \core.csr.currentInstruction[26] ;
 wire \core.csr.currentInstruction[27] ;
 wire \core.csr.currentInstruction[28] ;
 wire \core.csr.currentInstruction[29] ;
 wire \core.csr.currentInstruction[2] ;
 wire \core.csr.currentInstruction[30] ;
 wire \core.csr.currentInstruction[31] ;
 wire \core.csr.currentInstruction[3] ;
 wire \core.csr.currentInstruction[4] ;
 wire \core.csr.currentInstruction[5] ;
 wire \core.csr.currentInstruction[6] ;
 wire \core.csr.currentInstruction[7] ;
 wire \core.csr.currentInstruction[8] ;
 wire \core.csr.currentInstruction[9] ;
 wire \core.csr.cycleTimer.currentValue[0] ;
 wire \core.csr.cycleTimer.currentValue[10] ;
 wire \core.csr.cycleTimer.currentValue[11] ;
 wire \core.csr.cycleTimer.currentValue[12] ;
 wire \core.csr.cycleTimer.currentValue[13] ;
 wire \core.csr.cycleTimer.currentValue[14] ;
 wire \core.csr.cycleTimer.currentValue[15] ;
 wire \core.csr.cycleTimer.currentValue[16] ;
 wire \core.csr.cycleTimer.currentValue[17] ;
 wire \core.csr.cycleTimer.currentValue[18] ;
 wire \core.csr.cycleTimer.currentValue[19] ;
 wire \core.csr.cycleTimer.currentValue[1] ;
 wire \core.csr.cycleTimer.currentValue[20] ;
 wire \core.csr.cycleTimer.currentValue[21] ;
 wire \core.csr.cycleTimer.currentValue[22] ;
 wire \core.csr.cycleTimer.currentValue[23] ;
 wire \core.csr.cycleTimer.currentValue[24] ;
 wire \core.csr.cycleTimer.currentValue[25] ;
 wire \core.csr.cycleTimer.currentValue[26] ;
 wire \core.csr.cycleTimer.currentValue[27] ;
 wire \core.csr.cycleTimer.currentValue[28] ;
 wire \core.csr.cycleTimer.currentValue[29] ;
 wire \core.csr.cycleTimer.currentValue[2] ;
 wire \core.csr.cycleTimer.currentValue[30] ;
 wire \core.csr.cycleTimer.currentValue[31] ;
 wire \core.csr.cycleTimer.currentValue[32] ;
 wire \core.csr.cycleTimer.currentValue[33] ;
 wire \core.csr.cycleTimer.currentValue[34] ;
 wire \core.csr.cycleTimer.currentValue[35] ;
 wire \core.csr.cycleTimer.currentValue[36] ;
 wire \core.csr.cycleTimer.currentValue[37] ;
 wire \core.csr.cycleTimer.currentValue[38] ;
 wire \core.csr.cycleTimer.currentValue[39] ;
 wire \core.csr.cycleTimer.currentValue[3] ;
 wire \core.csr.cycleTimer.currentValue[40] ;
 wire \core.csr.cycleTimer.currentValue[41] ;
 wire \core.csr.cycleTimer.currentValue[42] ;
 wire \core.csr.cycleTimer.currentValue[43] ;
 wire \core.csr.cycleTimer.currentValue[44] ;
 wire \core.csr.cycleTimer.currentValue[45] ;
 wire \core.csr.cycleTimer.currentValue[46] ;
 wire \core.csr.cycleTimer.currentValue[47] ;
 wire \core.csr.cycleTimer.currentValue[48] ;
 wire \core.csr.cycleTimer.currentValue[49] ;
 wire \core.csr.cycleTimer.currentValue[4] ;
 wire \core.csr.cycleTimer.currentValue[50] ;
 wire \core.csr.cycleTimer.currentValue[51] ;
 wire \core.csr.cycleTimer.currentValue[52] ;
 wire \core.csr.cycleTimer.currentValue[53] ;
 wire \core.csr.cycleTimer.currentValue[54] ;
 wire \core.csr.cycleTimer.currentValue[55] ;
 wire \core.csr.cycleTimer.currentValue[56] ;
 wire \core.csr.cycleTimer.currentValue[57] ;
 wire \core.csr.cycleTimer.currentValue[58] ;
 wire \core.csr.cycleTimer.currentValue[59] ;
 wire \core.csr.cycleTimer.currentValue[5] ;
 wire \core.csr.cycleTimer.currentValue[60] ;
 wire \core.csr.cycleTimer.currentValue[61] ;
 wire \core.csr.cycleTimer.currentValue[62] ;
 wire \core.csr.cycleTimer.currentValue[63] ;
 wire \core.csr.cycleTimer.currentValue[6] ;
 wire \core.csr.cycleTimer.currentValue[7] ;
 wire \core.csr.cycleTimer.currentValue[8] ;
 wire \core.csr.cycleTimer.currentValue[9] ;
 wire \core.csr.inTrap ;
 wire \core.csr.instretTimer.currentValue[0] ;
 wire \core.csr.instretTimer.currentValue[10] ;
 wire \core.csr.instretTimer.currentValue[11] ;
 wire \core.csr.instretTimer.currentValue[12] ;
 wire \core.csr.instretTimer.currentValue[13] ;
 wire \core.csr.instretTimer.currentValue[14] ;
 wire \core.csr.instretTimer.currentValue[15] ;
 wire \core.csr.instretTimer.currentValue[16] ;
 wire \core.csr.instretTimer.currentValue[17] ;
 wire \core.csr.instretTimer.currentValue[18] ;
 wire \core.csr.instretTimer.currentValue[19] ;
 wire \core.csr.instretTimer.currentValue[1] ;
 wire \core.csr.instretTimer.currentValue[20] ;
 wire \core.csr.instretTimer.currentValue[21] ;
 wire \core.csr.instretTimer.currentValue[22] ;
 wire \core.csr.instretTimer.currentValue[23] ;
 wire \core.csr.instretTimer.currentValue[24] ;
 wire \core.csr.instretTimer.currentValue[25] ;
 wire \core.csr.instretTimer.currentValue[26] ;
 wire \core.csr.instretTimer.currentValue[27] ;
 wire \core.csr.instretTimer.currentValue[28] ;
 wire \core.csr.instretTimer.currentValue[29] ;
 wire \core.csr.instretTimer.currentValue[2] ;
 wire \core.csr.instretTimer.currentValue[30] ;
 wire \core.csr.instretTimer.currentValue[31] ;
 wire \core.csr.instretTimer.currentValue[32] ;
 wire \core.csr.instretTimer.currentValue[33] ;
 wire \core.csr.instretTimer.currentValue[34] ;
 wire \core.csr.instretTimer.currentValue[35] ;
 wire \core.csr.instretTimer.currentValue[36] ;
 wire \core.csr.instretTimer.currentValue[37] ;
 wire \core.csr.instretTimer.currentValue[38] ;
 wire \core.csr.instretTimer.currentValue[39] ;
 wire \core.csr.instretTimer.currentValue[3] ;
 wire \core.csr.instretTimer.currentValue[40] ;
 wire \core.csr.instretTimer.currentValue[41] ;
 wire \core.csr.instretTimer.currentValue[42] ;
 wire \core.csr.instretTimer.currentValue[43] ;
 wire \core.csr.instretTimer.currentValue[44] ;
 wire \core.csr.instretTimer.currentValue[45] ;
 wire \core.csr.instretTimer.currentValue[46] ;
 wire \core.csr.instretTimer.currentValue[47] ;
 wire \core.csr.instretTimer.currentValue[48] ;
 wire \core.csr.instretTimer.currentValue[49] ;
 wire \core.csr.instretTimer.currentValue[4] ;
 wire \core.csr.instretTimer.currentValue[50] ;
 wire \core.csr.instretTimer.currentValue[51] ;
 wire \core.csr.instretTimer.currentValue[52] ;
 wire \core.csr.instretTimer.currentValue[53] ;
 wire \core.csr.instretTimer.currentValue[54] ;
 wire \core.csr.instretTimer.currentValue[55] ;
 wire \core.csr.instretTimer.currentValue[56] ;
 wire \core.csr.instretTimer.currentValue[57] ;
 wire \core.csr.instretTimer.currentValue[58] ;
 wire \core.csr.instretTimer.currentValue[59] ;
 wire \core.csr.instretTimer.currentValue[5] ;
 wire \core.csr.instretTimer.currentValue[60] ;
 wire \core.csr.instretTimer.currentValue[61] ;
 wire \core.csr.instretTimer.currentValue[62] ;
 wire \core.csr.instretTimer.currentValue[63] ;
 wire \core.csr.instretTimer.currentValue[6] ;
 wire \core.csr.instretTimer.currentValue[7] ;
 wire \core.csr.instretTimer.currentValue[8] ;
 wire \core.csr.instretTimer.currentValue[9] ;
 wire \core.csr.instruction_memoryAddress[0] ;
 wire \core.csr.instruction_memoryAddress[10] ;
 wire \core.csr.instruction_memoryAddress[11] ;
 wire \core.csr.instruction_memoryAddress[12] ;
 wire \core.csr.instruction_memoryAddress[13] ;
 wire \core.csr.instruction_memoryAddress[14] ;
 wire \core.csr.instruction_memoryAddress[15] ;
 wire \core.csr.instruction_memoryAddress[16] ;
 wire \core.csr.instruction_memoryAddress[17] ;
 wire \core.csr.instruction_memoryAddress[18] ;
 wire \core.csr.instruction_memoryAddress[19] ;
 wire \core.csr.instruction_memoryAddress[1] ;
 wire \core.csr.instruction_memoryAddress[20] ;
 wire \core.csr.instruction_memoryAddress[21] ;
 wire \core.csr.instruction_memoryAddress[22] ;
 wire \core.csr.instruction_memoryAddress[23] ;
 wire \core.csr.instruction_memoryAddress[24] ;
 wire \core.csr.instruction_memoryAddress[25] ;
 wire \core.csr.instruction_memoryAddress[26] ;
 wire \core.csr.instruction_memoryAddress[27] ;
 wire \core.csr.instruction_memoryAddress[28] ;
 wire \core.csr.instruction_memoryAddress[29] ;
 wire \core.csr.instruction_memoryAddress[2] ;
 wire \core.csr.instruction_memoryAddress[30] ;
 wire \core.csr.instruction_memoryAddress[31] ;
 wire \core.csr.instruction_memoryAddress[3] ;
 wire \core.csr.instruction_memoryAddress[4] ;
 wire \core.csr.instruction_memoryAddress[5] ;
 wire \core.csr.instruction_memoryAddress[6] ;
 wire \core.csr.instruction_memoryAddress[7] ;
 wire \core.csr.instruction_memoryAddress[8] ;
 wire \core.csr.instruction_memoryAddress[9] ;
 wire \core.csr.mconfigptr.currentValue[0] ;
 wire \core.csr.mconfigptr.currentValue[10] ;
 wire \core.csr.mconfigptr.currentValue[11] ;
 wire \core.csr.mconfigptr.currentValue[12] ;
 wire \core.csr.mconfigptr.currentValue[13] ;
 wire \core.csr.mconfigptr.currentValue[14] ;
 wire \core.csr.mconfigptr.currentValue[15] ;
 wire \core.csr.mconfigptr.currentValue[16] ;
 wire \core.csr.mconfigptr.currentValue[17] ;
 wire \core.csr.mconfigptr.currentValue[18] ;
 wire \core.csr.mconfigptr.currentValue[19] ;
 wire \core.csr.mconfigptr.currentValue[1] ;
 wire \core.csr.mconfigptr.currentValue[20] ;
 wire \core.csr.mconfigptr.currentValue[21] ;
 wire \core.csr.mconfigptr.currentValue[22] ;
 wire \core.csr.mconfigptr.currentValue[23] ;
 wire \core.csr.mconfigptr.currentValue[24] ;
 wire \core.csr.mconfigptr.currentValue[25] ;
 wire \core.csr.mconfigptr.currentValue[26] ;
 wire \core.csr.mconfigptr.currentValue[27] ;
 wire \core.csr.mconfigptr.currentValue[28] ;
 wire \core.csr.mconfigptr.currentValue[29] ;
 wire \core.csr.mconfigptr.currentValue[2] ;
 wire \core.csr.mconfigptr.currentValue[30] ;
 wire \core.csr.mconfigptr.currentValue[31] ;
 wire \core.csr.mconfigptr.currentValue[3] ;
 wire \core.csr.mconfigptr.currentValue[4] ;
 wire \core.csr.mconfigptr.currentValue[5] ;
 wire \core.csr.mconfigptr.currentValue[6] ;
 wire \core.csr.mconfigptr.currentValue[7] ;
 wire \core.csr.mconfigptr.currentValue[8] ;
 wire \core.csr.mconfigptr.currentValue[9] ;
 wire \core.csr.trapReturnVector[0] ;
 wire \core.csr.trapReturnVector[10] ;
 wire \core.csr.trapReturnVector[11] ;
 wire \core.csr.trapReturnVector[12] ;
 wire \core.csr.trapReturnVector[13] ;
 wire \core.csr.trapReturnVector[14] ;
 wire \core.csr.trapReturnVector[15] ;
 wire \core.csr.trapReturnVector[16] ;
 wire \core.csr.trapReturnVector[17] ;
 wire \core.csr.trapReturnVector[18] ;
 wire \core.csr.trapReturnVector[19] ;
 wire \core.csr.trapReturnVector[1] ;
 wire \core.csr.trapReturnVector[20] ;
 wire \core.csr.trapReturnVector[21] ;
 wire \core.csr.trapReturnVector[22] ;
 wire \core.csr.trapReturnVector[23] ;
 wire \core.csr.trapReturnVector[24] ;
 wire \core.csr.trapReturnVector[25] ;
 wire \core.csr.trapReturnVector[26] ;
 wire \core.csr.trapReturnVector[27] ;
 wire \core.csr.trapReturnVector[28] ;
 wire \core.csr.trapReturnVector[29] ;
 wire \core.csr.trapReturnVector[2] ;
 wire \core.csr.trapReturnVector[30] ;
 wire \core.csr.trapReturnVector[31] ;
 wire \core.csr.trapReturnVector[3] ;
 wire \core.csr.trapReturnVector[4] ;
 wire \core.csr.trapReturnVector[5] ;
 wire \core.csr.trapReturnVector[6] ;
 wire \core.csr.trapReturnVector[7] ;
 wire \core.csr.trapReturnVector[8] ;
 wire \core.csr.trapReturnVector[9] ;
 wire \core.csr.traps.machineInterruptEnable ;
 wire \core.csr.traps.machinePreviousInterruptEnable ;
 wire \core.csr.traps.mcause.csrReadData[0] ;
 wire \core.csr.traps.mcause.csrReadData[10] ;
 wire \core.csr.traps.mcause.csrReadData[11] ;
 wire \core.csr.traps.mcause.csrReadData[12] ;
 wire \core.csr.traps.mcause.csrReadData[13] ;
 wire \core.csr.traps.mcause.csrReadData[14] ;
 wire \core.csr.traps.mcause.csrReadData[15] ;
 wire \core.csr.traps.mcause.csrReadData[16] ;
 wire \core.csr.traps.mcause.csrReadData[17] ;
 wire \core.csr.traps.mcause.csrReadData[18] ;
 wire \core.csr.traps.mcause.csrReadData[19] ;
 wire \core.csr.traps.mcause.csrReadData[1] ;
 wire \core.csr.traps.mcause.csrReadData[20] ;
 wire \core.csr.traps.mcause.csrReadData[21] ;
 wire \core.csr.traps.mcause.csrReadData[22] ;
 wire \core.csr.traps.mcause.csrReadData[23] ;
 wire \core.csr.traps.mcause.csrReadData[24] ;
 wire \core.csr.traps.mcause.csrReadData[25] ;
 wire \core.csr.traps.mcause.csrReadData[26] ;
 wire \core.csr.traps.mcause.csrReadData[27] ;
 wire \core.csr.traps.mcause.csrReadData[28] ;
 wire \core.csr.traps.mcause.csrReadData[29] ;
 wire \core.csr.traps.mcause.csrReadData[2] ;
 wire \core.csr.traps.mcause.csrReadData[30] ;
 wire \core.csr.traps.mcause.csrReadData[31] ;
 wire \core.csr.traps.mcause.csrReadData[3] ;
 wire \core.csr.traps.mcause.csrReadData[4] ;
 wire \core.csr.traps.mcause.csrReadData[5] ;
 wire \core.csr.traps.mcause.csrReadData[6] ;
 wire \core.csr.traps.mcause.csrReadData[7] ;
 wire \core.csr.traps.mcause.csrReadData[8] ;
 wire \core.csr.traps.mcause.csrReadData[9] ;
 wire \core.csr.traps.mie.currentValue[0] ;
 wire \core.csr.traps.mie.currentValue[10] ;
 wire \core.csr.traps.mie.currentValue[11] ;
 wire \core.csr.traps.mie.currentValue[12] ;
 wire \core.csr.traps.mie.currentValue[13] ;
 wire \core.csr.traps.mie.currentValue[14] ;
 wire \core.csr.traps.mie.currentValue[15] ;
 wire \core.csr.traps.mie.currentValue[16] ;
 wire \core.csr.traps.mie.currentValue[17] ;
 wire \core.csr.traps.mie.currentValue[18] ;
 wire \core.csr.traps.mie.currentValue[19] ;
 wire \core.csr.traps.mie.currentValue[1] ;
 wire \core.csr.traps.mie.currentValue[20] ;
 wire \core.csr.traps.mie.currentValue[21] ;
 wire \core.csr.traps.mie.currentValue[22] ;
 wire \core.csr.traps.mie.currentValue[23] ;
 wire \core.csr.traps.mie.currentValue[24] ;
 wire \core.csr.traps.mie.currentValue[25] ;
 wire \core.csr.traps.mie.currentValue[26] ;
 wire \core.csr.traps.mie.currentValue[27] ;
 wire \core.csr.traps.mie.currentValue[28] ;
 wire \core.csr.traps.mie.currentValue[29] ;
 wire \core.csr.traps.mie.currentValue[2] ;
 wire \core.csr.traps.mie.currentValue[30] ;
 wire \core.csr.traps.mie.currentValue[31] ;
 wire \core.csr.traps.mie.currentValue[3] ;
 wire \core.csr.traps.mie.currentValue[4] ;
 wire \core.csr.traps.mie.currentValue[5] ;
 wire \core.csr.traps.mie.currentValue[6] ;
 wire \core.csr.traps.mie.currentValue[7] ;
 wire \core.csr.traps.mie.currentValue[8] ;
 wire \core.csr.traps.mie.currentValue[9] ;
 wire \core.csr.traps.mip.csrReadData[0] ;
 wire \core.csr.traps.mip.csrReadData[10] ;
 wire \core.csr.traps.mip.csrReadData[11] ;
 wire \core.csr.traps.mip.csrReadData[12] ;
 wire \core.csr.traps.mip.csrReadData[13] ;
 wire \core.csr.traps.mip.csrReadData[14] ;
 wire \core.csr.traps.mip.csrReadData[15] ;
 wire \core.csr.traps.mip.csrReadData[16] ;
 wire \core.csr.traps.mip.csrReadData[17] ;
 wire \core.csr.traps.mip.csrReadData[18] ;
 wire \core.csr.traps.mip.csrReadData[19] ;
 wire \core.csr.traps.mip.csrReadData[1] ;
 wire \core.csr.traps.mip.csrReadData[20] ;
 wire \core.csr.traps.mip.csrReadData[21] ;
 wire \core.csr.traps.mip.csrReadData[22] ;
 wire \core.csr.traps.mip.csrReadData[23] ;
 wire \core.csr.traps.mip.csrReadData[24] ;
 wire \core.csr.traps.mip.csrReadData[25] ;
 wire \core.csr.traps.mip.csrReadData[26] ;
 wire \core.csr.traps.mip.csrReadData[27] ;
 wire \core.csr.traps.mip.csrReadData[28] ;
 wire \core.csr.traps.mip.csrReadData[29] ;
 wire \core.csr.traps.mip.csrReadData[2] ;
 wire \core.csr.traps.mip.csrReadData[30] ;
 wire \core.csr.traps.mip.csrReadData[31] ;
 wire \core.csr.traps.mip.csrReadData[3] ;
 wire \core.csr.traps.mip.csrReadData[4] ;
 wire \core.csr.traps.mip.csrReadData[5] ;
 wire \core.csr.traps.mip.csrReadData[6] ;
 wire \core.csr.traps.mip.csrReadData[7] ;
 wire \core.csr.traps.mip.csrReadData[8] ;
 wire \core.csr.traps.mip.csrReadData[9] ;
 wire \core.csr.traps.mscratch.currentValue[0] ;
 wire \core.csr.traps.mscratch.currentValue[10] ;
 wire \core.csr.traps.mscratch.currentValue[11] ;
 wire \core.csr.traps.mscratch.currentValue[12] ;
 wire \core.csr.traps.mscratch.currentValue[13] ;
 wire \core.csr.traps.mscratch.currentValue[14] ;
 wire \core.csr.traps.mscratch.currentValue[15] ;
 wire \core.csr.traps.mscratch.currentValue[16] ;
 wire \core.csr.traps.mscratch.currentValue[17] ;
 wire \core.csr.traps.mscratch.currentValue[18] ;
 wire \core.csr.traps.mscratch.currentValue[19] ;
 wire \core.csr.traps.mscratch.currentValue[1] ;
 wire \core.csr.traps.mscratch.currentValue[20] ;
 wire \core.csr.traps.mscratch.currentValue[21] ;
 wire \core.csr.traps.mscratch.currentValue[22] ;
 wire \core.csr.traps.mscratch.currentValue[23] ;
 wire \core.csr.traps.mscratch.currentValue[24] ;
 wire \core.csr.traps.mscratch.currentValue[25] ;
 wire \core.csr.traps.mscratch.currentValue[26] ;
 wire \core.csr.traps.mscratch.currentValue[27] ;
 wire \core.csr.traps.mscratch.currentValue[28] ;
 wire \core.csr.traps.mscratch.currentValue[29] ;
 wire \core.csr.traps.mscratch.currentValue[2] ;
 wire \core.csr.traps.mscratch.currentValue[30] ;
 wire \core.csr.traps.mscratch.currentValue[31] ;
 wire \core.csr.traps.mscratch.currentValue[3] ;
 wire \core.csr.traps.mscratch.currentValue[4] ;
 wire \core.csr.traps.mscratch.currentValue[5] ;
 wire \core.csr.traps.mscratch.currentValue[6] ;
 wire \core.csr.traps.mscratch.currentValue[7] ;
 wire \core.csr.traps.mscratch.currentValue[8] ;
 wire \core.csr.traps.mscratch.currentValue[9] ;
 wire \core.csr.traps.mtval.csrReadData[0] ;
 wire \core.csr.traps.mtval.csrReadData[10] ;
 wire \core.csr.traps.mtval.csrReadData[11] ;
 wire \core.csr.traps.mtval.csrReadData[12] ;
 wire \core.csr.traps.mtval.csrReadData[13] ;
 wire \core.csr.traps.mtval.csrReadData[14] ;
 wire \core.csr.traps.mtval.csrReadData[15] ;
 wire \core.csr.traps.mtval.csrReadData[16] ;
 wire \core.csr.traps.mtval.csrReadData[17] ;
 wire \core.csr.traps.mtval.csrReadData[18] ;
 wire \core.csr.traps.mtval.csrReadData[19] ;
 wire \core.csr.traps.mtval.csrReadData[1] ;
 wire \core.csr.traps.mtval.csrReadData[20] ;
 wire \core.csr.traps.mtval.csrReadData[21] ;
 wire \core.csr.traps.mtval.csrReadData[22] ;
 wire \core.csr.traps.mtval.csrReadData[23] ;
 wire \core.csr.traps.mtval.csrReadData[24] ;
 wire \core.csr.traps.mtval.csrReadData[25] ;
 wire \core.csr.traps.mtval.csrReadData[26] ;
 wire \core.csr.traps.mtval.csrReadData[27] ;
 wire \core.csr.traps.mtval.csrReadData[28] ;
 wire \core.csr.traps.mtval.csrReadData[29] ;
 wire \core.csr.traps.mtval.csrReadData[2] ;
 wire \core.csr.traps.mtval.csrReadData[30] ;
 wire \core.csr.traps.mtval.csrReadData[31] ;
 wire \core.csr.traps.mtval.csrReadData[3] ;
 wire \core.csr.traps.mtval.csrReadData[4] ;
 wire \core.csr.traps.mtval.csrReadData[5] ;
 wire \core.csr.traps.mtval.csrReadData[6] ;
 wire \core.csr.traps.mtval.csrReadData[7] ;
 wire \core.csr.traps.mtval.csrReadData[8] ;
 wire \core.csr.traps.mtval.csrReadData[9] ;
 wire \core.csr.traps.mtvec.csrReadData[0] ;
 wire \core.csr.traps.mtvec.csrReadData[10] ;
 wire \core.csr.traps.mtvec.csrReadData[11] ;
 wire \core.csr.traps.mtvec.csrReadData[12] ;
 wire \core.csr.traps.mtvec.csrReadData[13] ;
 wire \core.csr.traps.mtvec.csrReadData[14] ;
 wire \core.csr.traps.mtvec.csrReadData[15] ;
 wire \core.csr.traps.mtvec.csrReadData[16] ;
 wire \core.csr.traps.mtvec.csrReadData[17] ;
 wire \core.csr.traps.mtvec.csrReadData[18] ;
 wire \core.csr.traps.mtvec.csrReadData[19] ;
 wire \core.csr.traps.mtvec.csrReadData[1] ;
 wire \core.csr.traps.mtvec.csrReadData[20] ;
 wire \core.csr.traps.mtvec.csrReadData[21] ;
 wire \core.csr.traps.mtvec.csrReadData[22] ;
 wire \core.csr.traps.mtvec.csrReadData[23] ;
 wire \core.csr.traps.mtvec.csrReadData[24] ;
 wire \core.csr.traps.mtvec.csrReadData[25] ;
 wire \core.csr.traps.mtvec.csrReadData[26] ;
 wire \core.csr.traps.mtvec.csrReadData[27] ;
 wire \core.csr.traps.mtvec.csrReadData[28] ;
 wire \core.csr.traps.mtvec.csrReadData[29] ;
 wire \core.csr.traps.mtvec.csrReadData[2] ;
 wire \core.csr.traps.mtvec.csrReadData[30] ;
 wire \core.csr.traps.mtvec.csrReadData[31] ;
 wire \core.csr.traps.mtvec.csrReadData[3] ;
 wire \core.csr.traps.mtvec.csrReadData[4] ;
 wire \core.csr.traps.mtvec.csrReadData[5] ;
 wire \core.csr.traps.mtvec.csrReadData[6] ;
 wire \core.csr.traps.mtvec.csrReadData[7] ;
 wire \core.csr.traps.mtvec.csrReadData[8] ;
 wire \core.csr.traps.mtvec.csrReadData[9] ;
 wire \core.fetchProgramCounter[0] ;
 wire \core.fetchProgramCounter[10] ;
 wire \core.fetchProgramCounter[11] ;
 wire \core.fetchProgramCounter[12] ;
 wire \core.fetchProgramCounter[13] ;
 wire \core.fetchProgramCounter[14] ;
 wire \core.fetchProgramCounter[15] ;
 wire \core.fetchProgramCounter[16] ;
 wire \core.fetchProgramCounter[17] ;
 wire \core.fetchProgramCounter[18] ;
 wire \core.fetchProgramCounter[19] ;
 wire \core.fetchProgramCounter[1] ;
 wire \core.fetchProgramCounter[20] ;
 wire \core.fetchProgramCounter[21] ;
 wire \core.fetchProgramCounter[22] ;
 wire \core.fetchProgramCounter[23] ;
 wire \core.fetchProgramCounter[24] ;
 wire \core.fetchProgramCounter[25] ;
 wire \core.fetchProgramCounter[26] ;
 wire \core.fetchProgramCounter[27] ;
 wire \core.fetchProgramCounter[28] ;
 wire \core.fetchProgramCounter[29] ;
 wire \core.fetchProgramCounter[2] ;
 wire \core.fetchProgramCounter[30] ;
 wire \core.fetchProgramCounter[31] ;
 wire \core.fetchProgramCounter[3] ;
 wire \core.fetchProgramCounter[4] ;
 wire \core.fetchProgramCounter[5] ;
 wire \core.fetchProgramCounter[6] ;
 wire \core.fetchProgramCounter[7] ;
 wire \core.fetchProgramCounter[8] ;
 wire \core.fetchProgramCounter[9] ;
 wire \core.management_interruptEnable ;
 wire \core.management_pipeStartup ;
 wire \core.management_run ;
 wire \core.memoryOperationCompleted ;
 wire \core.pipe0_currentInstruction[0] ;
 wire \core.pipe0_currentInstruction[10] ;
 wire \core.pipe0_currentInstruction[11] ;
 wire \core.pipe0_currentInstruction[12] ;
 wire \core.pipe0_currentInstruction[13] ;
 wire \core.pipe0_currentInstruction[14] ;
 wire \core.pipe0_currentInstruction[15] ;
 wire \core.pipe0_currentInstruction[16] ;
 wire \core.pipe0_currentInstruction[17] ;
 wire \core.pipe0_currentInstruction[18] ;
 wire \core.pipe0_currentInstruction[19] ;
 wire \core.pipe0_currentInstruction[1] ;
 wire \core.pipe0_currentInstruction[20] ;
 wire \core.pipe0_currentInstruction[21] ;
 wire \core.pipe0_currentInstruction[22] ;
 wire \core.pipe0_currentInstruction[23] ;
 wire \core.pipe0_currentInstruction[24] ;
 wire \core.pipe0_currentInstruction[25] ;
 wire \core.pipe0_currentInstruction[26] ;
 wire \core.pipe0_currentInstruction[27] ;
 wire \core.pipe0_currentInstruction[28] ;
 wire \core.pipe0_currentInstruction[29] ;
 wire \core.pipe0_currentInstruction[2] ;
 wire \core.pipe0_currentInstruction[30] ;
 wire \core.pipe0_currentInstruction[31] ;
 wire \core.pipe0_currentInstruction[3] ;
 wire \core.pipe0_currentInstruction[4] ;
 wire \core.pipe0_currentInstruction[5] ;
 wire \core.pipe0_currentInstruction[6] ;
 wire \core.pipe0_currentInstruction[7] ;
 wire \core.pipe0_currentInstruction[8] ;
 wire \core.pipe0_currentInstruction[9] ;
 wire \core.pipe0_fetch.cachedInstruction[0] ;
 wire \core.pipe0_fetch.cachedInstruction[10] ;
 wire \core.pipe0_fetch.cachedInstruction[11] ;
 wire \core.pipe0_fetch.cachedInstruction[12] ;
 wire \core.pipe0_fetch.cachedInstruction[13] ;
 wire \core.pipe0_fetch.cachedInstruction[14] ;
 wire \core.pipe0_fetch.cachedInstruction[15] ;
 wire \core.pipe0_fetch.cachedInstruction[16] ;
 wire \core.pipe0_fetch.cachedInstruction[17] ;
 wire \core.pipe0_fetch.cachedInstruction[18] ;
 wire \core.pipe0_fetch.cachedInstruction[19] ;
 wire \core.pipe0_fetch.cachedInstruction[1] ;
 wire \core.pipe0_fetch.cachedInstruction[20] ;
 wire \core.pipe0_fetch.cachedInstruction[21] ;
 wire \core.pipe0_fetch.cachedInstruction[22] ;
 wire \core.pipe0_fetch.cachedInstruction[23] ;
 wire \core.pipe0_fetch.cachedInstruction[24] ;
 wire \core.pipe0_fetch.cachedInstruction[25] ;
 wire \core.pipe0_fetch.cachedInstruction[26] ;
 wire \core.pipe0_fetch.cachedInstruction[27] ;
 wire \core.pipe0_fetch.cachedInstruction[28] ;
 wire \core.pipe0_fetch.cachedInstruction[29] ;
 wire \core.pipe0_fetch.cachedInstruction[2] ;
 wire \core.pipe0_fetch.cachedInstruction[30] ;
 wire \core.pipe0_fetch.cachedInstruction[31] ;
 wire \core.pipe0_fetch.cachedInstruction[3] ;
 wire \core.pipe0_fetch.cachedInstruction[4] ;
 wire \core.pipe0_fetch.cachedInstruction[5] ;
 wire \core.pipe0_fetch.cachedInstruction[6] ;
 wire \core.pipe0_fetch.cachedInstruction[7] ;
 wire \core.pipe0_fetch.cachedInstruction[8] ;
 wire \core.pipe0_fetch.cachedInstruction[9] ;
 wire \core.pipe0_fetch.currentPipeStall ;
 wire \core.pipe0_fetch.instructionCached ;
 wire \core.pipe1_csrData[0] ;
 wire \core.pipe1_csrData[10] ;
 wire \core.pipe1_csrData[11] ;
 wire \core.pipe1_csrData[12] ;
 wire \core.pipe1_csrData[13] ;
 wire \core.pipe1_csrData[14] ;
 wire \core.pipe1_csrData[15] ;
 wire \core.pipe1_csrData[16] ;
 wire \core.pipe1_csrData[17] ;
 wire \core.pipe1_csrData[18] ;
 wire \core.pipe1_csrData[19] ;
 wire \core.pipe1_csrData[1] ;
 wire \core.pipe1_csrData[20] ;
 wire \core.pipe1_csrData[21] ;
 wire \core.pipe1_csrData[22] ;
 wire \core.pipe1_csrData[23] ;
 wire \core.pipe1_csrData[24] ;
 wire \core.pipe1_csrData[25] ;
 wire \core.pipe1_csrData[26] ;
 wire \core.pipe1_csrData[27] ;
 wire \core.pipe1_csrData[28] ;
 wire \core.pipe1_csrData[29] ;
 wire \core.pipe1_csrData[2] ;
 wire \core.pipe1_csrData[30] ;
 wire \core.pipe1_csrData[31] ;
 wire \core.pipe1_csrData[3] ;
 wire \core.pipe1_csrData[4] ;
 wire \core.pipe1_csrData[5] ;
 wire \core.pipe1_csrData[6] ;
 wire \core.pipe1_csrData[7] ;
 wire \core.pipe1_csrData[8] ;
 wire \core.pipe1_csrData[9] ;
 wire \core.pipe1_loadResult[0] ;
 wire \core.pipe1_loadResult[10] ;
 wire \core.pipe1_loadResult[11] ;
 wire \core.pipe1_loadResult[12] ;
 wire \core.pipe1_loadResult[13] ;
 wire \core.pipe1_loadResult[14] ;
 wire \core.pipe1_loadResult[15] ;
 wire \core.pipe1_loadResult[16] ;
 wire \core.pipe1_loadResult[17] ;
 wire \core.pipe1_loadResult[18] ;
 wire \core.pipe1_loadResult[19] ;
 wire \core.pipe1_loadResult[1] ;
 wire \core.pipe1_loadResult[20] ;
 wire \core.pipe1_loadResult[21] ;
 wire \core.pipe1_loadResult[22] ;
 wire \core.pipe1_loadResult[23] ;
 wire \core.pipe1_loadResult[24] ;
 wire \core.pipe1_loadResult[25] ;
 wire \core.pipe1_loadResult[26] ;
 wire \core.pipe1_loadResult[27] ;
 wire \core.pipe1_loadResult[28] ;
 wire \core.pipe1_loadResult[29] ;
 wire \core.pipe1_loadResult[2] ;
 wire \core.pipe1_loadResult[30] ;
 wire \core.pipe1_loadResult[31] ;
 wire \core.pipe1_loadResult[3] ;
 wire \core.pipe1_loadResult[4] ;
 wire \core.pipe1_loadResult[5] ;
 wire \core.pipe1_loadResult[6] ;
 wire \core.pipe1_loadResult[7] ;
 wire \core.pipe1_loadResult[8] ;
 wire \core.pipe1_loadResult[9] ;
 wire \core.pipe1_operation.currentPipeStall ;
 wire \core.pipe1_resultRegister[0] ;
 wire \core.pipe1_resultRegister[10] ;
 wire \core.pipe1_resultRegister[11] ;
 wire \core.pipe1_resultRegister[12] ;
 wire \core.pipe1_resultRegister[13] ;
 wire \core.pipe1_resultRegister[14] ;
 wire \core.pipe1_resultRegister[15] ;
 wire \core.pipe1_resultRegister[16] ;
 wire \core.pipe1_resultRegister[17] ;
 wire \core.pipe1_resultRegister[18] ;
 wire \core.pipe1_resultRegister[19] ;
 wire \core.pipe1_resultRegister[1] ;
 wire \core.pipe1_resultRegister[20] ;
 wire \core.pipe1_resultRegister[21] ;
 wire \core.pipe1_resultRegister[22] ;
 wire \core.pipe1_resultRegister[23] ;
 wire \core.pipe1_resultRegister[24] ;
 wire \core.pipe1_resultRegister[25] ;
 wire \core.pipe1_resultRegister[26] ;
 wire \core.pipe1_resultRegister[27] ;
 wire \core.pipe1_resultRegister[28] ;
 wire \core.pipe1_resultRegister[29] ;
 wire \core.pipe1_resultRegister[2] ;
 wire \core.pipe1_resultRegister[30] ;
 wire \core.pipe1_resultRegister[31] ;
 wire \core.pipe1_resultRegister[3] ;
 wire \core.pipe1_resultRegister[4] ;
 wire \core.pipe1_resultRegister[5] ;
 wire \core.pipe1_resultRegister[6] ;
 wire \core.pipe1_resultRegister[7] ;
 wire \core.pipe1_resultRegister[8] ;
 wire \core.pipe1_resultRegister[9] ;
 wire \core.pipe2_stall ;
 wire \core.registers[0][0] ;
 wire \core.registers[0][10] ;
 wire \core.registers[0][11] ;
 wire \core.registers[0][12] ;
 wire \core.registers[0][13] ;
 wire \core.registers[0][14] ;
 wire \core.registers[0][15] ;
 wire \core.registers[0][16] ;
 wire \core.registers[0][17] ;
 wire \core.registers[0][18] ;
 wire \core.registers[0][19] ;
 wire \core.registers[0][1] ;
 wire \core.registers[0][20] ;
 wire \core.registers[0][21] ;
 wire \core.registers[0][22] ;
 wire \core.registers[0][23] ;
 wire \core.registers[0][24] ;
 wire \core.registers[0][25] ;
 wire \core.registers[0][26] ;
 wire \core.registers[0][27] ;
 wire \core.registers[0][28] ;
 wire \core.registers[0][29] ;
 wire \core.registers[0][2] ;
 wire \core.registers[0][30] ;
 wire \core.registers[0][31] ;
 wire \core.registers[0][3] ;
 wire \core.registers[0][4] ;
 wire \core.registers[0][5] ;
 wire \core.registers[0][6] ;
 wire \core.registers[0][7] ;
 wire \core.registers[0][8] ;
 wire \core.registers[0][9] ;
 wire \core.registers[10][0] ;
 wire \core.registers[10][10] ;
 wire \core.registers[10][11] ;
 wire \core.registers[10][12] ;
 wire \core.registers[10][13] ;
 wire \core.registers[10][14] ;
 wire \core.registers[10][15] ;
 wire \core.registers[10][16] ;
 wire \core.registers[10][17] ;
 wire \core.registers[10][18] ;
 wire \core.registers[10][19] ;
 wire \core.registers[10][1] ;
 wire \core.registers[10][20] ;
 wire \core.registers[10][21] ;
 wire \core.registers[10][22] ;
 wire \core.registers[10][23] ;
 wire \core.registers[10][24] ;
 wire \core.registers[10][25] ;
 wire \core.registers[10][26] ;
 wire \core.registers[10][27] ;
 wire \core.registers[10][28] ;
 wire \core.registers[10][29] ;
 wire \core.registers[10][2] ;
 wire \core.registers[10][30] ;
 wire \core.registers[10][31] ;
 wire \core.registers[10][3] ;
 wire \core.registers[10][4] ;
 wire \core.registers[10][5] ;
 wire \core.registers[10][6] ;
 wire \core.registers[10][7] ;
 wire \core.registers[10][8] ;
 wire \core.registers[10][9] ;
 wire \core.registers[11][0] ;
 wire \core.registers[11][10] ;
 wire \core.registers[11][11] ;
 wire \core.registers[11][12] ;
 wire \core.registers[11][13] ;
 wire \core.registers[11][14] ;
 wire \core.registers[11][15] ;
 wire \core.registers[11][16] ;
 wire \core.registers[11][17] ;
 wire \core.registers[11][18] ;
 wire \core.registers[11][19] ;
 wire \core.registers[11][1] ;
 wire \core.registers[11][20] ;
 wire \core.registers[11][21] ;
 wire \core.registers[11][22] ;
 wire \core.registers[11][23] ;
 wire \core.registers[11][24] ;
 wire \core.registers[11][25] ;
 wire \core.registers[11][26] ;
 wire \core.registers[11][27] ;
 wire \core.registers[11][28] ;
 wire \core.registers[11][29] ;
 wire \core.registers[11][2] ;
 wire \core.registers[11][30] ;
 wire \core.registers[11][31] ;
 wire \core.registers[11][3] ;
 wire \core.registers[11][4] ;
 wire \core.registers[11][5] ;
 wire \core.registers[11][6] ;
 wire \core.registers[11][7] ;
 wire \core.registers[11][8] ;
 wire \core.registers[11][9] ;
 wire \core.registers[12][0] ;
 wire \core.registers[12][10] ;
 wire \core.registers[12][11] ;
 wire \core.registers[12][12] ;
 wire \core.registers[12][13] ;
 wire \core.registers[12][14] ;
 wire \core.registers[12][15] ;
 wire \core.registers[12][16] ;
 wire \core.registers[12][17] ;
 wire \core.registers[12][18] ;
 wire \core.registers[12][19] ;
 wire \core.registers[12][1] ;
 wire \core.registers[12][20] ;
 wire \core.registers[12][21] ;
 wire \core.registers[12][22] ;
 wire \core.registers[12][23] ;
 wire \core.registers[12][24] ;
 wire \core.registers[12][25] ;
 wire \core.registers[12][26] ;
 wire \core.registers[12][27] ;
 wire \core.registers[12][28] ;
 wire \core.registers[12][29] ;
 wire \core.registers[12][2] ;
 wire \core.registers[12][30] ;
 wire \core.registers[12][31] ;
 wire \core.registers[12][3] ;
 wire \core.registers[12][4] ;
 wire \core.registers[12][5] ;
 wire \core.registers[12][6] ;
 wire \core.registers[12][7] ;
 wire \core.registers[12][8] ;
 wire \core.registers[12][9] ;
 wire \core.registers[13][0] ;
 wire \core.registers[13][10] ;
 wire \core.registers[13][11] ;
 wire \core.registers[13][12] ;
 wire \core.registers[13][13] ;
 wire \core.registers[13][14] ;
 wire \core.registers[13][15] ;
 wire \core.registers[13][16] ;
 wire \core.registers[13][17] ;
 wire \core.registers[13][18] ;
 wire \core.registers[13][19] ;
 wire \core.registers[13][1] ;
 wire \core.registers[13][20] ;
 wire \core.registers[13][21] ;
 wire \core.registers[13][22] ;
 wire \core.registers[13][23] ;
 wire \core.registers[13][24] ;
 wire \core.registers[13][25] ;
 wire \core.registers[13][26] ;
 wire \core.registers[13][27] ;
 wire \core.registers[13][28] ;
 wire \core.registers[13][29] ;
 wire \core.registers[13][2] ;
 wire \core.registers[13][30] ;
 wire \core.registers[13][31] ;
 wire \core.registers[13][3] ;
 wire \core.registers[13][4] ;
 wire \core.registers[13][5] ;
 wire \core.registers[13][6] ;
 wire \core.registers[13][7] ;
 wire \core.registers[13][8] ;
 wire \core.registers[13][9] ;
 wire \core.registers[14][0] ;
 wire \core.registers[14][10] ;
 wire \core.registers[14][11] ;
 wire \core.registers[14][12] ;
 wire \core.registers[14][13] ;
 wire \core.registers[14][14] ;
 wire \core.registers[14][15] ;
 wire \core.registers[14][16] ;
 wire \core.registers[14][17] ;
 wire \core.registers[14][18] ;
 wire \core.registers[14][19] ;
 wire \core.registers[14][1] ;
 wire \core.registers[14][20] ;
 wire \core.registers[14][21] ;
 wire \core.registers[14][22] ;
 wire \core.registers[14][23] ;
 wire \core.registers[14][24] ;
 wire \core.registers[14][25] ;
 wire \core.registers[14][26] ;
 wire \core.registers[14][27] ;
 wire \core.registers[14][28] ;
 wire \core.registers[14][29] ;
 wire \core.registers[14][2] ;
 wire \core.registers[14][30] ;
 wire \core.registers[14][31] ;
 wire \core.registers[14][3] ;
 wire \core.registers[14][4] ;
 wire \core.registers[14][5] ;
 wire \core.registers[14][6] ;
 wire \core.registers[14][7] ;
 wire \core.registers[14][8] ;
 wire \core.registers[14][9] ;
 wire \core.registers[15][0] ;
 wire \core.registers[15][10] ;
 wire \core.registers[15][11] ;
 wire \core.registers[15][12] ;
 wire \core.registers[15][13] ;
 wire \core.registers[15][14] ;
 wire \core.registers[15][15] ;
 wire \core.registers[15][16] ;
 wire \core.registers[15][17] ;
 wire \core.registers[15][18] ;
 wire \core.registers[15][19] ;
 wire \core.registers[15][1] ;
 wire \core.registers[15][20] ;
 wire \core.registers[15][21] ;
 wire \core.registers[15][22] ;
 wire \core.registers[15][23] ;
 wire \core.registers[15][24] ;
 wire \core.registers[15][25] ;
 wire \core.registers[15][26] ;
 wire \core.registers[15][27] ;
 wire \core.registers[15][28] ;
 wire \core.registers[15][29] ;
 wire \core.registers[15][2] ;
 wire \core.registers[15][30] ;
 wire \core.registers[15][31] ;
 wire \core.registers[15][3] ;
 wire \core.registers[15][4] ;
 wire \core.registers[15][5] ;
 wire \core.registers[15][6] ;
 wire \core.registers[15][7] ;
 wire \core.registers[15][8] ;
 wire \core.registers[15][9] ;
 wire \core.registers[16][0] ;
 wire \core.registers[16][10] ;
 wire \core.registers[16][11] ;
 wire \core.registers[16][12] ;
 wire \core.registers[16][13] ;
 wire \core.registers[16][14] ;
 wire \core.registers[16][15] ;
 wire \core.registers[16][16] ;
 wire \core.registers[16][17] ;
 wire \core.registers[16][18] ;
 wire \core.registers[16][19] ;
 wire \core.registers[16][1] ;
 wire \core.registers[16][20] ;
 wire \core.registers[16][21] ;
 wire \core.registers[16][22] ;
 wire \core.registers[16][23] ;
 wire \core.registers[16][24] ;
 wire \core.registers[16][25] ;
 wire \core.registers[16][26] ;
 wire \core.registers[16][27] ;
 wire \core.registers[16][28] ;
 wire \core.registers[16][29] ;
 wire \core.registers[16][2] ;
 wire \core.registers[16][30] ;
 wire \core.registers[16][31] ;
 wire \core.registers[16][3] ;
 wire \core.registers[16][4] ;
 wire \core.registers[16][5] ;
 wire \core.registers[16][6] ;
 wire \core.registers[16][7] ;
 wire \core.registers[16][8] ;
 wire \core.registers[16][9] ;
 wire \core.registers[17][0] ;
 wire \core.registers[17][10] ;
 wire \core.registers[17][11] ;
 wire \core.registers[17][12] ;
 wire \core.registers[17][13] ;
 wire \core.registers[17][14] ;
 wire \core.registers[17][15] ;
 wire \core.registers[17][16] ;
 wire \core.registers[17][17] ;
 wire \core.registers[17][18] ;
 wire \core.registers[17][19] ;
 wire \core.registers[17][1] ;
 wire \core.registers[17][20] ;
 wire \core.registers[17][21] ;
 wire \core.registers[17][22] ;
 wire \core.registers[17][23] ;
 wire \core.registers[17][24] ;
 wire \core.registers[17][25] ;
 wire \core.registers[17][26] ;
 wire \core.registers[17][27] ;
 wire \core.registers[17][28] ;
 wire \core.registers[17][29] ;
 wire \core.registers[17][2] ;
 wire \core.registers[17][30] ;
 wire \core.registers[17][31] ;
 wire \core.registers[17][3] ;
 wire \core.registers[17][4] ;
 wire \core.registers[17][5] ;
 wire \core.registers[17][6] ;
 wire \core.registers[17][7] ;
 wire \core.registers[17][8] ;
 wire \core.registers[17][9] ;
 wire \core.registers[18][0] ;
 wire \core.registers[18][10] ;
 wire \core.registers[18][11] ;
 wire \core.registers[18][12] ;
 wire \core.registers[18][13] ;
 wire \core.registers[18][14] ;
 wire \core.registers[18][15] ;
 wire \core.registers[18][16] ;
 wire \core.registers[18][17] ;
 wire \core.registers[18][18] ;
 wire \core.registers[18][19] ;
 wire \core.registers[18][1] ;
 wire \core.registers[18][20] ;
 wire \core.registers[18][21] ;
 wire \core.registers[18][22] ;
 wire \core.registers[18][23] ;
 wire \core.registers[18][24] ;
 wire \core.registers[18][25] ;
 wire \core.registers[18][26] ;
 wire \core.registers[18][27] ;
 wire \core.registers[18][28] ;
 wire \core.registers[18][29] ;
 wire \core.registers[18][2] ;
 wire \core.registers[18][30] ;
 wire \core.registers[18][31] ;
 wire \core.registers[18][3] ;
 wire \core.registers[18][4] ;
 wire \core.registers[18][5] ;
 wire \core.registers[18][6] ;
 wire \core.registers[18][7] ;
 wire \core.registers[18][8] ;
 wire \core.registers[18][9] ;
 wire \core.registers[19][0] ;
 wire \core.registers[19][10] ;
 wire \core.registers[19][11] ;
 wire \core.registers[19][12] ;
 wire \core.registers[19][13] ;
 wire \core.registers[19][14] ;
 wire \core.registers[19][15] ;
 wire \core.registers[19][16] ;
 wire \core.registers[19][17] ;
 wire \core.registers[19][18] ;
 wire \core.registers[19][19] ;
 wire \core.registers[19][1] ;
 wire \core.registers[19][20] ;
 wire \core.registers[19][21] ;
 wire \core.registers[19][22] ;
 wire \core.registers[19][23] ;
 wire \core.registers[19][24] ;
 wire \core.registers[19][25] ;
 wire \core.registers[19][26] ;
 wire \core.registers[19][27] ;
 wire \core.registers[19][28] ;
 wire \core.registers[19][29] ;
 wire \core.registers[19][2] ;
 wire \core.registers[19][30] ;
 wire \core.registers[19][31] ;
 wire \core.registers[19][3] ;
 wire \core.registers[19][4] ;
 wire \core.registers[19][5] ;
 wire \core.registers[19][6] ;
 wire \core.registers[19][7] ;
 wire \core.registers[19][8] ;
 wire \core.registers[19][9] ;
 wire \core.registers[1][0] ;
 wire \core.registers[1][10] ;
 wire \core.registers[1][11] ;
 wire \core.registers[1][12] ;
 wire \core.registers[1][13] ;
 wire \core.registers[1][14] ;
 wire \core.registers[1][15] ;
 wire \core.registers[1][16] ;
 wire \core.registers[1][17] ;
 wire \core.registers[1][18] ;
 wire \core.registers[1][19] ;
 wire \core.registers[1][1] ;
 wire \core.registers[1][20] ;
 wire \core.registers[1][21] ;
 wire \core.registers[1][22] ;
 wire \core.registers[1][23] ;
 wire \core.registers[1][24] ;
 wire \core.registers[1][25] ;
 wire \core.registers[1][26] ;
 wire \core.registers[1][27] ;
 wire \core.registers[1][28] ;
 wire \core.registers[1][29] ;
 wire \core.registers[1][2] ;
 wire \core.registers[1][30] ;
 wire \core.registers[1][31] ;
 wire \core.registers[1][3] ;
 wire \core.registers[1][4] ;
 wire \core.registers[1][5] ;
 wire \core.registers[1][6] ;
 wire \core.registers[1][7] ;
 wire \core.registers[1][8] ;
 wire \core.registers[1][9] ;
 wire \core.registers[20][0] ;
 wire \core.registers[20][10] ;
 wire \core.registers[20][11] ;
 wire \core.registers[20][12] ;
 wire \core.registers[20][13] ;
 wire \core.registers[20][14] ;
 wire \core.registers[20][15] ;
 wire \core.registers[20][16] ;
 wire \core.registers[20][17] ;
 wire \core.registers[20][18] ;
 wire \core.registers[20][19] ;
 wire \core.registers[20][1] ;
 wire \core.registers[20][20] ;
 wire \core.registers[20][21] ;
 wire \core.registers[20][22] ;
 wire \core.registers[20][23] ;
 wire \core.registers[20][24] ;
 wire \core.registers[20][25] ;
 wire \core.registers[20][26] ;
 wire \core.registers[20][27] ;
 wire \core.registers[20][28] ;
 wire \core.registers[20][29] ;
 wire \core.registers[20][2] ;
 wire \core.registers[20][30] ;
 wire \core.registers[20][31] ;
 wire \core.registers[20][3] ;
 wire \core.registers[20][4] ;
 wire \core.registers[20][5] ;
 wire \core.registers[20][6] ;
 wire \core.registers[20][7] ;
 wire \core.registers[20][8] ;
 wire \core.registers[20][9] ;
 wire \core.registers[21][0] ;
 wire \core.registers[21][10] ;
 wire \core.registers[21][11] ;
 wire \core.registers[21][12] ;
 wire \core.registers[21][13] ;
 wire \core.registers[21][14] ;
 wire \core.registers[21][15] ;
 wire \core.registers[21][16] ;
 wire \core.registers[21][17] ;
 wire \core.registers[21][18] ;
 wire \core.registers[21][19] ;
 wire \core.registers[21][1] ;
 wire \core.registers[21][20] ;
 wire \core.registers[21][21] ;
 wire \core.registers[21][22] ;
 wire \core.registers[21][23] ;
 wire \core.registers[21][24] ;
 wire \core.registers[21][25] ;
 wire \core.registers[21][26] ;
 wire \core.registers[21][27] ;
 wire \core.registers[21][28] ;
 wire \core.registers[21][29] ;
 wire \core.registers[21][2] ;
 wire \core.registers[21][30] ;
 wire \core.registers[21][31] ;
 wire \core.registers[21][3] ;
 wire \core.registers[21][4] ;
 wire \core.registers[21][5] ;
 wire \core.registers[21][6] ;
 wire \core.registers[21][7] ;
 wire \core.registers[21][8] ;
 wire \core.registers[21][9] ;
 wire \core.registers[22][0] ;
 wire \core.registers[22][10] ;
 wire \core.registers[22][11] ;
 wire \core.registers[22][12] ;
 wire \core.registers[22][13] ;
 wire \core.registers[22][14] ;
 wire \core.registers[22][15] ;
 wire \core.registers[22][16] ;
 wire \core.registers[22][17] ;
 wire \core.registers[22][18] ;
 wire \core.registers[22][19] ;
 wire \core.registers[22][1] ;
 wire \core.registers[22][20] ;
 wire \core.registers[22][21] ;
 wire \core.registers[22][22] ;
 wire \core.registers[22][23] ;
 wire \core.registers[22][24] ;
 wire \core.registers[22][25] ;
 wire \core.registers[22][26] ;
 wire \core.registers[22][27] ;
 wire \core.registers[22][28] ;
 wire \core.registers[22][29] ;
 wire \core.registers[22][2] ;
 wire \core.registers[22][30] ;
 wire \core.registers[22][31] ;
 wire \core.registers[22][3] ;
 wire \core.registers[22][4] ;
 wire \core.registers[22][5] ;
 wire \core.registers[22][6] ;
 wire \core.registers[22][7] ;
 wire \core.registers[22][8] ;
 wire \core.registers[22][9] ;
 wire \core.registers[23][0] ;
 wire \core.registers[23][10] ;
 wire \core.registers[23][11] ;
 wire \core.registers[23][12] ;
 wire \core.registers[23][13] ;
 wire \core.registers[23][14] ;
 wire \core.registers[23][15] ;
 wire \core.registers[23][16] ;
 wire \core.registers[23][17] ;
 wire \core.registers[23][18] ;
 wire \core.registers[23][19] ;
 wire \core.registers[23][1] ;
 wire \core.registers[23][20] ;
 wire \core.registers[23][21] ;
 wire \core.registers[23][22] ;
 wire \core.registers[23][23] ;
 wire \core.registers[23][24] ;
 wire \core.registers[23][25] ;
 wire \core.registers[23][26] ;
 wire \core.registers[23][27] ;
 wire \core.registers[23][28] ;
 wire \core.registers[23][29] ;
 wire \core.registers[23][2] ;
 wire \core.registers[23][30] ;
 wire \core.registers[23][31] ;
 wire \core.registers[23][3] ;
 wire \core.registers[23][4] ;
 wire \core.registers[23][5] ;
 wire \core.registers[23][6] ;
 wire \core.registers[23][7] ;
 wire \core.registers[23][8] ;
 wire \core.registers[23][9] ;
 wire \core.registers[24][0] ;
 wire \core.registers[24][10] ;
 wire \core.registers[24][11] ;
 wire \core.registers[24][12] ;
 wire \core.registers[24][13] ;
 wire \core.registers[24][14] ;
 wire \core.registers[24][15] ;
 wire \core.registers[24][16] ;
 wire \core.registers[24][17] ;
 wire \core.registers[24][18] ;
 wire \core.registers[24][19] ;
 wire \core.registers[24][1] ;
 wire \core.registers[24][20] ;
 wire \core.registers[24][21] ;
 wire \core.registers[24][22] ;
 wire \core.registers[24][23] ;
 wire \core.registers[24][24] ;
 wire \core.registers[24][25] ;
 wire \core.registers[24][26] ;
 wire \core.registers[24][27] ;
 wire \core.registers[24][28] ;
 wire \core.registers[24][29] ;
 wire \core.registers[24][2] ;
 wire \core.registers[24][30] ;
 wire \core.registers[24][31] ;
 wire \core.registers[24][3] ;
 wire \core.registers[24][4] ;
 wire \core.registers[24][5] ;
 wire \core.registers[24][6] ;
 wire \core.registers[24][7] ;
 wire \core.registers[24][8] ;
 wire \core.registers[24][9] ;
 wire \core.registers[25][0] ;
 wire \core.registers[25][10] ;
 wire \core.registers[25][11] ;
 wire \core.registers[25][12] ;
 wire \core.registers[25][13] ;
 wire \core.registers[25][14] ;
 wire \core.registers[25][15] ;
 wire \core.registers[25][16] ;
 wire \core.registers[25][17] ;
 wire \core.registers[25][18] ;
 wire \core.registers[25][19] ;
 wire \core.registers[25][1] ;
 wire \core.registers[25][20] ;
 wire \core.registers[25][21] ;
 wire \core.registers[25][22] ;
 wire \core.registers[25][23] ;
 wire \core.registers[25][24] ;
 wire \core.registers[25][25] ;
 wire \core.registers[25][26] ;
 wire \core.registers[25][27] ;
 wire \core.registers[25][28] ;
 wire \core.registers[25][29] ;
 wire \core.registers[25][2] ;
 wire \core.registers[25][30] ;
 wire \core.registers[25][31] ;
 wire \core.registers[25][3] ;
 wire \core.registers[25][4] ;
 wire \core.registers[25][5] ;
 wire \core.registers[25][6] ;
 wire \core.registers[25][7] ;
 wire \core.registers[25][8] ;
 wire \core.registers[25][9] ;
 wire \core.registers[26][0] ;
 wire \core.registers[26][10] ;
 wire \core.registers[26][11] ;
 wire \core.registers[26][12] ;
 wire \core.registers[26][13] ;
 wire \core.registers[26][14] ;
 wire \core.registers[26][15] ;
 wire \core.registers[26][16] ;
 wire \core.registers[26][17] ;
 wire \core.registers[26][18] ;
 wire \core.registers[26][19] ;
 wire \core.registers[26][1] ;
 wire \core.registers[26][20] ;
 wire \core.registers[26][21] ;
 wire \core.registers[26][22] ;
 wire \core.registers[26][23] ;
 wire \core.registers[26][24] ;
 wire \core.registers[26][25] ;
 wire \core.registers[26][26] ;
 wire \core.registers[26][27] ;
 wire \core.registers[26][28] ;
 wire \core.registers[26][29] ;
 wire \core.registers[26][2] ;
 wire \core.registers[26][30] ;
 wire \core.registers[26][31] ;
 wire \core.registers[26][3] ;
 wire \core.registers[26][4] ;
 wire \core.registers[26][5] ;
 wire \core.registers[26][6] ;
 wire \core.registers[26][7] ;
 wire \core.registers[26][8] ;
 wire \core.registers[26][9] ;
 wire \core.registers[27][0] ;
 wire \core.registers[27][10] ;
 wire \core.registers[27][11] ;
 wire \core.registers[27][12] ;
 wire \core.registers[27][13] ;
 wire \core.registers[27][14] ;
 wire \core.registers[27][15] ;
 wire \core.registers[27][16] ;
 wire \core.registers[27][17] ;
 wire \core.registers[27][18] ;
 wire \core.registers[27][19] ;
 wire \core.registers[27][1] ;
 wire \core.registers[27][20] ;
 wire \core.registers[27][21] ;
 wire \core.registers[27][22] ;
 wire \core.registers[27][23] ;
 wire \core.registers[27][24] ;
 wire \core.registers[27][25] ;
 wire \core.registers[27][26] ;
 wire \core.registers[27][27] ;
 wire \core.registers[27][28] ;
 wire \core.registers[27][29] ;
 wire \core.registers[27][2] ;
 wire \core.registers[27][30] ;
 wire \core.registers[27][31] ;
 wire \core.registers[27][3] ;
 wire \core.registers[27][4] ;
 wire \core.registers[27][5] ;
 wire \core.registers[27][6] ;
 wire \core.registers[27][7] ;
 wire \core.registers[27][8] ;
 wire \core.registers[27][9] ;
 wire \core.registers[28][0] ;
 wire \core.registers[28][10] ;
 wire \core.registers[28][11] ;
 wire \core.registers[28][12] ;
 wire \core.registers[28][13] ;
 wire \core.registers[28][14] ;
 wire \core.registers[28][15] ;
 wire \core.registers[28][16] ;
 wire \core.registers[28][17] ;
 wire \core.registers[28][18] ;
 wire \core.registers[28][19] ;
 wire \core.registers[28][1] ;
 wire \core.registers[28][20] ;
 wire \core.registers[28][21] ;
 wire \core.registers[28][22] ;
 wire \core.registers[28][23] ;
 wire \core.registers[28][24] ;
 wire \core.registers[28][25] ;
 wire \core.registers[28][26] ;
 wire \core.registers[28][27] ;
 wire \core.registers[28][28] ;
 wire \core.registers[28][29] ;
 wire \core.registers[28][2] ;
 wire \core.registers[28][30] ;
 wire \core.registers[28][31] ;
 wire \core.registers[28][3] ;
 wire \core.registers[28][4] ;
 wire \core.registers[28][5] ;
 wire \core.registers[28][6] ;
 wire \core.registers[28][7] ;
 wire \core.registers[28][8] ;
 wire \core.registers[28][9] ;
 wire \core.registers[29][0] ;
 wire \core.registers[29][10] ;
 wire \core.registers[29][11] ;
 wire \core.registers[29][12] ;
 wire \core.registers[29][13] ;
 wire \core.registers[29][14] ;
 wire \core.registers[29][15] ;
 wire \core.registers[29][16] ;
 wire \core.registers[29][17] ;
 wire \core.registers[29][18] ;
 wire \core.registers[29][19] ;
 wire \core.registers[29][1] ;
 wire \core.registers[29][20] ;
 wire \core.registers[29][21] ;
 wire \core.registers[29][22] ;
 wire \core.registers[29][23] ;
 wire \core.registers[29][24] ;
 wire \core.registers[29][25] ;
 wire \core.registers[29][26] ;
 wire \core.registers[29][27] ;
 wire \core.registers[29][28] ;
 wire \core.registers[29][29] ;
 wire \core.registers[29][2] ;
 wire \core.registers[29][30] ;
 wire \core.registers[29][31] ;
 wire \core.registers[29][3] ;
 wire \core.registers[29][4] ;
 wire \core.registers[29][5] ;
 wire \core.registers[29][6] ;
 wire \core.registers[29][7] ;
 wire \core.registers[29][8] ;
 wire \core.registers[29][9] ;
 wire \core.registers[2][0] ;
 wire \core.registers[2][10] ;
 wire \core.registers[2][11] ;
 wire \core.registers[2][12] ;
 wire \core.registers[2][13] ;
 wire \core.registers[2][14] ;
 wire \core.registers[2][15] ;
 wire \core.registers[2][16] ;
 wire \core.registers[2][17] ;
 wire \core.registers[2][18] ;
 wire \core.registers[2][19] ;
 wire \core.registers[2][1] ;
 wire \core.registers[2][20] ;
 wire \core.registers[2][21] ;
 wire \core.registers[2][22] ;
 wire \core.registers[2][23] ;
 wire \core.registers[2][24] ;
 wire \core.registers[2][25] ;
 wire \core.registers[2][26] ;
 wire \core.registers[2][27] ;
 wire \core.registers[2][28] ;
 wire \core.registers[2][29] ;
 wire \core.registers[2][2] ;
 wire \core.registers[2][30] ;
 wire \core.registers[2][31] ;
 wire \core.registers[2][3] ;
 wire \core.registers[2][4] ;
 wire \core.registers[2][5] ;
 wire \core.registers[2][6] ;
 wire \core.registers[2][7] ;
 wire \core.registers[2][8] ;
 wire \core.registers[2][9] ;
 wire \core.registers[30][0] ;
 wire \core.registers[30][10] ;
 wire \core.registers[30][11] ;
 wire \core.registers[30][12] ;
 wire \core.registers[30][13] ;
 wire \core.registers[30][14] ;
 wire \core.registers[30][15] ;
 wire \core.registers[30][16] ;
 wire \core.registers[30][17] ;
 wire \core.registers[30][18] ;
 wire \core.registers[30][19] ;
 wire \core.registers[30][1] ;
 wire \core.registers[30][20] ;
 wire \core.registers[30][21] ;
 wire \core.registers[30][22] ;
 wire \core.registers[30][23] ;
 wire \core.registers[30][24] ;
 wire \core.registers[30][25] ;
 wire \core.registers[30][26] ;
 wire \core.registers[30][27] ;
 wire \core.registers[30][28] ;
 wire \core.registers[30][29] ;
 wire \core.registers[30][2] ;
 wire \core.registers[30][30] ;
 wire \core.registers[30][31] ;
 wire \core.registers[30][3] ;
 wire \core.registers[30][4] ;
 wire \core.registers[30][5] ;
 wire \core.registers[30][6] ;
 wire \core.registers[30][7] ;
 wire \core.registers[30][8] ;
 wire \core.registers[30][9] ;
 wire \core.registers[31][0] ;
 wire \core.registers[31][10] ;
 wire \core.registers[31][11] ;
 wire \core.registers[31][12] ;
 wire \core.registers[31][13] ;
 wire \core.registers[31][14] ;
 wire \core.registers[31][15] ;
 wire \core.registers[31][16] ;
 wire \core.registers[31][17] ;
 wire \core.registers[31][18] ;
 wire \core.registers[31][19] ;
 wire \core.registers[31][1] ;
 wire \core.registers[31][20] ;
 wire \core.registers[31][21] ;
 wire \core.registers[31][22] ;
 wire \core.registers[31][23] ;
 wire \core.registers[31][24] ;
 wire \core.registers[31][25] ;
 wire \core.registers[31][26] ;
 wire \core.registers[31][27] ;
 wire \core.registers[31][28] ;
 wire \core.registers[31][29] ;
 wire \core.registers[31][2] ;
 wire \core.registers[31][30] ;
 wire \core.registers[31][31] ;
 wire \core.registers[31][3] ;
 wire \core.registers[31][4] ;
 wire \core.registers[31][5] ;
 wire \core.registers[31][6] ;
 wire \core.registers[31][7] ;
 wire \core.registers[31][8] ;
 wire \core.registers[31][9] ;
 wire \core.registers[3][0] ;
 wire \core.registers[3][10] ;
 wire \core.registers[3][11] ;
 wire \core.registers[3][12] ;
 wire \core.registers[3][13] ;
 wire \core.registers[3][14] ;
 wire \core.registers[3][15] ;
 wire \core.registers[3][16] ;
 wire \core.registers[3][17] ;
 wire \core.registers[3][18] ;
 wire \core.registers[3][19] ;
 wire \core.registers[3][1] ;
 wire \core.registers[3][20] ;
 wire \core.registers[3][21] ;
 wire \core.registers[3][22] ;
 wire \core.registers[3][23] ;
 wire \core.registers[3][24] ;
 wire \core.registers[3][25] ;
 wire \core.registers[3][26] ;
 wire \core.registers[3][27] ;
 wire \core.registers[3][28] ;
 wire \core.registers[3][29] ;
 wire \core.registers[3][2] ;
 wire \core.registers[3][30] ;
 wire \core.registers[3][31] ;
 wire \core.registers[3][3] ;
 wire \core.registers[3][4] ;
 wire \core.registers[3][5] ;
 wire \core.registers[3][6] ;
 wire \core.registers[3][7] ;
 wire \core.registers[3][8] ;
 wire \core.registers[3][9] ;
 wire \core.registers[4][0] ;
 wire \core.registers[4][10] ;
 wire \core.registers[4][11] ;
 wire \core.registers[4][12] ;
 wire \core.registers[4][13] ;
 wire \core.registers[4][14] ;
 wire \core.registers[4][15] ;
 wire \core.registers[4][16] ;
 wire \core.registers[4][17] ;
 wire \core.registers[4][18] ;
 wire \core.registers[4][19] ;
 wire \core.registers[4][1] ;
 wire \core.registers[4][20] ;
 wire \core.registers[4][21] ;
 wire \core.registers[4][22] ;
 wire \core.registers[4][23] ;
 wire \core.registers[4][24] ;
 wire \core.registers[4][25] ;
 wire \core.registers[4][26] ;
 wire \core.registers[4][27] ;
 wire \core.registers[4][28] ;
 wire \core.registers[4][29] ;
 wire \core.registers[4][2] ;
 wire \core.registers[4][30] ;
 wire \core.registers[4][31] ;
 wire \core.registers[4][3] ;
 wire \core.registers[4][4] ;
 wire \core.registers[4][5] ;
 wire \core.registers[4][6] ;
 wire \core.registers[4][7] ;
 wire \core.registers[4][8] ;
 wire \core.registers[4][9] ;
 wire \core.registers[5][0] ;
 wire \core.registers[5][10] ;
 wire \core.registers[5][11] ;
 wire \core.registers[5][12] ;
 wire \core.registers[5][13] ;
 wire \core.registers[5][14] ;
 wire \core.registers[5][15] ;
 wire \core.registers[5][16] ;
 wire \core.registers[5][17] ;
 wire \core.registers[5][18] ;
 wire \core.registers[5][19] ;
 wire \core.registers[5][1] ;
 wire \core.registers[5][20] ;
 wire \core.registers[5][21] ;
 wire \core.registers[5][22] ;
 wire \core.registers[5][23] ;
 wire \core.registers[5][24] ;
 wire \core.registers[5][25] ;
 wire \core.registers[5][26] ;
 wire \core.registers[5][27] ;
 wire \core.registers[5][28] ;
 wire \core.registers[5][29] ;
 wire \core.registers[5][2] ;
 wire \core.registers[5][30] ;
 wire \core.registers[5][31] ;
 wire \core.registers[5][3] ;
 wire \core.registers[5][4] ;
 wire \core.registers[5][5] ;
 wire \core.registers[5][6] ;
 wire \core.registers[5][7] ;
 wire \core.registers[5][8] ;
 wire \core.registers[5][9] ;
 wire \core.registers[6][0] ;
 wire \core.registers[6][10] ;
 wire \core.registers[6][11] ;
 wire \core.registers[6][12] ;
 wire \core.registers[6][13] ;
 wire \core.registers[6][14] ;
 wire \core.registers[6][15] ;
 wire \core.registers[6][16] ;
 wire \core.registers[6][17] ;
 wire \core.registers[6][18] ;
 wire \core.registers[6][19] ;
 wire \core.registers[6][1] ;
 wire \core.registers[6][20] ;
 wire \core.registers[6][21] ;
 wire \core.registers[6][22] ;
 wire \core.registers[6][23] ;
 wire \core.registers[6][24] ;
 wire \core.registers[6][25] ;
 wire \core.registers[6][26] ;
 wire \core.registers[6][27] ;
 wire \core.registers[6][28] ;
 wire \core.registers[6][29] ;
 wire \core.registers[6][2] ;
 wire \core.registers[6][30] ;
 wire \core.registers[6][31] ;
 wire \core.registers[6][3] ;
 wire \core.registers[6][4] ;
 wire \core.registers[6][5] ;
 wire \core.registers[6][6] ;
 wire \core.registers[6][7] ;
 wire \core.registers[6][8] ;
 wire \core.registers[6][9] ;
 wire \core.registers[7][0] ;
 wire \core.registers[7][10] ;
 wire \core.registers[7][11] ;
 wire \core.registers[7][12] ;
 wire \core.registers[7][13] ;
 wire \core.registers[7][14] ;
 wire \core.registers[7][15] ;
 wire \core.registers[7][16] ;
 wire \core.registers[7][17] ;
 wire \core.registers[7][18] ;
 wire \core.registers[7][19] ;
 wire \core.registers[7][1] ;
 wire \core.registers[7][20] ;
 wire \core.registers[7][21] ;
 wire \core.registers[7][22] ;
 wire \core.registers[7][23] ;
 wire \core.registers[7][24] ;
 wire \core.registers[7][25] ;
 wire \core.registers[7][26] ;
 wire \core.registers[7][27] ;
 wire \core.registers[7][28] ;
 wire \core.registers[7][29] ;
 wire \core.registers[7][2] ;
 wire \core.registers[7][30] ;
 wire \core.registers[7][31] ;
 wire \core.registers[7][3] ;
 wire \core.registers[7][4] ;
 wire \core.registers[7][5] ;
 wire \core.registers[7][6] ;
 wire \core.registers[7][7] ;
 wire \core.registers[7][8] ;
 wire \core.registers[7][9] ;
 wire \core.registers[8][0] ;
 wire \core.registers[8][10] ;
 wire \core.registers[8][11] ;
 wire \core.registers[8][12] ;
 wire \core.registers[8][13] ;
 wire \core.registers[8][14] ;
 wire \core.registers[8][15] ;
 wire \core.registers[8][16] ;
 wire \core.registers[8][17] ;
 wire \core.registers[8][18] ;
 wire \core.registers[8][19] ;
 wire \core.registers[8][1] ;
 wire \core.registers[8][20] ;
 wire \core.registers[8][21] ;
 wire \core.registers[8][22] ;
 wire \core.registers[8][23] ;
 wire \core.registers[8][24] ;
 wire \core.registers[8][25] ;
 wire \core.registers[8][26] ;
 wire \core.registers[8][27] ;
 wire \core.registers[8][28] ;
 wire \core.registers[8][29] ;
 wire \core.registers[8][2] ;
 wire \core.registers[8][30] ;
 wire \core.registers[8][31] ;
 wire \core.registers[8][3] ;
 wire \core.registers[8][4] ;
 wire \core.registers[8][5] ;
 wire \core.registers[8][6] ;
 wire \core.registers[8][7] ;
 wire \core.registers[8][8] ;
 wire \core.registers[8][9] ;
 wire \core.registers[9][0] ;
 wire \core.registers[9][10] ;
 wire \core.registers[9][11] ;
 wire \core.registers[9][12] ;
 wire \core.registers[9][13] ;
 wire \core.registers[9][14] ;
 wire \core.registers[9][15] ;
 wire \core.registers[9][16] ;
 wire \core.registers[9][17] ;
 wire \core.registers[9][18] ;
 wire \core.registers[9][19] ;
 wire \core.registers[9][1] ;
 wire \core.registers[9][20] ;
 wire \core.registers[9][21] ;
 wire \core.registers[9][22] ;
 wire \core.registers[9][23] ;
 wire \core.registers[9][24] ;
 wire \core.registers[9][25] ;
 wire \core.registers[9][26] ;
 wire \core.registers[9][27] ;
 wire \core.registers[9][28] ;
 wire \core.registers[9][29] ;
 wire \core.registers[9][2] ;
 wire \core.registers[9][30] ;
 wire \core.registers[9][31] ;
 wire \core.registers[9][3] ;
 wire \core.registers[9][4] ;
 wire \core.registers[9][5] ;
 wire \core.registers[9][6] ;
 wire \core.registers[9][7] ;
 wire \core.registers[9][8] ;
 wire \core.registers[9][9] ;
 wire \core.useCachedLoad ;
 wire \coreManagement.control[1] ;
 wire \coreWBInterface.readDataBuffered[0] ;
 wire \coreWBInterface.readDataBuffered[10] ;
 wire \coreWBInterface.readDataBuffered[11] ;
 wire \coreWBInterface.readDataBuffered[12] ;
 wire \coreWBInterface.readDataBuffered[13] ;
 wire \coreWBInterface.readDataBuffered[14] ;
 wire \coreWBInterface.readDataBuffered[15] ;
 wire \coreWBInterface.readDataBuffered[16] ;
 wire \coreWBInterface.readDataBuffered[17] ;
 wire \coreWBInterface.readDataBuffered[18] ;
 wire \coreWBInterface.readDataBuffered[19] ;
 wire \coreWBInterface.readDataBuffered[1] ;
 wire \coreWBInterface.readDataBuffered[20] ;
 wire \coreWBInterface.readDataBuffered[21] ;
 wire \coreWBInterface.readDataBuffered[22] ;
 wire \coreWBInterface.readDataBuffered[23] ;
 wire \coreWBInterface.readDataBuffered[24] ;
 wire \coreWBInterface.readDataBuffered[25] ;
 wire \coreWBInterface.readDataBuffered[26] ;
 wire \coreWBInterface.readDataBuffered[27] ;
 wire \coreWBInterface.readDataBuffered[28] ;
 wire \coreWBInterface.readDataBuffered[29] ;
 wire \coreWBInterface.readDataBuffered[2] ;
 wire \coreWBInterface.readDataBuffered[30] ;
 wire \coreWBInterface.readDataBuffered[31] ;
 wire \coreWBInterface.readDataBuffered[3] ;
 wire \coreWBInterface.readDataBuffered[4] ;
 wire \coreWBInterface.readDataBuffered[5] ;
 wire \coreWBInterface.readDataBuffered[6] ;
 wire \coreWBInterface.readDataBuffered[7] ;
 wire \coreWBInterface.readDataBuffered[8] ;
 wire \coreWBInterface.readDataBuffered[9] ;
 wire \coreWBInterface.state[0] ;
 wire \coreWBInterface.state[1] ;
 wire \coreWBInterface.stb ;
 wire \jtag.dataBSRRegister.data[0] ;
 wire \jtag.dataBSRRegister.data[10] ;
 wire \jtag.dataBSRRegister.data[11] ;
 wire \jtag.dataBSRRegister.data[12] ;
 wire \jtag.dataBSRRegister.data[13] ;
 wire \jtag.dataBSRRegister.data[14] ;
 wire \jtag.dataBSRRegister.data[15] ;
 wire \jtag.dataBSRRegister.data[16] ;
 wire \jtag.dataBSRRegister.data[17] ;
 wire \jtag.dataBSRRegister.data[18] ;
 wire \jtag.dataBSRRegister.data[19] ;
 wire \jtag.dataBSRRegister.data[1] ;
 wire \jtag.dataBSRRegister.data[20] ;
 wire \jtag.dataBSRRegister.data[21] ;
 wire \jtag.dataBSRRegister.data[22] ;
 wire \jtag.dataBSRRegister.data[23] ;
 wire \jtag.dataBSRRegister.data[24] ;
 wire \jtag.dataBSRRegister.data[25] ;
 wire \jtag.dataBSRRegister.data[26] ;
 wire \jtag.dataBSRRegister.data[27] ;
 wire \jtag.dataBSRRegister.data[28] ;
 wire \jtag.dataBSRRegister.data[29] ;
 wire \jtag.dataBSRRegister.data[2] ;
 wire \jtag.dataBSRRegister.data[30] ;
 wire \jtag.dataBSRRegister.data[31] ;
 wire \jtag.dataBSRRegister.data[3] ;
 wire \jtag.dataBSRRegister.data[4] ;
 wire \jtag.dataBSRRegister.data[5] ;
 wire \jtag.dataBSRRegister.data[6] ;
 wire \jtag.dataBSRRegister.data[7] ;
 wire \jtag.dataBSRRegister.data[8] ;
 wire \jtag.dataBSRRegister.data[9] ;
 wire \jtag.dataBypassRegister.data ;
 wire \jtag.dataIDRegister.data[0] ;
 wire \jtag.dataIDRegister.data[10] ;
 wire \jtag.dataIDRegister.data[11] ;
 wire \jtag.dataIDRegister.data[12] ;
 wire \jtag.dataIDRegister.data[13] ;
 wire \jtag.dataIDRegister.data[14] ;
 wire \jtag.dataIDRegister.data[15] ;
 wire \jtag.dataIDRegister.data[16] ;
 wire \jtag.dataIDRegister.data[17] ;
 wire \jtag.dataIDRegister.data[18] ;
 wire \jtag.dataIDRegister.data[19] ;
 wire \jtag.dataIDRegister.data[1] ;
 wire \jtag.dataIDRegister.data[20] ;
 wire \jtag.dataIDRegister.data[21] ;
 wire \jtag.dataIDRegister.data[22] ;
 wire \jtag.dataIDRegister.data[23] ;
 wire \jtag.dataIDRegister.data[24] ;
 wire \jtag.dataIDRegister.data[25] ;
 wire \jtag.dataIDRegister.data[26] ;
 wire \jtag.dataIDRegister.data[27] ;
 wire \jtag.dataIDRegister.data[28] ;
 wire \jtag.dataIDRegister.data[29] ;
 wire \jtag.dataIDRegister.data[2] ;
 wire \jtag.dataIDRegister.data[30] ;
 wire \jtag.dataIDRegister.data[31] ;
 wire \jtag.dataIDRegister.data[3] ;
 wire \jtag.dataIDRegister.data[4] ;
 wire \jtag.dataIDRegister.data[5] ;
 wire \jtag.dataIDRegister.data[6] ;
 wire \jtag.dataIDRegister.data[7] ;
 wire \jtag.dataIDRegister.data[8] ;
 wire \jtag.dataIDRegister.data[9] ;
 wire \jtag.instructionRegister.data[0] ;
 wire \jtag.instructionRegister.data[1] ;
 wire \jtag.instructionRegister.data[2] ;
 wire \jtag.instructionRegister.data[3] ;
 wire \jtag.instructionRegister.data[4] ;
 wire \jtag.managementAddress[0] ;
 wire \jtag.managementAddress[10] ;
 wire \jtag.managementAddress[11] ;
 wire \jtag.managementAddress[12] ;
 wire \jtag.managementAddress[13] ;
 wire \jtag.managementAddress[14] ;
 wire \jtag.managementAddress[15] ;
 wire \jtag.managementAddress[16] ;
 wire \jtag.managementAddress[17] ;
 wire \jtag.managementAddress[18] ;
 wire \jtag.managementAddress[19] ;
 wire \jtag.managementAddress[1] ;
 wire \jtag.managementAddress[2] ;
 wire \jtag.managementAddress[3] ;
 wire \jtag.managementAddress[4] ;
 wire \jtag.managementAddress[5] ;
 wire \jtag.managementAddress[6] ;
 wire \jtag.managementAddress[7] ;
 wire \jtag.managementAddress[8] ;
 wire \jtag.managementAddress[9] ;
 wire \jtag.managementReadData[0] ;
 wire \jtag.managementReadData[10] ;
 wire \jtag.managementReadData[11] ;
 wire \jtag.managementReadData[12] ;
 wire \jtag.managementReadData[13] ;
 wire \jtag.managementReadData[14] ;
 wire \jtag.managementReadData[15] ;
 wire \jtag.managementReadData[16] ;
 wire \jtag.managementReadData[17] ;
 wire \jtag.managementReadData[18] ;
 wire \jtag.managementReadData[19] ;
 wire \jtag.managementReadData[1] ;
 wire \jtag.managementReadData[20] ;
 wire \jtag.managementReadData[21] ;
 wire \jtag.managementReadData[22] ;
 wire \jtag.managementReadData[23] ;
 wire \jtag.managementReadData[24] ;
 wire \jtag.managementReadData[25] ;
 wire \jtag.managementReadData[26] ;
 wire \jtag.managementReadData[27] ;
 wire \jtag.managementReadData[28] ;
 wire \jtag.managementReadData[29] ;
 wire \jtag.managementReadData[2] ;
 wire \jtag.managementReadData[30] ;
 wire \jtag.managementReadData[31] ;
 wire \jtag.managementReadData[3] ;
 wire \jtag.managementReadData[4] ;
 wire \jtag.managementReadData[5] ;
 wire \jtag.managementReadData[6] ;
 wire \jtag.managementReadData[7] ;
 wire \jtag.managementReadData[8] ;
 wire \jtag.managementReadData[9] ;
 wire \jtag.managementState[0] ;
 wire \jtag.managementState[1] ;
 wire \jtag.managementState[2] ;
 wire \jtag.state[0] ;
 wire \jtag.state[1] ;
 wire \jtag.state[2] ;
 wire \jtag.state[3] ;
 wire \jtag.tckRisingEdge ;
 wire \jtag.tckState ;
 wire \localMemoryInterface.coreReadReady ;
 wire \localMemoryInterface.lastCoreByteSelect[0] ;
 wire \localMemoryInterface.lastCoreByteSelect[1] ;
 wire \localMemoryInterface.lastCoreByteSelect[2] ;
 wire \localMemoryInterface.lastCoreByteSelect[3] ;
 wire \localMemoryInterface.lastRBankSelect ;
 wire \localMemoryInterface.lastRWBankSelect ;
 wire \localMemoryInterface.lastWBByteSelect[0] ;
 wire \localMemoryInterface.lastWBByteSelect[1] ;
 wire \localMemoryInterface.lastWBByteSelect[2] ;
 wire \localMemoryInterface.lastWBByteSelect[3] ;
 wire \localMemoryInterface.wbReadReady ;
 wire \memoryController.last_data_enableLocalMemory ;
 wire \memoryController.last_data_enableWB ;
 wire \memoryController.last_instruction_enableLocalMemory ;
 wire \memoryController.last_instruction_enableWB ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \wbSRAMInterface.currentAddress[0] ;
 wire \wbSRAMInterface.currentAddress[10] ;
 wire \wbSRAMInterface.currentAddress[11] ;
 wire \wbSRAMInterface.currentAddress[12] ;
 wire \wbSRAMInterface.currentAddress[13] ;
 wire \wbSRAMInterface.currentAddress[14] ;
 wire \wbSRAMInterface.currentAddress[15] ;
 wire \wbSRAMInterface.currentAddress[16] ;
 wire \wbSRAMInterface.currentAddress[17] ;
 wire \wbSRAMInterface.currentAddress[18] ;
 wire \wbSRAMInterface.currentAddress[19] ;
 wire \wbSRAMInterface.currentAddress[1] ;
 wire \wbSRAMInterface.currentAddress[20] ;
 wire \wbSRAMInterface.currentAddress[21] ;
 wire \wbSRAMInterface.currentAddress[22] ;
 wire \wbSRAMInterface.currentAddress[23] ;
 wire \wbSRAMInterface.currentAddress[2] ;
 wire \wbSRAMInterface.currentAddress[3] ;
 wire \wbSRAMInterface.currentAddress[4] ;
 wire \wbSRAMInterface.currentAddress[5] ;
 wire \wbSRAMInterface.currentAddress[6] ;
 wire \wbSRAMInterface.currentAddress[7] ;
 wire \wbSRAMInterface.currentAddress[8] ;
 wire \wbSRAMInterface.currentAddress[9] ;
 wire \wbSRAMInterface.currentByteSelect[0] ;
 wire \wbSRAMInterface.currentByteSelect[1] ;
 wire \wbSRAMInterface.currentByteSelect[2] ;
 wire \wbSRAMInterface.currentByteSelect[3] ;
 wire \wbSRAMInterface.state[0] ;
 wire \wbSRAMInterface.state[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_07346_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_07378_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_07394_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_07399_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_07492_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_07874_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_07886_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_08345_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_08379_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_08379_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_02246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_08402_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_08407_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_08437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_08437_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_08495_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_08506_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_08506_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_08509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_08509_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_08510_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_08510_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_08513_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_08513_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_08514_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(_08515_));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_08520_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(_08520_));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_08523_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(_08523_));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(_08523_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_08529_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_08533_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_08541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_08541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_08541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(_08541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(_08541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(_08544_));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(_08563_));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(_08574_));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(_08577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_08577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_08584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_08594_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_08594_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_08598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_08602_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_08610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_08610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_08614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_08618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_08618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_08618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(_08618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(_08618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(_08618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_08618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_08623_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_08636_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(_08650_));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(_08650_));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(_09110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(\core.csr.currentInstruction[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(\core.csr.currentInstruction[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(\core.csr.currentInstruction[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(\core.csr.currentInstruction[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(\core.csr.currentInstruction[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(\core.csr.currentInstruction[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(\core.csr.currentInstruction[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(\core.csr.currentInstruction[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(\core.csr.currentInstruction[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(\core.csr.currentInstruction[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(\core.csr.currentInstruction[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(\core.csr.currentInstruction[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(\core.csr.currentInstruction[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(\core.fetchProgramCounter[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(\core.pipe0_currentInstruction[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(\core.pipe0_currentInstruction[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(\core.pipe0_currentInstruction[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(\core.pipe0_currentInstruction[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(\core.pipe0_currentInstruction[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(\core.pipe0_currentInstruction[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(\core.pipe0_currentInstruction[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(\core.pipe0_currentInstruction[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(\core.pipe0_currentInstruction[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_02346_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(\core.pipe0_currentInstruction[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(\core.pipe0_currentInstruction[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(\core.pipe1_resultRegister[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(\core.pipe1_resultRegister[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(\core.pipe1_resultRegister[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(\core.pipe1_resultRegister[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(\core.pipe1_resultRegister[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(\core.pipe1_resultRegister[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(\core.pipe1_resultRegister[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(\core.registers[0][23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00572_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(\core.registers[0][27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(\coreWBInterface.readDataBuffered[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(\coreWBInterface.readDataBuffered[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(\coreWBInterface.readDataBuffered[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(\coreWBInterface.readDataBuffered[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(\coreWBInterface.readDataBuffered[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(\jtag.dataIDRegister.data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_02415_));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_02478_));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(\wbSRAMInterface.currentAddress[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(\wbSRAMInterface.currentAddress[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(\wbSRAMInterface.currentByteSelect[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_02609_));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(\wbSRAMInterface.currentByteSelect[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(\wbSRAMInterface.currentByteSelect[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00574_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_02688_));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(net1473));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(net1746));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(net1746));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(net1776));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(net1815));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(net1819));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(net1831));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(net1831));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(net1852));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(net1852));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_03119_));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(net1852));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(net1852));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(net1852));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(net1852));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(net1867));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(net1867));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(net1871));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(net1871));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(_02037_));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(_02100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(_02269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_03129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(_02415_));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(_02451_));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(_02469_));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(_02609_));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(_02687_));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(_02759_));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(_02795_));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_02058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_03139_));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(_03283_));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(_03290_));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(_03311_));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(_03348_));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(_03362_));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(_03593_));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_03194_));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(_03794_));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(_03802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(_03802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_414 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA_415 (.DIODE(_03806_));
 sky130_fd_sc_hd__diode_2 ANTENNA_416 (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA_417 (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA_418 (.DIODE(_04128_));
 sky130_fd_sc_hd__diode_2 ANTENNA_419 (.DIODE(_04537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA_420 (.DIODE(_04641_));
 sky130_fd_sc_hd__diode_2 ANTENNA_421 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_422 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA_423 (.DIODE(_05292_));
 sky130_fd_sc_hd__diode_2 ANTENNA_424 (.DIODE(_05375_));
 sky130_fd_sc_hd__diode_2 ANTENNA_425 (.DIODE(_05726_));
 sky130_fd_sc_hd__diode_2 ANTENNA_426 (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA_427 (.DIODE(_07241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_428 (.DIODE(_07273_));
 sky130_fd_sc_hd__diode_2 ANTENNA_429 (.DIODE(_07865_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_03227_));
 sky130_fd_sc_hd__diode_2 ANTENNA_430 (.DIODE(_08052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_431 (.DIODE(_08508_));
 sky130_fd_sc_hd__diode_2 ANTENNA_432 (.DIODE(_08512_));
 sky130_fd_sc_hd__diode_2 ANTENNA_433 (.DIODE(_08525_));
 sky130_fd_sc_hd__diode_2 ANTENNA_434 (.DIODE(_08529_));
 sky130_fd_sc_hd__diode_2 ANTENNA_435 (.DIODE(_08551_));
 sky130_fd_sc_hd__diode_2 ANTENNA_436 (.DIODE(_08566_));
 sky130_fd_sc_hd__diode_2 ANTENNA_437 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_438 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_439 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA_440 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_441 (.DIODE(_08571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_442 (.DIODE(_08574_));
 sky130_fd_sc_hd__diode_2 ANTENNA_443 (.DIODE(_08574_));
 sky130_fd_sc_hd__diode_2 ANTENNA_444 (.DIODE(_08598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_445 (.DIODE(_08598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_446 (.DIODE(_08598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_447 (.DIODE(_08598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_448 (.DIODE(_08610_));
 sky130_fd_sc_hd__diode_2 ANTENNA_449 (.DIODE(_08614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_03234_));
 sky130_fd_sc_hd__diode_2 ANTENNA_450 (.DIODE(_08614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_451 (.DIODE(_08614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_452 (.DIODE(_08650_));
 sky130_fd_sc_hd__diode_2 ANTENNA_453 (.DIODE(\core.csr.currentInstruction[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_454 (.DIODE(\core.csr.currentInstruction[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_455 (.DIODE(\core.csr.currentInstruction[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_456 (.DIODE(\core.csr.currentInstruction[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_457 (.DIODE(\core.csr.currentInstruction[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_458 (.DIODE(\core.csr.currentInstruction[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_459 (.DIODE(\core.csr.currentInstruction[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA_460 (.DIODE(\core.fetchProgramCounter[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_461 (.DIODE(\core.fetchProgramCounter[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_462 (.DIODE(\core.fetchProgramCounter[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_463 (.DIODE(\core.pipe0_currentInstruction[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_464 (.DIODE(\coreWBInterface.readDataBuffered[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_465 (.DIODE(\coreWBInterface.readDataBuffered[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_466 (.DIODE(\coreWBInterface.readDataBuffered[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_467 (.DIODE(\coreWBInterface.readDataBuffered[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_468 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_469 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA_470 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_471 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_472 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_473 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_474 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_475 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_476 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_477 (.DIODE(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_478 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_479 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_03261_));
 sky130_fd_sc_hd__diode_2 ANTENNA_480 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_481 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_482 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_483 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_484 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_485 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_486 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_487 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_488 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_489 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_03269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_490 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_491 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_492 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_493 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_494 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_495 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_496 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_497 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_498 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_499 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_02093_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_03297_));
 sky130_fd_sc_hd__diode_2 ANTENNA_500 (.DIODE(\wbSRAMInterface.currentAddress[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_501 (.DIODE(\wbSRAMInterface.currentByteSelect[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_502 (.DIODE(\wbSRAMInterface.currentByteSelect[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_503 (.DIODE(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_504 (.DIODE(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_505 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_506 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_507 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_508 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_509 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_03304_));
 sky130_fd_sc_hd__diode_2 ANTENNA_510 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_511 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_512 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_513 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_514 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_515 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_516 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_517 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_518 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_519 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_03320_));
 sky130_fd_sc_hd__diode_2 ANTENNA_520 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_521 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_522 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_523 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_524 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_525 (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_526 (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_527 (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA_528 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_529 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_03327_));
 sky130_fd_sc_hd__diode_2 ANTENNA_530 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_531 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_532 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_533 (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_534 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_535 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA_536 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_537 (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA_538 (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA_539 (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_03334_));
 sky130_fd_sc_hd__diode_2 ANTENNA_540 (.DIODE(net1477));
 sky130_fd_sc_hd__diode_2 ANTENNA_541 (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA_542 (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA_543 (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA_544 (.DIODE(net1714));
 sky130_fd_sc_hd__diode_2 ANTENNA_545 (.DIODE(net1829));
 sky130_fd_sc_hd__diode_2 ANTENNA_546 (.DIODE(net1852));
 sky130_fd_sc_hd__diode_2 ANTENNA_547 (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_548 (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_549 (.DIODE(_02100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_03341_));
 sky130_fd_sc_hd__diode_2 ANTENNA_550 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_551 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_552 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_553 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_554 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_555 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_556 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_557 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_558 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_559 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_03355_));
 sky130_fd_sc_hd__diode_2 ANTENNA_560 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_561 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_562 (.DIODE(_02240_));
 sky130_fd_sc_hd__diode_2 ANTENNA_563 (.DIODE(_02384_));
 sky130_fd_sc_hd__diode_2 ANTENNA_564 (.DIODE(_06112_));
 sky130_fd_sc_hd__diode_2 ANTENNA_565 (.DIODE(_08376_));
 sky130_fd_sc_hd__diode_2 ANTENNA_566 (.DIODE(_08376_));
 sky130_fd_sc_hd__diode_2 ANTENNA_567 (.DIODE(_08512_));
 sky130_fd_sc_hd__diode_2 ANTENNA_568 (.DIODE(_08566_));
 sky130_fd_sc_hd__diode_2 ANTENNA_569 (.DIODE(_08618_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_03363_));
 sky130_fd_sc_hd__diode_2 ANTENNA_570 (.DIODE(\core.csr.currentInstruction[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_571 (.DIODE(\coreWBInterface.readDataBuffered[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_572 (.DIODE(\coreWBInterface.readDataBuffered[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_573 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_574 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_575 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_576 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_577 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_578 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_579 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA_580 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_581 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_582 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_583 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_584 (.DIODE(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_585 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_586 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_587 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_588 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_589 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA_590 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_591 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_592 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_593 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_594 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_595 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_596 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_597 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_598 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_599 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_02157_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA_600 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_601 (.DIODE(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_602 (.DIODE(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_603 (.DIODE(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_604 (.DIODE(\wbSRAMInterface.currentByteSelect[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_605 (.DIODE(\wbSRAMInterface.currentByteSelect[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_606 (.DIODE(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_607 (.DIODE(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_608 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_609 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_03608_));
 sky130_fd_sc_hd__diode_2 ANTENNA_610 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_611 (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA_612 (.DIODE(net1666));
 sky130_fd_sc_hd__diode_2 ANTENNA_613 (.DIODE(net1666));
 sky130_fd_sc_hd__diode_2 ANTENNA_614 (.DIODE(_08614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_615 (.DIODE(_08614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_616 (.DIODE(_08614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_617 (.DIODE(_08614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_618 (.DIODE(_08614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_619 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA_620 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_621 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_622 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_623 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_624 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_625 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_626 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_627 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_628 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_629 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_03786_));
 sky130_fd_sc_hd__diode_2 ANTENNA_630 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_631 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_632 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_633 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_634 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_635 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_636 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_637 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_638 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_639 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_03810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_640 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_641 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_642 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_643 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_644 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_645 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_646 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_647 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_648 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_649 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_03810_));
 sky130_fd_sc_hd__diode_2 ANTENNA_650 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_651 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_652 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_653 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_654 (.DIODE(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_655 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_03882_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_03890_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_04295_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_04415_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_02212_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_04560_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_04663_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_04782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_04859_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_05627_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_06365_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_06445_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_06481_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_06600_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_02234_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_06720_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_06945_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_06953_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_07067_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_07190_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_07315_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_07315_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_07346_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_07346_));
 sky130_fd_sc_hd__conb_1 ExperiarCore_2007 (.LO(net2007));
 sky130_fd_sc_hd__decap_6 FILLER_0_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_997 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _09477_ (.A(net1883),
    .Y(_04391_));
 sky130_fd_sc_hd__inv_2 _09478_ (.A(\core.csr.traps.mtval.csrReadData[1] ),
    .Y(_04392_));
 sky130_fd_sc_hd__inv_2 _09479_ (.A(\core.csr.traps.mtvec.csrReadData[6] ),
    .Y(_04393_));
 sky130_fd_sc_hd__inv_2 _09480_ (.A(\core.csr.traps.mtvec.csrReadData[2] ),
    .Y(_04394_));
 sky130_fd_sc_hd__inv_2 _09481_ (.A(\core.csr.traps.mcause.csrReadData[0] ),
    .Y(_04395_));
 sky130_fd_sc_hd__inv_2 _09482_ (.A(\core.csr.mconfigptr.currentValue[8] ),
    .Y(_04396_));
 sky130_fd_sc_hd__inv_2 _09483_ (.A(\jtag.managementState[0] ),
    .Y(_04397_));
 sky130_fd_sc_hd__clkinv_4 _09484_ (.A(net1781),
    .Y(_04398_));
 sky130_fd_sc_hd__inv_2 _09485_ (.A(net1780),
    .Y(_04399_));
 sky130_fd_sc_hd__inv_2 _09486_ (.A(net409),
    .Y(_04400_));
 sky130_fd_sc_hd__inv_4 _09487_ (.A(net1806),
    .Y(_04401_));
 sky130_fd_sc_hd__inv_4 _09488_ (.A(net1767),
    .Y(_04402_));
 sky130_fd_sc_hd__inv_2 _09489_ (.A(net474),
    .Y(_04403_));
 sky130_fd_sc_hd__inv_2 _09490_ (.A(\core.csr.instruction_memoryAddress[29] ),
    .Y(_04404_));
 sky130_fd_sc_hd__inv_2 _09491_ (.A(\core.csr.instruction_memoryAddress[22] ),
    .Y(_04405_));
 sky130_fd_sc_hd__clkinv_2 _09492_ (.A(net479),
    .Y(_04406_));
 sky130_fd_sc_hd__inv_2 _09493_ (.A(\core.csr.instruction_memoryAddress[5] ),
    .Y(_04407_));
 sky130_fd_sc_hd__inv_2 _09494_ (.A(\core.csr.instruction_memoryAddress[4] ),
    .Y(_04408_));
 sky130_fd_sc_hd__inv_2 _09495_ (.A(net1813),
    .Y(_04409_));
 sky130_fd_sc_hd__inv_2 _09496_ (.A(\core.fetchProgramCounter[16] ),
    .Y(_04410_));
 sky130_fd_sc_hd__inv_2 _09497_ (.A(\core.fetchProgramCounter[11] ),
    .Y(_04411_));
 sky130_fd_sc_hd__inv_2 _09498_ (.A(\core.fetchProgramCounter[1] ),
    .Y(_04412_));
 sky130_fd_sc_hd__inv_2 _09499_ (.A(\core.pipe0_fetch.instructionCached ),
    .Y(_04413_));
 sky130_fd_sc_hd__inv_6 _09500_ (.A(\core.pipe0_currentInstruction[29] ),
    .Y(_04414_));
 sky130_fd_sc_hd__inv_12 _09501_ (.A(net1828),
    .Y(_04415_));
 sky130_fd_sc_hd__inv_6 _09502_ (.A(net1834),
    .Y(_04416_));
 sky130_fd_sc_hd__inv_6 _09503_ (.A(net1845),
    .Y(_04417_));
 sky130_fd_sc_hd__clkinv_8 _09504_ (.A(net1851),
    .Y(_04418_));
 sky130_fd_sc_hd__inv_2 _09505_ (.A(net1857),
    .Y(_04419_));
 sky130_fd_sc_hd__inv_2 _09506_ (.A(net1865),
    .Y(_04420_));
 sky130_fd_sc_hd__inv_2 _09507_ (.A(net1872),
    .Y(_04421_));
 sky130_fd_sc_hd__inv_2 _09508_ (.A(\core.pipe0_currentInstruction[15] ),
    .Y(_04422_));
 sky130_fd_sc_hd__inv_8 _09509_ (.A(net1879),
    .Y(_04423_));
 sky130_fd_sc_hd__inv_2 _09510_ (.A(\core.csr.currentInstruction[9] ),
    .Y(_04424_));
 sky130_fd_sc_hd__inv_2 _09511_ (.A(\core.csr.currentInstruction[7] ),
    .Y(_04425_));
 sky130_fd_sc_hd__inv_2 _09512_ (.A(\core.csr.currentInstruction[6] ),
    .Y(_04426_));
 sky130_fd_sc_hd__inv_2 _09513_ (.A(\core.csr.currentInstruction[3] ),
    .Y(_04427_));
 sky130_fd_sc_hd__inv_2 _09514_ (.A(\core.csr.currentInstruction[2] ),
    .Y(_04428_));
 sky130_fd_sc_hd__clkinv_8 _09515_ (.A(net2001),
    .Y(_04429_));
 sky130_fd_sc_hd__inv_6 _09516_ (.A(\memoryController.last_data_enableLocalMemory ),
    .Y(_04430_));
 sky130_fd_sc_hd__inv_6 _09517_ (.A(\memoryController.last_instruction_enableLocalMemory ),
    .Y(_04431_));
 sky130_fd_sc_hd__inv_2 _09518_ (.A(net43),
    .Y(_04432_));
 sky130_fd_sc_hd__inv_2 _09519_ (.A(net54),
    .Y(_04433_));
 sky130_fd_sc_hd__inv_2 _09520_ (.A(net65),
    .Y(_04434_));
 sky130_fd_sc_hd__inv_2 _09521_ (.A(net105),
    .Y(_04435_));
 sky130_fd_sc_hd__inv_2 _09522_ (.A(net106),
    .Y(_04436_));
 sky130_fd_sc_hd__inv_2 _09523_ (.A(net44),
    .Y(_04437_));
 sky130_fd_sc_hd__inv_2 _09524_ (.A(net45),
    .Y(_04438_));
 sky130_fd_sc_hd__inv_2 _09525_ (.A(net46),
    .Y(_04439_));
 sky130_fd_sc_hd__inv_2 _09526_ (.A(net47),
    .Y(_04440_));
 sky130_fd_sc_hd__inv_2 _09527_ (.A(net48),
    .Y(_04441_));
 sky130_fd_sc_hd__inv_2 _09528_ (.A(net49),
    .Y(_04442_));
 sky130_fd_sc_hd__inv_2 _09529_ (.A(net189),
    .Y(_04443_));
 sky130_fd_sc_hd__inv_2 _09530_ (.A(net771),
    .Y(_04444_));
 sky130_fd_sc_hd__and2b_1 _09531_ (.A_N(\coreWBInterface.state[1] ),
    .B(\coreWBInterface.state[0] ),
    .X(net371));
 sky130_fd_sc_hd__and2b_1 _09532_ (.A_N(\core.cancelStall ),
    .B(\core.pipe0_fetch.currentPipeStall ),
    .X(_04445_));
 sky130_fd_sc_hd__nand2b_2 _09533_ (.A_N(\core.cancelStall ),
    .B(\core.pipe0_fetch.currentPipeStall ),
    .Y(_04446_));
 sky130_fd_sc_hd__nor2_2 _09534_ (.A(\core.pipe0_currentInstruction[4] ),
    .B(net1667),
    .Y(_04447_));
 sky130_fd_sc_hd__nand2_2 _09535_ (.A(\core.pipe0_currentInstruction[5] ),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__and3_2 _09536_ (.A(\core.pipe0_currentInstruction[6] ),
    .B(\core.pipe0_currentInstruction[5] ),
    .C(_04447_),
    .X(_04449_));
 sky130_fd_sc_hd__nand2_4 _09537_ (.A(\core.pipe0_currentInstruction[1] ),
    .B(\core.pipe0_currentInstruction[0] ),
    .Y(_04450_));
 sky130_fd_sc_hd__and3_2 _09538_ (.A(\core.pipe0_currentInstruction[2] ),
    .B(\core.pipe0_currentInstruction[1] ),
    .C(\core.pipe0_currentInstruction[0] ),
    .X(_04451_));
 sky130_fd_sc_hd__and2_2 _09539_ (.A(\core.pipe0_currentInstruction[3] ),
    .B(_04451_),
    .X(_04452_));
 sky130_fd_sc_hd__and2_1 _09540_ (.A(_04449_),
    .B(_04452_),
    .X(_04453_));
 sky130_fd_sc_hd__nand2_4 _09541_ (.A(_04449_),
    .B(_04452_),
    .Y(_04454_));
 sky130_fd_sc_hd__nor2_4 _09542_ (.A(\core.pipe0_currentInstruction[3] ),
    .B(net1668),
    .Y(_04455_));
 sky130_fd_sc_hd__nand2_4 _09543_ (.A(_04451_),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__nor2_2 _09544_ (.A(\core.pipe0_currentInstruction[6] ),
    .B(\core.pipe0_currentInstruction[5] ),
    .Y(_04457_));
 sky130_fd_sc_hd__nand2_2 _09545_ (.A(\core.pipe0_currentInstruction[4] ),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__nor2_4 _09546_ (.A(_04456_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__or2_4 _09547_ (.A(_04456_),
    .B(_04458_),
    .X(_04460_));
 sky130_fd_sc_hd__and4b_2 _09548_ (.A_N(\core.pipe0_currentInstruction[2] ),
    .B(\core.pipe0_currentInstruction[1] ),
    .C(\core.pipe0_currentInstruction[0] ),
    .D(_04455_),
    .X(_04461_));
 sky130_fd_sc_hd__or4_4 _09549_ (.A(\core.pipe0_currentInstruction[3] ),
    .B(\core.pipe0_currentInstruction[2] ),
    .C(net1667),
    .D(_04450_),
    .X(_04462_));
 sky130_fd_sc_hd__nand2_8 _09550_ (.A(net1880),
    .B(net1662),
    .Y(_04463_));
 sky130_fd_sc_hd__or2_2 _09551_ (.A(net1878),
    .B(net1882),
    .X(_04464_));
 sky130_fd_sc_hd__nor2_2 _09552_ (.A(_04463_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__a31o_4 _09553_ (.A1(net1880),
    .A2(net1666),
    .A3(_04464_),
    .B1(_04462_),
    .X(_04466_));
 sky130_fd_sc_hd__nor4_4 _09554_ (.A(net1879),
    .B(\core.pipe0_currentInstruction[6] ),
    .C(_04448_),
    .D(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__or4_4 _09555_ (.A(net1878),
    .B(\core.pipe0_currentInstruction[6] ),
    .C(_04448_),
    .D(_04466_),
    .X(_04468_));
 sky130_fd_sc_hd__or2_2 _09556_ (.A(_04458_),
    .B(_04462_),
    .X(_04469_));
 sky130_fd_sc_hd__or3_1 _09557_ (.A(\core.pipe0_currentInstruction[29] ),
    .B(net1819),
    .C(net1820),
    .X(_04470_));
 sky130_fd_sc_hd__or3_4 _09558_ (.A(net1815),
    .B(net1817),
    .C(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__or3b_1 _09559_ (.A(net1821),
    .B(net1822),
    .C_N(net1817),
    .X(_04472_));
 sky130_fd_sc_hd__or4_1 _09560_ (.A(net1815),
    .B(net1667),
    .C(_04470_),
    .D(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__or4_1 _09561_ (.A(net1815),
    .B(net1667),
    .C(_04470_),
    .D(_04472_),
    .X(_04474_));
 sky130_fd_sc_hd__o32a_2 _09562_ (.A1(net1821),
    .A2(net1822),
    .A3(_04471_),
    .B1(_04473_),
    .B2(_04423_),
    .X(_04475_));
 sky130_fd_sc_hd__and3b_4 _09563_ (.A_N(net1880),
    .B(net1881),
    .C(net1662),
    .X(_04476_));
 sky130_fd_sc_hd__or3b_4 _09564_ (.A(net1880),
    .B(net1668),
    .C_N(net1881),
    .X(_04477_));
 sky130_fd_sc_hd__a21oi_4 _09565_ (.A1(_04475_),
    .A2(_04476_),
    .B1(_04469_),
    .Y(_04478_));
 sky130_fd_sc_hd__nor3b_4 _09566_ (.A(_04466_),
    .B(\core.pipe0_currentInstruction[4] ),
    .C_N(_04457_),
    .Y(_04479_));
 sky130_fd_sc_hd__or3b_4 _09567_ (.A(_04466_),
    .B(\core.pipe0_currentInstruction[4] ),
    .C_N(_04457_),
    .X(_04480_));
 sky130_fd_sc_hd__or2_4 _09568_ (.A(_04478_),
    .B(net1274),
    .X(_04481_));
 sky130_fd_sc_hd__nor2_8 _09569_ (.A(net1275),
    .B(net1274),
    .Y(_04482_));
 sky130_fd_sc_hd__nand2_4 _09570_ (.A(_04468_),
    .B(_04480_),
    .Y(_04483_));
 sky130_fd_sc_hd__nor2_8 _09571_ (.A(_04478_),
    .B(net1241),
    .Y(_04484_));
 sky130_fd_sc_hd__or2_1 _09572_ (.A(_04478_),
    .B(net1241),
    .X(_04485_));
 sky130_fd_sc_hd__a21oi_1 _09573_ (.A1(net1815),
    .A2(net1192),
    .B1(net1285),
    .Y(_04486_));
 sky130_fd_sc_hd__nand2b_4 _09574_ (.A_N(net1884),
    .B(\core.csr.currentInstruction[12] ),
    .Y(_04487_));
 sky130_fd_sc_hd__nor2_4 _09575_ (.A(net1885),
    .B(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__or4bb_1 _09576_ (.A(net1883),
    .B(net1885),
    .C_N(\core.csr.currentInstruction[12] ),
    .D_N(\core.csr.currentInstruction[14] ),
    .X(_04489_));
 sky130_fd_sc_hd__o21ba_2 _09577_ (.A1(net1885),
    .A2(\core.csr.currentInstruction[12] ),
    .B1_N(net1883),
    .X(_04490_));
 sky130_fd_sc_hd__o211a_1 _09578_ (.A1(\core.csr.currentInstruction[14] ),
    .A2(_04490_),
    .B1(_04489_),
    .C1(\core.csr.currentInstruction[30] ),
    .X(_04491_));
 sky130_fd_sc_hd__or2_2 _09579_ (.A(\core.csr.currentInstruction[27] ),
    .B(\core.csr.currentInstruction[26] ),
    .X(_04492_));
 sky130_fd_sc_hd__or4_2 _09580_ (.A(\core.csr.currentInstruction[31] ),
    .B(\core.csr.currentInstruction[29] ),
    .C(\core.csr.currentInstruction[28] ),
    .D(\core.csr.currentInstruction[25] ),
    .X(_04493_));
 sky130_fd_sc_hd__o32ai_4 _09581_ (.A1(_04491_),
    .A2(_04492_),
    .A3(_04493_),
    .B1(_04488_),
    .B2(\core.csr.currentInstruction[5] ),
    .Y(_04494_));
 sky130_fd_sc_hd__and3b_2 _09582_ (.A_N(net1884),
    .B(\core.csr.currentInstruction[1] ),
    .C(\core.csr.currentInstruction[0] ),
    .X(_04495_));
 sky130_fd_sc_hd__and3_1 _09583_ (.A(_04427_),
    .B(_04428_),
    .C(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__or3b_4 _09584_ (.A(\core.csr.currentInstruction[3] ),
    .B(\core.csr.currentInstruction[2] ),
    .C_N(_04495_),
    .X(_04497_));
 sky130_fd_sc_hd__and4_4 _09585_ (.A(_04426_),
    .B(\core.csr.currentInstruction[4] ),
    .C(_04494_),
    .D(_04496_),
    .X(_04498_));
 sky130_fd_sc_hd__inv_2 _09586_ (.A(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__and4bb_1 _09587_ (.A_N(net1884),
    .B_N(\core.csr.currentInstruction[4] ),
    .C(\core.csr.currentInstruction[5] ),
    .D(\core.csr.currentInstruction[6] ),
    .X(_04500_));
 sky130_fd_sc_hd__and4_1 _09588_ (.A(\core.csr.currentInstruction[3] ),
    .B(\core.csr.currentInstruction[2] ),
    .C(_04495_),
    .D(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__o21a_1 _09589_ (.A1(\core.csr.currentInstruction[14] ),
    .A2(net1885),
    .B1(_04391_),
    .X(_04502_));
 sky130_fd_sc_hd__o21bai_4 _09590_ (.A1(\core.csr.currentInstruction[14] ),
    .A2(net1885),
    .B1_N(net1883),
    .Y(_04503_));
 sky130_fd_sc_hd__nand2_1 _09591_ (.A(_04487_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__and3_1 _09592_ (.A(_04487_),
    .B(_04500_),
    .C(_04503_),
    .X(_04505_));
 sky130_fd_sc_hd__a31o_1 _09593_ (.A1(_04391_),
    .A2(_04426_),
    .A3(\core.csr.currentInstruction[4] ),
    .B1(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__a41o_2 _09594_ (.A1(_04427_),
    .A2(\core.csr.currentInstruction[2] ),
    .A3(_04495_),
    .A4(_04506_),
    .B1(_04501_),
    .X(_04507_));
 sky130_fd_sc_hd__inv_2 _09595_ (.A(net1271),
    .Y(_04508_));
 sky130_fd_sc_hd__or2_1 _09596_ (.A(_04498_),
    .B(net1271),
    .X(_04509_));
 sky130_fd_sc_hd__and2b_4 _09597_ (.A_N(net1883),
    .B(\core.csr.currentInstruction[7] ),
    .X(_04510_));
 sky130_fd_sc_hd__nand2b_4 _09598_ (.A_N(net1883),
    .B(\core.csr.currentInstruction[8] ),
    .Y(_04511_));
 sky130_fd_sc_hd__nand2b_4 _09599_ (.A_N(_04510_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__nand2b_4 _09600_ (.A_N(net1883),
    .B(\core.csr.currentInstruction[11] ),
    .Y(_04513_));
 sky130_fd_sc_hd__nand2b_4 _09601_ (.A_N(net1883),
    .B(\core.csr.currentInstruction[10] ),
    .Y(_04514_));
 sky130_fd_sc_hd__nand2b_4 _09602_ (.A_N(net1883),
    .B(\core.csr.currentInstruction[9] ),
    .Y(_04515_));
 sky130_fd_sc_hd__nand3_4 _09603_ (.A(_04513_),
    .B(_04514_),
    .C(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__or3_2 _09604_ (.A(_04488_),
    .B(_04512_),
    .C(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__and4_1 _09605_ (.A(_04391_),
    .B(\core.csr.currentInstruction[6] ),
    .C(\core.csr.currentInstruction[5] ),
    .D(\core.csr.currentInstruction[4] ),
    .X(_04518_));
 sky130_fd_sc_hd__nand2_1 _09606_ (.A(_04496_),
    .B(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__and3b_4 _09607_ (.A_N(_04519_),
    .B(_04517_),
    .C(_04504_),
    .X(_04520_));
 sky130_fd_sc_hd__o31a_4 _09608_ (.A1(\core.csr.currentInstruction[6] ),
    .A2(\core.csr.currentInstruction[5] ),
    .A3(\core.csr.currentInstruction[4] ),
    .B1(_04391_),
    .X(_04521_));
 sky130_fd_sc_hd__or4b_4 _09609_ (.A(net1883),
    .B(\core.csr.currentInstruction[14] ),
    .C(\core.csr.currentInstruction[12] ),
    .D_N(net1885),
    .X(_04522_));
 sky130_fd_sc_hd__and3_2 _09610_ (.A(_04391_),
    .B(net1885),
    .C(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__or3_4 _09611_ (.A(_04497_),
    .B(_04521_),
    .C(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__or3_4 _09612_ (.A(_04497_),
    .B(_04521_),
    .C(_04523_),
    .X(_04525_));
 sky130_fd_sc_hd__or3b_4 _09613_ (.A(net1239),
    .B(net1270),
    .C_N(_04524_),
    .X(_04526_));
 sky130_fd_sc_hd__and2_4 _09614_ (.A(net1831),
    .B(net1664),
    .X(_04527_));
 sky130_fd_sc_hd__nand2_8 _09615_ (.A(net1831),
    .B(net1663),
    .Y(_04528_));
 sky130_fd_sc_hd__nor2_1 _09616_ (.A(_04514_),
    .B(net1637),
    .Y(_04529_));
 sky130_fd_sc_hd__nor2_2 _09617_ (.A(net1743),
    .B(net1667),
    .Y(_04530_));
 sky130_fd_sc_hd__nand2_8 _09618_ (.A(net1846),
    .B(net1663),
    .Y(_04531_));
 sky130_fd_sc_hd__a2bb2o_1 _09619_ (.A1_N(_04511_),
    .A2_N(net1623),
    .B1(net1637),
    .B2(_04514_),
    .X(_04532_));
 sky130_fd_sc_hd__a211o_1 _09620_ (.A1(_04511_),
    .A2(net1623),
    .B1(_04532_),
    .C1(_04529_),
    .X(_04533_));
 sky130_fd_sc_hd__nor2_1 _09621_ (.A(net1746),
    .B(net1667),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_1 _09622_ (.A(net1836),
    .B(net1663),
    .Y(_04535_));
 sky130_fd_sc_hd__xnor2_1 _09623_ (.A(_04515_),
    .B(net1591),
    .Y(_04536_));
 sky130_fd_sc_hd__nor2_8 _09624_ (.A(net1752),
    .B(net1668),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_8 _09625_ (.A(net1827),
    .B(net1663),
    .Y(_04538_));
 sky130_fd_sc_hd__xnor2_1 _09626_ (.A(_04513_),
    .B(net1573),
    .Y(_04539_));
 sky130_fd_sc_hd__nor2_1 _09627_ (.A(net1730),
    .B(net1667),
    .Y(_04540_));
 sky130_fd_sc_hd__nand2_1 _09628_ (.A(net1850),
    .B(net1663),
    .Y(_04541_));
 sky130_fd_sc_hd__xnor2_1 _09629_ (.A(_04510_),
    .B(net1499),
    .Y(_04542_));
 sky130_fd_sc_hd__or4_1 _09630_ (.A(_04533_),
    .B(_04536_),
    .C(_04539_),
    .D(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__and2b_4 _09631_ (.A_N(_04543_),
    .B(_04526_),
    .X(_04544_));
 sky130_fd_sc_hd__nand2b_4 _09632_ (.A_N(_04543_),
    .B(_04526_),
    .Y(_04545_));
 sky130_fd_sc_hd__a22o_1 _09633_ (.A1(\core.pipe1_resultRegister[23] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[23] ),
    .X(_04546_));
 sky130_fd_sc_hd__or4b_1 _09634_ (.A(net1884),
    .B(\core.csr.currentInstruction[6] ),
    .C(\core.csr.currentInstruction[4] ),
    .D_N(\core.csr.currentInstruction[5] ),
    .X(_04547_));
 sky130_fd_sc_hd__a211o_4 _09635_ (.A1(_04502_),
    .A2(_04522_),
    .B1(_04547_),
    .C1(_04497_),
    .X(_04548_));
 sky130_fd_sc_hd__nand2_1 _09636_ (.A(_04524_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__a21oi_4 _09637_ (.A1(_04525_),
    .A2(_04548_),
    .B1(_04522_),
    .Y(_04550_));
 sky130_fd_sc_hd__nand2_8 _09638_ (.A(_04401_),
    .B(net1810),
    .Y(_04551_));
 sky130_fd_sc_hd__a21bo_1 _09639_ (.A1(net1810),
    .A2(_04490_),
    .B1_N(_04522_),
    .X(_04552_));
 sky130_fd_sc_hd__nand2_1 _09640_ (.A(net1806),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__a21o_1 _09641_ (.A1(_04525_),
    .A2(_04548_),
    .B1(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__a2bb2oi_4 _09642_ (.A1_N(net1806),
    .A2_N(_04550_),
    .B1(_04551_),
    .B2(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__nor2_1 _09643_ (.A(_04524_),
    .B(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__and2_4 _09644_ (.A(net1806),
    .B(net1810),
    .X(_04557_));
 sky130_fd_sc_hd__nand2_8 _09645_ (.A(net1807),
    .B(net1811),
    .Y(_04558_));
 sky130_fd_sc_hd__nand2_2 _09646_ (.A(\localMemoryInterface.lastCoreByteSelect[3] ),
    .B(\localMemoryInterface.coreReadReady ),
    .Y(_04559_));
 sky130_fd_sc_hd__mux2_8 _09647_ (.A0(net131),
    .A1(net166),
    .S(net1805),
    .X(_04560_));
 sky130_fd_sc_hd__nand2b_4 _09648_ (.A_N(\memoryController.last_data_enableLocalMemory ),
    .B(\memoryController.last_data_enableWB ),
    .Y(_04561_));
 sky130_fd_sc_hd__or3b_4 _09649_ (.A(\coreWBInterface.readDataBuffered[31] ),
    .B(\memoryController.last_data_enableLocalMemory ),
    .C_N(\memoryController.last_data_enableWB ),
    .X(_04562_));
 sky130_fd_sc_hd__o31a_1 _09650_ (.A1(net1674),
    .A2(net1661),
    .A3(_04560_),
    .B1(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__nand2_1 _09651_ (.A(\core.pipe1_loadResult[31] ),
    .B(net1813),
    .Y(_04564_));
 sky130_fd_sc_hd__o311ai_4 _09652_ (.A1(net1673),
    .A2(net1661),
    .A3(_04560_),
    .B1(_04562_),
    .C1(net1757),
    .Y(_04565_));
 sky130_fd_sc_hd__nand2_1 _09653_ (.A(_04564_),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__a21oi_1 _09654_ (.A1(_04564_),
    .A2(_04565_),
    .B1(_04558_),
    .Y(_04567_));
 sky130_fd_sc_hd__nand2_4 _09655_ (.A(\localMemoryInterface.coreReadReady ),
    .B(\localMemoryInterface.lastCoreByteSelect[0] ),
    .Y(_04568_));
 sky130_fd_sc_hd__mux2_8 _09656_ (.A0(net168),
    .A1(net139),
    .S(net1805),
    .X(_04569_));
 sky130_fd_sc_hd__o32a_1 _09657_ (.A1(net1674),
    .A2(net1656),
    .A3(_04569_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[7] ),
    .X(_04570_));
 sky130_fd_sc_hd__nor2_8 _09658_ (.A(net1807),
    .B(net1811),
    .Y(_04571_));
 sky130_fd_sc_hd__or2_4 _09659_ (.A(net1808),
    .B(net1811),
    .X(_04572_));
 sky130_fd_sc_hd__or2_1 _09660_ (.A(\core.pipe1_loadResult[7] ),
    .B(net1758),
    .X(_04573_));
 sky130_fd_sc_hd__o211a_1 _09661_ (.A1(net1813),
    .A2(_04570_),
    .B1(_04571_),
    .C1(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__nand2_2 _09662_ (.A(\localMemoryInterface.coreReadReady ),
    .B(\localMemoryInterface.lastCoreByteSelect[1] ),
    .Y(_04575_));
 sky130_fd_sc_hd__mux2_8 _09663_ (.A0(net113),
    .A1(net148),
    .S(net1805),
    .X(_04576_));
 sky130_fd_sc_hd__or3_1 _09664_ (.A(net1675),
    .B(net1653),
    .C(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__or3b_4 _09665_ (.A(\coreWBInterface.readDataBuffered[15] ),
    .B(\memoryController.last_data_enableLocalMemory ),
    .C_N(\memoryController.last_data_enableWB ),
    .X(_04578_));
 sky130_fd_sc_hd__nand2_1 _09666_ (.A(\core.pipe1_loadResult[15] ),
    .B(net1813),
    .Y(_04579_));
 sky130_fd_sc_hd__o311ai_4 _09667_ (.A1(net1673),
    .A2(net1654),
    .A3(_04576_),
    .B1(_04578_),
    .C1(net1758),
    .Y(_04580_));
 sky130_fd_sc_hd__a21oi_1 _09668_ (.A1(_04579_),
    .A2(_04580_),
    .B1(_04551_),
    .Y(_04581_));
 sky130_fd_sc_hd__or2_4 _09669_ (.A(_04401_),
    .B(net1810),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_4 _09670_ (.A(\localMemoryInterface.coreReadReady ),
    .B(\localMemoryInterface.lastCoreByteSelect[2] ),
    .Y(_04583_));
 sky130_fd_sc_hd__mux2_8 _09671_ (.A0(net122),
    .A1(net157),
    .S(net1805),
    .X(_04584_));
 sky130_fd_sc_hd__or3_1 _09672_ (.A(net1675),
    .B(net1652),
    .C(_04584_),
    .X(_04585_));
 sky130_fd_sc_hd__or3b_4 _09673_ (.A(\coreWBInterface.readDataBuffered[23] ),
    .B(\memoryController.last_data_enableLocalMemory ),
    .C_N(\memoryController.last_data_enableWB ),
    .X(_04586_));
 sky130_fd_sc_hd__nand2_1 _09674_ (.A(\core.pipe1_loadResult[23] ),
    .B(net1812),
    .Y(_04587_));
 sky130_fd_sc_hd__o311ai_4 _09675_ (.A1(net1673),
    .A2(net1651),
    .A3(_04584_),
    .B1(_04586_),
    .C1(net1757),
    .Y(_04588_));
 sky130_fd_sc_hd__nand2_2 _09676_ (.A(_04587_),
    .B(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__a21oi_1 _09677_ (.A1(_04587_),
    .A2(_04588_),
    .B1(_04582_),
    .Y(_04590_));
 sky130_fd_sc_hd__or4_4 _09678_ (.A(_04567_),
    .B(_04574_),
    .C(_04581_),
    .D(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__a21o_1 _09679_ (.A1(_04587_),
    .A2(_04588_),
    .B1(net1807),
    .X(_04592_));
 sky130_fd_sc_hd__and3_1 _09680_ (.A(_04571_),
    .B(_04579_),
    .C(_04580_),
    .X(_04593_));
 sky130_fd_sc_hd__and3_1 _09681_ (.A(net1808),
    .B(_04564_),
    .C(_04565_),
    .X(_04594_));
 sky130_fd_sc_hd__a211oi_2 _09682_ (.A1(net1811),
    .A2(_04592_),
    .B1(_04593_),
    .C1(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__o221a_4 _09683_ (.A1(_04490_),
    .A2(_04591_),
    .B1(_04595_),
    .B2(_04487_),
    .C1(_04503_),
    .X(_04596_));
 sky130_fd_sc_hd__and2_1 _09684_ (.A(_04550_),
    .B(_04571_),
    .X(_04597_));
 sky130_fd_sc_hd__a21o_4 _09685_ (.A1(_04589_),
    .A2(net1234),
    .B1(net1236),
    .X(_04598_));
 sky130_fd_sc_hd__nor4_4 _09686_ (.A(_04497_),
    .B(_04521_),
    .C(_04523_),
    .D(_04555_),
    .Y(_04599_));
 sky130_fd_sc_hd__a21o_1 _09687_ (.A1(net1188),
    .A2(_04598_),
    .B1(_04546_),
    .X(_04600_));
 sky130_fd_sc_hd__nand2_2 _09688_ (.A(net1580),
    .B(net1498),
    .Y(_04601_));
 sky130_fd_sc_hd__or4_4 _09689_ (.A(net1637),
    .B(net1623),
    .C(net1573),
    .D(net1339),
    .X(_04602_));
 sky130_fd_sc_hd__or2_1 _09690_ (.A(\core.registers[1][23] ),
    .B(net1494),
    .X(_04603_));
 sky130_fd_sc_hd__or2_1 _09691_ (.A(\core.registers[6][23] ),
    .B(net1511),
    .X(_04604_));
 sky130_fd_sc_hd__or2_1 _09692_ (.A(\core.registers[17][23] ),
    .B(net1495),
    .X(_04605_));
 sky130_fd_sc_hd__or2_1 _09693_ (.A(\core.registers[29][23] ),
    .B(net1493),
    .X(_04606_));
 sky130_fd_sc_hd__o211a_1 _09694_ (.A1(\core.registers[28][23] ),
    .A2(net1513),
    .B1(_04606_),
    .C1(net1736),
    .X(_04607_));
 sky130_fd_sc_hd__nor2_8 _09695_ (.A(net1742),
    .B(net1851),
    .Y(_04608_));
 sky130_fd_sc_hd__a31o_1 _09696_ (.A1(net1840),
    .A2(net1720),
    .A3(\core.registers[30][23] ),
    .B1(net1748),
    .X(_04609_));
 sky130_fd_sc_hd__a31o_1 _09697_ (.A1(net1840),
    .A2(\core.registers[31][23] ),
    .A3(net1513),
    .B1(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__mux2_1 _09698_ (.A0(\core.registers[8][23] ),
    .A1(\core.registers[9][23] ),
    .S(net1509),
    .X(_04611_));
 sky130_fd_sc_hd__mux2_1 _09699_ (.A0(\core.registers[10][23] ),
    .A1(\core.registers[11][23] ),
    .S(net1509),
    .X(_04612_));
 sky130_fd_sc_hd__mux2_1 _09700_ (.A0(\core.registers[24][23] ),
    .A1(\core.registers[25][23] ),
    .S(net1509),
    .X(_04613_));
 sky130_fd_sc_hd__a221o_1 _09701_ (.A1(net1720),
    .A2(\core.registers[26][23] ),
    .B1(\core.registers[27][23] ),
    .B2(net1509),
    .C1(net1735),
    .X(_04614_));
 sky130_fd_sc_hd__mux2_1 _09702_ (.A0(\core.registers[12][23] ),
    .A1(\core.registers[13][23] ),
    .S(net1509),
    .X(_04615_));
 sky130_fd_sc_hd__mux2_1 _09703_ (.A0(\core.registers[14][23] ),
    .A1(\core.registers[15][23] ),
    .S(net1509),
    .X(_04616_));
 sky130_fd_sc_hd__mux2_1 _09704_ (.A0(_04615_),
    .A1(_04616_),
    .S(net1612),
    .X(_04617_));
 sky130_fd_sc_hd__o221a_1 _09705_ (.A1(_04607_),
    .A2(_04610_),
    .B1(_04617_),
    .B2(net1823),
    .C1(net1832),
    .X(_04618_));
 sky130_fd_sc_hd__mux2_1 _09706_ (.A0(_04611_),
    .A1(_04612_),
    .S(net1612),
    .X(_04619_));
 sky130_fd_sc_hd__o21a_1 _09707_ (.A1(net1838),
    .A2(_04613_),
    .B1(_04614_),
    .X(_04620_));
 sky130_fd_sc_hd__mux2_1 _09708_ (.A0(_04619_),
    .A1(_04620_),
    .S(net1823),
    .X(_04621_));
 sky130_fd_sc_hd__a211o_2 _09709_ (.A1(net1744),
    .A2(_04621_),
    .B1(_04618_),
    .C1(net1631),
    .X(_04622_));
 sky130_fd_sc_hd__o211a_1 _09710_ (.A1(net1720),
    .A2(\core.registers[7][23] ),
    .B1(net1613),
    .C1(_04604_),
    .X(_04623_));
 sky130_fd_sc_hd__mux2_1 _09711_ (.A0(\core.registers[4][23] ),
    .A1(\core.registers[5][23] ),
    .S(net1512),
    .X(_04624_));
 sky130_fd_sc_hd__a211o_1 _09712_ (.A1(net1597),
    .A2(_04624_),
    .B1(_04623_),
    .C1(net1576),
    .X(_04625_));
 sky130_fd_sc_hd__o211a_1 _09713_ (.A1(\core.registers[0][23] ),
    .A2(net1521),
    .B1(_04603_),
    .C1(net1601),
    .X(_04626_));
 sky130_fd_sc_hd__mux2_1 _09714_ (.A0(\core.registers[2][23] ),
    .A1(\core.registers[3][23] ),
    .S(net1520),
    .X(_04627_));
 sky130_fd_sc_hd__a211o_1 _09715_ (.A1(net1616),
    .A2(_04627_),
    .B1(_04626_),
    .C1(net1587),
    .X(_04628_));
 sky130_fd_sc_hd__o211a_1 _09716_ (.A1(\core.registers[16][23] ),
    .A2(net1511),
    .B1(_04605_),
    .C1(net1597),
    .X(_04629_));
 sky130_fd_sc_hd__mux2_1 _09717_ (.A0(\core.registers[18][23] ),
    .A1(\core.registers[19][23] ),
    .S(net1511),
    .X(_04630_));
 sky130_fd_sc_hd__a211o_1 _09718_ (.A1(net1612),
    .A2(_04630_),
    .B1(_04629_),
    .C1(net1587),
    .X(_04631_));
 sky130_fd_sc_hd__mux2_1 _09719_ (.A0(\core.registers[22][23] ),
    .A1(\core.registers[23][23] ),
    .S(net1509),
    .X(_04632_));
 sky130_fd_sc_hd__mux2_1 _09720_ (.A0(\core.registers[20][23] ),
    .A1(\core.registers[21][23] ),
    .S(net1510),
    .X(_04633_));
 sky130_fd_sc_hd__mux2_1 _09721_ (.A0(_04632_),
    .A1(_04633_),
    .S(net1597),
    .X(_04634_));
 sky130_fd_sc_hd__o211a_1 _09722_ (.A1(net1576),
    .A2(_04634_),
    .B1(_04631_),
    .C1(net1571),
    .X(_04635_));
 sky130_fd_sc_hd__a311o_1 _09723_ (.A1(net1567),
    .A2(_04625_),
    .A3(_04628_),
    .B1(_04635_),
    .C1(net1635),
    .X(_04636_));
 sky130_fd_sc_hd__a21o_1 _09724_ (.A1(_04622_),
    .A2(_04636_),
    .B1(net1157),
    .X(_04637_));
 sky130_fd_sc_hd__o211ai_2 _09725_ (.A1(net1153),
    .A2(net1152),
    .B1(net1263),
    .C1(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__o21ai_1 _09726_ (.A1(net1192),
    .A2(_04638_),
    .B1(net1161),
    .Y(_04639_));
 sky130_fd_sc_hd__o21a_1 _09727_ (.A1(net1831),
    .A2(net1278),
    .B1(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__and2_4 _09728_ (.A(\core.pipe0_currentInstruction[18] ),
    .B(net1665),
    .X(_04641_));
 sky130_fd_sc_hd__nand2_8 _09729_ (.A(\core.pipe0_currentInstruction[18] ),
    .B(net1665),
    .Y(_04642_));
 sky130_fd_sc_hd__nor2_2 _09730_ (.A(net1708),
    .B(net1667),
    .Y(_04643_));
 sky130_fd_sc_hd__nand2_2 _09731_ (.A(net1877),
    .B(net1663),
    .Y(_04644_));
 sky130_fd_sc_hd__nor2_8 _09732_ (.A(net1716),
    .B(net1667),
    .Y(_04645_));
 sky130_fd_sc_hd__nand2_8 _09733_ (.A(net1860),
    .B(net1663),
    .Y(_04646_));
 sky130_fd_sc_hd__nor2_8 _09734_ (.A(net1715),
    .B(net1667),
    .Y(_04647_));
 sky130_fd_sc_hd__nand2_8 _09735_ (.A(net1866),
    .B(net1663),
    .Y(_04648_));
 sky130_fd_sc_hd__nor2_8 _09736_ (.A(net1694),
    .B(net1668),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_2 _09737_ (.A(\core.pipe0_currentInstruction[15] ),
    .B(net1665),
    .Y(_04650_));
 sky130_fd_sc_hd__nand2_8 _09738_ (.A(net1440),
    .B(net1378),
    .Y(_04651_));
 sky130_fd_sc_hd__and4b_2 _09739_ (.A_N(net1334),
    .B(net1462),
    .C(net1477),
    .D(net1488),
    .X(_04652_));
 sky130_fd_sc_hd__xnor2_1 _09740_ (.A(_04511_),
    .B(net1483),
    .Y(_04653_));
 sky130_fd_sc_hd__nor2_1 _09741_ (.A(_04515_),
    .B(net1454),
    .Y(_04654_));
 sky130_fd_sc_hd__and3_1 _09742_ (.A(net1866),
    .B(net1665),
    .C(_04515_),
    .X(_04655_));
 sky130_fd_sc_hd__o22a_1 _09743_ (.A1(_04514_),
    .A2(net1492),
    .B1(net1377),
    .B2(_04510_),
    .X(_04656_));
 sky130_fd_sc_hd__xnor2_1 _09744_ (.A(_04513_),
    .B(_04645_),
    .Y(_04657_));
 sky130_fd_sc_hd__a22o_1 _09745_ (.A1(_04514_),
    .A2(net1492),
    .B1(net1377),
    .B2(_04510_),
    .X(_04658_));
 sky130_fd_sc_hd__or4b_1 _09746_ (.A(_04653_),
    .B(_04657_),
    .C(_04658_),
    .D_N(_04656_),
    .X(_04659_));
 sky130_fd_sc_hd__or4b_4 _09747_ (.A(_04654_),
    .B(_04659_),
    .C(_04655_),
    .D_N(_04526_),
    .X(_04660_));
 sky130_fd_sc_hd__nor2_4 _09748_ (.A(_04652_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__and2b_1 _09749_ (.A_N(_04652_),
    .B(_04660_),
    .X(_04662_));
 sky130_fd_sc_hd__nand2b_4 _09750_ (.A_N(_04652_),
    .B(_04660_),
    .Y(_04663_));
 sky130_fd_sc_hd__o22a_1 _09751_ (.A1(net1679),
    .A2(\core.registers[23][23] ),
    .B1(net1385),
    .B2(\core.registers[22][23] ),
    .X(_04664_));
 sky130_fd_sc_hd__or3_1 _09752_ (.A(net1679),
    .B(\core.registers[19][23] ),
    .C(net1442),
    .X(_04665_));
 sky130_fd_sc_hd__o221a_1 _09753_ (.A1(\core.registers[18][23] ),
    .A2(net1331),
    .B1(_04664_),
    .B2(net1431),
    .C1(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__mux4_1 _09754_ (.A0(\core.registers[16][23] ),
    .A1(\core.registers[17][23] ),
    .A2(\core.registers[20][23] ),
    .A3(\core.registers[21][23] ),
    .S0(net1385),
    .S1(net1442),
    .X(_04667_));
 sky130_fd_sc_hd__mux2_1 _09755_ (.A0(_04666_),
    .A1(_04667_),
    .S(net1465),
    .X(_04668_));
 sky130_fd_sc_hd__o22a_1 _09756_ (.A1(net1680),
    .A2(\core.registers[7][23] ),
    .B1(net1392),
    .B2(\core.registers[6][23] ),
    .X(_04669_));
 sky130_fd_sc_hd__or3_1 _09757_ (.A(net1680),
    .B(\core.registers[3][23] ),
    .C(net1443),
    .X(_04670_));
 sky130_fd_sc_hd__o221a_1 _09758_ (.A1(\core.registers[2][23] ),
    .A2(net1333),
    .B1(_04669_),
    .B2(net1433),
    .C1(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__mux4_1 _09759_ (.A0(\core.registers[0][23] ),
    .A1(\core.registers[1][23] ),
    .A2(\core.registers[4][23] ),
    .A3(\core.registers[5][23] ),
    .S0(net1393),
    .S1(net1443),
    .X(_04672_));
 sky130_fd_sc_hd__mux2_1 _09760_ (.A0(_04671_),
    .A1(_04672_),
    .S(net1466),
    .X(_04673_));
 sky130_fd_sc_hd__mux2_1 _09761_ (.A0(_04668_),
    .A1(_04673_),
    .S(net1460),
    .X(_04674_));
 sky130_fd_sc_hd__a221o_1 _09762_ (.A1(net1679),
    .A2(\core.registers[26][23] ),
    .B1(\core.registers[27][23] ),
    .B2(net1383),
    .C1(net1704),
    .X(_04675_));
 sky130_fd_sc_hd__mux2_1 _09763_ (.A0(\core.registers[24][23] ),
    .A1(\core.registers[25][23] ),
    .S(net1383),
    .X(_04676_));
 sky130_fd_sc_hd__o21ai_1 _09764_ (.A1(net1868),
    .A2(_04676_),
    .B1(_04675_),
    .Y(_04677_));
 sky130_fd_sc_hd__a221o_1 _09765_ (.A1(net1679),
    .A2(\core.registers[10][23] ),
    .B1(\core.registers[11][23] ),
    .B2(net1383),
    .C1(net1705),
    .X(_04678_));
 sky130_fd_sc_hd__a21o_1 _09766_ (.A1(\core.registers[8][23] ),
    .A2(net1373),
    .B1(net1869),
    .X(_04679_));
 sky130_fd_sc_hd__a21o_1 _09767_ (.A1(\core.registers[9][23] ),
    .A2(net1383),
    .B1(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__a21oi_1 _09768_ (.A1(_04678_),
    .A2(_04680_),
    .B1(net1854),
    .Y(_04681_));
 sky130_fd_sc_hd__a211o_1 _09769_ (.A1(net1854),
    .A2(_04677_),
    .B1(_04681_),
    .C1(net1862),
    .X(_04682_));
 sky130_fd_sc_hd__mux2_1 _09770_ (.A0(\core.registers[12][23] ),
    .A1(\core.registers[13][23] ),
    .S(net1383),
    .X(_04683_));
 sky130_fd_sc_hd__mux2_1 _09771_ (.A0(\core.registers[14][23] ),
    .A1(\core.registers[15][23] ),
    .S(net1383),
    .X(_04684_));
 sky130_fd_sc_hd__mux2_1 _09772_ (.A0(_04683_),
    .A1(_04684_),
    .S(net1480),
    .X(_04685_));
 sky130_fd_sc_hd__a221o_1 _09773_ (.A1(net1681),
    .A2(\core.registers[30][23] ),
    .B1(\core.registers[31][23] ),
    .B2(net1384),
    .C1(net1705),
    .X(_04686_));
 sky130_fd_sc_hd__mux2_1 _09774_ (.A0(\core.registers[28][23] ),
    .A1(\core.registers[29][23] ),
    .S(net1384),
    .X(_04687_));
 sky130_fd_sc_hd__o21a_1 _09775_ (.A1(net1869),
    .A2(_04687_),
    .B1(_04686_),
    .X(_04688_));
 sky130_fd_sc_hd__mux2_1 _09776_ (.A0(_04685_),
    .A1(_04688_),
    .S(net1854),
    .X(_04689_));
 sky130_fd_sc_hd__a21oi_1 _09777_ (.A1(net1863),
    .A2(_04689_),
    .B1(net1484),
    .Y(_04690_));
 sky130_fd_sc_hd__o2bb2a_2 _09778_ (.A1_N(_04682_),
    .A2_N(_04690_),
    .B1(net1489),
    .B2(_04674_),
    .X(_04691_));
 sky130_fd_sc_hd__a22o_2 _09779_ (.A1(net1152),
    .A2(net1068),
    .B1(net1065),
    .B2(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__mux2_8 _09780_ (.A0(net465),
    .A1(_04692_),
    .S(net1276),
    .X(_04693_));
 sky130_fd_sc_hd__or2_4 _09781_ (.A(_04640_),
    .B(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__clkinv_2 _09782_ (.A(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__and2_4 _09783_ (.A(_04640_),
    .B(_04693_),
    .X(_04696_));
 sky130_fd_sc_hd__nor2_8 _09784_ (.A(_04695_),
    .B(_04696_),
    .Y(_04697_));
 sky130_fd_sc_hd__a22o_1 _09785_ (.A1(\core.pipe1_resultRegister[22] ),
    .A2(net1239),
    .B1(net1270),
    .B2(\core.pipe1_csrData[22] ),
    .X(_04698_));
 sky130_fd_sc_hd__mux2_8 _09786_ (.A0(net121),
    .A1(net156),
    .S(net1805),
    .X(_04699_));
 sky130_fd_sc_hd__o32a_1 _09787_ (.A1(net1675),
    .A2(net1651),
    .A3(_04699_),
    .B1(net1659),
    .B2(\coreWBInterface.readDataBuffered[22] ),
    .X(_04700_));
 sky130_fd_sc_hd__mux2_2 _09788_ (.A0(\core.pipe1_loadResult[22] ),
    .A1(_04700_),
    .S(net1757),
    .X(_04701_));
 sky130_fd_sc_hd__a21o_2 _09789_ (.A1(net1235),
    .A2(_04701_),
    .B1(net1237),
    .X(_04702_));
 sky130_fd_sc_hd__a21o_4 _09790_ (.A1(net1191),
    .A2(_04702_),
    .B1(_04698_),
    .X(_04703_));
 sky130_fd_sc_hd__mux2_1 _09791_ (.A0(\core.registers[8][22] ),
    .A1(\core.registers[9][22] ),
    .S(net1528),
    .X(_04704_));
 sky130_fd_sc_hd__mux2_1 _09792_ (.A0(\core.registers[10][22] ),
    .A1(\core.registers[11][22] ),
    .S(net1528),
    .X(_04705_));
 sky130_fd_sc_hd__mux2_1 _09793_ (.A0(\core.registers[24][22] ),
    .A1(\core.registers[25][22] ),
    .S(net1528),
    .X(_04706_));
 sky130_fd_sc_hd__a221o_1 _09794_ (.A1(net1723),
    .A2(\core.registers[26][22] ),
    .B1(\core.registers[27][22] ),
    .B2(net1528),
    .C1(net1737),
    .X(_04707_));
 sky130_fd_sc_hd__or2_1 _09795_ (.A(\core.registers[29][22] ),
    .B(net1497),
    .X(_04708_));
 sky130_fd_sc_hd__o211a_1 _09796_ (.A1(\core.registers[28][22] ),
    .A2(net1528),
    .B1(_04708_),
    .C1(net1737),
    .X(_04709_));
 sky130_fd_sc_hd__a31o_1 _09797_ (.A1(net1841),
    .A2(net1723),
    .A3(\core.registers[30][22] ),
    .B1(net1749),
    .X(_04710_));
 sky130_fd_sc_hd__a31o_1 _09798_ (.A1(net1841),
    .A2(\core.registers[31][22] ),
    .A3(net1528),
    .B1(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__or2_1 _09799_ (.A(\core.registers[1][22] ),
    .B(net1497),
    .X(_04712_));
 sky130_fd_sc_hd__or2_1 _09800_ (.A(\core.registers[6][22] ),
    .B(net1527),
    .X(_04713_));
 sky130_fd_sc_hd__or2_1 _09801_ (.A(\core.registers[17][22] ),
    .B(net1497),
    .X(_04714_));
 sky130_fd_sc_hd__mux2_1 _09802_ (.A0(\core.registers[12][22] ),
    .A1(\core.registers[13][22] ),
    .S(net1529),
    .X(_04715_));
 sky130_fd_sc_hd__mux2_1 _09803_ (.A0(\core.registers[14][22] ),
    .A1(\core.registers[15][22] ),
    .S(net1529),
    .X(_04716_));
 sky130_fd_sc_hd__mux2_1 _09804_ (.A0(_04715_),
    .A1(_04716_),
    .S(net1618),
    .X(_04717_));
 sky130_fd_sc_hd__o221a_1 _09805_ (.A1(_04709_),
    .A2(_04711_),
    .B1(_04717_),
    .B2(net1825),
    .C1(net1833),
    .X(_04718_));
 sky130_fd_sc_hd__mux2_1 _09806_ (.A0(_04704_),
    .A1(_04705_),
    .S(net1618),
    .X(_04719_));
 sky130_fd_sc_hd__o21a_1 _09807_ (.A1(net1842),
    .A2(_04706_),
    .B1(_04707_),
    .X(_04720_));
 sky130_fd_sc_hd__mux2_1 _09808_ (.A0(_04719_),
    .A1(_04720_),
    .S(net1825),
    .X(_04721_));
 sky130_fd_sc_hd__a211o_1 _09809_ (.A1(net1745),
    .A2(_04721_),
    .B1(_04718_),
    .C1(net1632),
    .X(_04722_));
 sky130_fd_sc_hd__o211a_1 _09810_ (.A1(net1722),
    .A2(\core.registers[7][22] ),
    .B1(net1617),
    .C1(_04713_),
    .X(_04723_));
 sky130_fd_sc_hd__mux2_1 _09811_ (.A0(\core.registers[4][22] ),
    .A1(\core.registers[5][22] ),
    .S(net1530),
    .X(_04724_));
 sky130_fd_sc_hd__a211o_1 _09812_ (.A1(net1603),
    .A2(_04724_),
    .B1(_04723_),
    .C1(net1577),
    .X(_04725_));
 sky130_fd_sc_hd__o211a_1 _09813_ (.A1(\core.registers[0][22] ),
    .A2(net1530),
    .B1(_04712_),
    .C1(net1604),
    .X(_04726_));
 sky130_fd_sc_hd__mux2_1 _09814_ (.A0(\core.registers[2][22] ),
    .A1(\core.registers[3][22] ),
    .S(net1526),
    .X(_04727_));
 sky130_fd_sc_hd__a211o_1 _09815_ (.A1(net1619),
    .A2(_04727_),
    .B1(_04726_),
    .C1(net1588),
    .X(_04728_));
 sky130_fd_sc_hd__o211a_1 _09816_ (.A1(\core.registers[16][22] ),
    .A2(net1530),
    .B1(_04714_),
    .C1(net1602),
    .X(_04729_));
 sky130_fd_sc_hd__mux2_1 _09817_ (.A0(\core.registers[18][22] ),
    .A1(\core.registers[19][22] ),
    .S(net1530),
    .X(_04730_));
 sky130_fd_sc_hd__a211o_1 _09818_ (.A1(net1618),
    .A2(_04730_),
    .B1(_04729_),
    .C1(net1589),
    .X(_04731_));
 sky130_fd_sc_hd__mux2_1 _09819_ (.A0(\core.registers[22][22] ),
    .A1(\core.registers[23][22] ),
    .S(net1528),
    .X(_04732_));
 sky130_fd_sc_hd__mux2_1 _09820_ (.A0(\core.registers[20][22] ),
    .A1(\core.registers[21][22] ),
    .S(net1526),
    .X(_04733_));
 sky130_fd_sc_hd__mux2_1 _09821_ (.A0(_04732_),
    .A1(_04733_),
    .S(net1602),
    .X(_04734_));
 sky130_fd_sc_hd__o211a_1 _09822_ (.A1(net1578),
    .A2(_04734_),
    .B1(_04731_),
    .C1(net1572),
    .X(_04735_));
 sky130_fd_sc_hd__a311o_1 _09823_ (.A1(net1568),
    .A2(_04725_),
    .A3(_04728_),
    .B1(_04735_),
    .C1(net1636),
    .X(_04736_));
 sky130_fd_sc_hd__a21o_2 _09824_ (.A1(_04722_),
    .A2(_04736_),
    .B1(net1158),
    .X(_04737_));
 sky130_fd_sc_hd__o211ai_4 _09825_ (.A1(net1154),
    .A2(_04703_),
    .B1(_04737_),
    .C1(net1264),
    .Y(_04738_));
 sky130_fd_sc_hd__o21a_1 _09826_ (.A1(net1192),
    .A2(_04738_),
    .B1(net1161),
    .X(_04739_));
 sky130_fd_sc_hd__a21oi_2 _09827_ (.A1(net1744),
    .A2(net1285),
    .B1(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__o22a_1 _09828_ (.A1(net1686),
    .A2(\core.registers[23][22] ),
    .B1(net1401),
    .B2(\core.registers[22][22] ),
    .X(_04741_));
 sky130_fd_sc_hd__or3_1 _09829_ (.A(net1686),
    .B(\core.registers[19][22] ),
    .C(net1448),
    .X(_04742_));
 sky130_fd_sc_hd__o221a_1 _09830_ (.A1(\core.registers[18][22] ),
    .A2(net1332),
    .B1(_04741_),
    .B2(net1436),
    .C1(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__mux4_1 _09831_ (.A0(\core.registers[16][22] ),
    .A1(\core.registers[17][22] ),
    .A2(\core.registers[20][22] ),
    .A3(\core.registers[21][22] ),
    .S0(net1397),
    .S1(net1447),
    .X(_04744_));
 sky130_fd_sc_hd__mux2_1 _09832_ (.A0(_04743_),
    .A1(_04744_),
    .S(net1470),
    .X(_04745_));
 sky130_fd_sc_hd__o22a_1 _09833_ (.A1(net1684),
    .A2(\core.registers[7][22] ),
    .B1(net1397),
    .B2(\core.registers[6][22] ),
    .X(_04746_));
 sky130_fd_sc_hd__or3_1 _09834_ (.A(net1685),
    .B(\core.registers[3][22] ),
    .C(net1447),
    .X(_04747_));
 sky130_fd_sc_hd__o221a_1 _09835_ (.A1(\core.registers[2][22] ),
    .A2(net1332),
    .B1(_04746_),
    .B2(net1435),
    .C1(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__mux4_1 _09836_ (.A0(\core.registers[0][22] ),
    .A1(\core.registers[1][22] ),
    .A2(\core.registers[4][22] ),
    .A3(\core.registers[5][22] ),
    .S0(net1401),
    .S1(net1448),
    .X(_04749_));
 sky130_fd_sc_hd__mux2_1 _09837_ (.A0(_04748_),
    .A1(_04749_),
    .S(net1469),
    .X(_04750_));
 sky130_fd_sc_hd__mux2_1 _09838_ (.A0(_04745_),
    .A1(_04750_),
    .S(net1461),
    .X(_04751_));
 sky130_fd_sc_hd__or2_1 _09839_ (.A(net1490),
    .B(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__mux2_1 _09840_ (.A0(\core.registers[14][22] ),
    .A1(\core.registers[15][22] ),
    .S(net1399),
    .X(_04753_));
 sky130_fd_sc_hd__mux2_1 _09841_ (.A0(\core.registers[12][22] ),
    .A1(\core.registers[13][22] ),
    .S(net1400),
    .X(_04754_));
 sky130_fd_sc_hd__mux2_1 _09842_ (.A0(_04753_),
    .A1(_04754_),
    .S(net1470),
    .X(_04755_));
 sky130_fd_sc_hd__mux2_1 _09843_ (.A0(\core.registers[28][22] ),
    .A1(\core.registers[29][22] ),
    .S(net1399),
    .X(_04756_));
 sky130_fd_sc_hd__a221o_1 _09844_ (.A1(net1686),
    .A2(\core.registers[30][22] ),
    .B1(\core.registers[31][22] ),
    .B2(net1399),
    .C1(net1706),
    .X(_04757_));
 sky130_fd_sc_hd__o21ai_1 _09845_ (.A1(net1870),
    .A2(_04756_),
    .B1(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__nand2_1 _09846_ (.A(net1855),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__o211a_1 _09847_ (.A1(net1861),
    .A2(_04755_),
    .B1(_04759_),
    .C1(net1867),
    .X(_04760_));
 sky130_fd_sc_hd__a221o_1 _09848_ (.A1(net1686),
    .A2(\core.registers[26][22] ),
    .B1(\core.registers[27][22] ),
    .B2(net1399),
    .C1(net1706),
    .X(_04761_));
 sky130_fd_sc_hd__mux2_1 _09849_ (.A0(\core.registers[24][22] ),
    .A1(\core.registers[25][22] ),
    .S(net1399),
    .X(_04762_));
 sky130_fd_sc_hd__o21a_1 _09850_ (.A1(net1870),
    .A2(_04762_),
    .B1(_04761_),
    .X(_04763_));
 sky130_fd_sc_hd__or2_1 _09851_ (.A(\core.registers[9][22] ),
    .B(net1374),
    .X(_04764_));
 sky130_fd_sc_hd__o21a_1 _09852_ (.A1(\core.registers[8][22] ),
    .A2(net1399),
    .B1(net1706),
    .X(_04765_));
 sky130_fd_sc_hd__a22o_1 _09853_ (.A1(net1686),
    .A2(\core.registers[10][22] ),
    .B1(\core.registers[11][22] ),
    .B2(net1399),
    .X(_04766_));
 sky130_fd_sc_hd__a221o_1 _09854_ (.A1(_04764_),
    .A2(_04765_),
    .B1(_04766_),
    .B2(net1870),
    .C1(net1861),
    .X(_04767_));
 sky130_fd_sc_hd__o211a_1 _09855_ (.A1(net1716),
    .A2(_04763_),
    .B1(_04767_),
    .C1(net1715),
    .X(_04768_));
 sky130_fd_sc_hd__o31a_4 _09856_ (.A1(net1486),
    .A2(_04760_),
    .A3(_04768_),
    .B1(_04752_),
    .X(_04769_));
 sky130_fd_sc_hd__a22o_4 _09857_ (.A1(net1069),
    .A2(_04703_),
    .B1(_04769_),
    .B2(net1067),
    .X(_04770_));
 sky130_fd_sc_hd__mux2_8 _09858_ (.A0(net464),
    .A1(_04770_),
    .S(net1276),
    .X(_04771_));
 sky130_fd_sc_hd__and2b_1 _09859_ (.A_N(_04740_),
    .B(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__or2_2 _09860_ (.A(_04740_),
    .B(_04771_),
    .X(_04773_));
 sky130_fd_sc_hd__and2_2 _09861_ (.A(_04740_),
    .B(_04771_),
    .X(_04774_));
 sky130_fd_sc_hd__inv_2 _09862_ (.A(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__nand2_1 _09863_ (.A(_04773_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__inv_2 _09864_ (.A(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__a22o_1 _09865_ (.A1(\core.pipe1_resultRegister[21] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[21] ),
    .X(_04778_));
 sky130_fd_sc_hd__mux2_8 _09866_ (.A0(net120),
    .A1(net155),
    .S(net1805),
    .X(_04779_));
 sky130_fd_sc_hd__o32a_1 _09867_ (.A1(net1673),
    .A2(net1651),
    .A3(_04779_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[21] ),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_2 _09868_ (.A0(\core.pipe1_loadResult[21] ),
    .A1(_04780_),
    .S(net1757),
    .X(_04781_));
 sky130_fd_sc_hd__a21o_4 _09869_ (.A1(net1234),
    .A2(_04781_),
    .B1(net1237),
    .X(_04782_));
 sky130_fd_sc_hd__a21o_1 _09870_ (.A1(net1188),
    .A2(_04782_),
    .B1(_04778_),
    .X(_04783_));
 sky130_fd_sc_hd__or2_1 _09871_ (.A(\core.registers[1][21] ),
    .B(net1494),
    .X(_04784_));
 sky130_fd_sc_hd__or2_1 _09872_ (.A(\core.registers[6][21] ),
    .B(net1517),
    .X(_04785_));
 sky130_fd_sc_hd__or2_1 _09873_ (.A(\core.registers[17][21] ),
    .B(net1494),
    .X(_04786_));
 sky130_fd_sc_hd__or2_1 _09874_ (.A(\core.registers[29][21] ),
    .B(net1493),
    .X(_04787_));
 sky130_fd_sc_hd__o211a_1 _09875_ (.A1(\core.registers[28][21] ),
    .A2(net1508),
    .B1(_04787_),
    .C1(net1735),
    .X(_04788_));
 sky130_fd_sc_hd__a31o_1 _09876_ (.A1(net1839),
    .A2(net1719),
    .A3(\core.registers[30][21] ),
    .B1(net1748),
    .X(_04789_));
 sky130_fd_sc_hd__a31o_1 _09877_ (.A1(net1839),
    .A2(\core.registers[31][21] ),
    .A3(net1507),
    .B1(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__mux2_1 _09878_ (.A0(\core.registers[8][21] ),
    .A1(\core.registers[9][21] ),
    .S(net1506),
    .X(_04791_));
 sky130_fd_sc_hd__mux2_1 _09879_ (.A0(\core.registers[10][21] ),
    .A1(\core.registers[11][21] ),
    .S(net1506),
    .X(_04792_));
 sky130_fd_sc_hd__mux2_1 _09880_ (.A0(\core.registers[24][21] ),
    .A1(\core.registers[25][21] ),
    .S(net1507),
    .X(_04793_));
 sky130_fd_sc_hd__a221o_1 _09881_ (.A1(net1719),
    .A2(\core.registers[26][21] ),
    .B1(\core.registers[27][21] ),
    .B2(net1507),
    .C1(net1735),
    .X(_04794_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(\core.registers[12][21] ),
    .A1(\core.registers[13][21] ),
    .S(net1506),
    .X(_04795_));
 sky130_fd_sc_hd__mux2_1 _09883_ (.A0(\core.registers[14][21] ),
    .A1(\core.registers[15][21] ),
    .S(net1506),
    .X(_04796_));
 sky130_fd_sc_hd__mux2_1 _09884_ (.A0(_04795_),
    .A1(_04796_),
    .S(net1613),
    .X(_04797_));
 sky130_fd_sc_hd__o221a_1 _09885_ (.A1(_04788_),
    .A2(_04790_),
    .B1(_04797_),
    .B2(net1823),
    .C1(net1832),
    .X(_04798_));
 sky130_fd_sc_hd__mux2_1 _09886_ (.A0(_04791_),
    .A1(_04792_),
    .S(net1611),
    .X(_04799_));
 sky130_fd_sc_hd__o21a_1 _09887_ (.A1(net1838),
    .A2(_04793_),
    .B1(_04794_),
    .X(_04800_));
 sky130_fd_sc_hd__mux2_1 _09888_ (.A0(_04799_),
    .A1(_04800_),
    .S(net1823),
    .X(_04801_));
 sky130_fd_sc_hd__a211o_2 _09889_ (.A1(net1744),
    .A2(_04801_),
    .B1(_04798_),
    .C1(net1631),
    .X(_04802_));
 sky130_fd_sc_hd__o211a_1 _09890_ (.A1(net1721),
    .A2(\core.registers[7][21] ),
    .B1(net1615),
    .C1(_04785_),
    .X(_04803_));
 sky130_fd_sc_hd__mux2_1 _09891_ (.A0(\core.registers[4][21] ),
    .A1(\core.registers[5][21] ),
    .S(net1517),
    .X(_04804_));
 sky130_fd_sc_hd__a211o_1 _09892_ (.A1(net1599),
    .A2(_04804_),
    .B1(_04803_),
    .C1(net1575),
    .X(_04805_));
 sky130_fd_sc_hd__o211a_1 _09893_ (.A1(\core.registers[0][21] ),
    .A2(net1517),
    .B1(_04784_),
    .C1(net1599),
    .X(_04806_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(\core.registers[2][21] ),
    .A1(\core.registers[3][21] ),
    .S(net1517),
    .X(_04807_));
 sky130_fd_sc_hd__a211o_1 _09895_ (.A1(net1615),
    .A2(_04807_),
    .B1(_04806_),
    .C1(net1586),
    .X(_04808_));
 sky130_fd_sc_hd__o211a_1 _09896_ (.A1(\core.registers[16][21] ),
    .A2(net1515),
    .B1(_04786_),
    .C1(net1600),
    .X(_04809_));
 sky130_fd_sc_hd__mux2_1 _09897_ (.A0(\core.registers[18][21] ),
    .A1(\core.registers[19][21] ),
    .S(net1515),
    .X(_04810_));
 sky130_fd_sc_hd__a211o_1 _09898_ (.A1(net1614),
    .A2(_04810_),
    .B1(_04809_),
    .C1(net1586),
    .X(_04811_));
 sky130_fd_sc_hd__mux2_1 _09899_ (.A0(\core.registers[22][21] ),
    .A1(\core.registers[23][21] ),
    .S(net1515),
    .X(_04812_));
 sky130_fd_sc_hd__mux2_1 _09900_ (.A0(\core.registers[20][21] ),
    .A1(\core.registers[21][21] ),
    .S(net1515),
    .X(_04813_));
 sky130_fd_sc_hd__mux2_1 _09901_ (.A0(_04812_),
    .A1(_04813_),
    .S(net1600),
    .X(_04814_));
 sky130_fd_sc_hd__o211a_1 _09902_ (.A1(net1575),
    .A2(_04814_),
    .B1(_04811_),
    .C1(net1571),
    .X(_04815_));
 sky130_fd_sc_hd__a311o_1 _09903_ (.A1(net1567),
    .A2(_04805_),
    .A3(_04808_),
    .B1(_04815_),
    .C1(net1635),
    .X(_04816_));
 sky130_fd_sc_hd__a21o_2 _09904_ (.A1(_04802_),
    .A2(_04816_),
    .B1(net1157),
    .X(_04817_));
 sky130_fd_sc_hd__o211ai_4 _09905_ (.A1(net1153),
    .A2(net1144),
    .B1(_04817_),
    .C1(net1263),
    .Y(_04818_));
 sky130_fd_sc_hd__o21a_1 _09906_ (.A1(net1192),
    .A2(_04818_),
    .B1(net1161),
    .X(_04819_));
 sky130_fd_sc_hd__a21oi_2 _09907_ (.A1(net1738),
    .A2(net1285),
    .B1(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__o22a_1 _09908_ (.A1(net1682),
    .A2(\core.registers[23][21] ),
    .B1(net1389),
    .B2(\core.registers[22][21] ),
    .X(_04821_));
 sky130_fd_sc_hd__or3_1 _09909_ (.A(net1682),
    .B(\core.registers[19][21] ),
    .C(net1445),
    .X(_04822_));
 sky130_fd_sc_hd__o221a_1 _09910_ (.A1(\core.registers[18][21] ),
    .A2(net1331),
    .B1(_04821_),
    .B2(net1434),
    .C1(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__mux4_1 _09911_ (.A0(\core.registers[16][21] ),
    .A1(\core.registers[17][21] ),
    .A2(\core.registers[20][21] ),
    .A3(\core.registers[21][21] ),
    .S0(net1388),
    .S1(net1445),
    .X(_04824_));
 sky130_fd_sc_hd__mux2_1 _09912_ (.A0(_04823_),
    .A1(_04824_),
    .S(net1467),
    .X(_04825_));
 sky130_fd_sc_hd__o22a_1 _09913_ (.A1(net1682),
    .A2(\core.registers[7][21] ),
    .B1(net1390),
    .B2(\core.registers[6][21] ),
    .X(_04826_));
 sky130_fd_sc_hd__or3_1 _09914_ (.A(net1682),
    .B(\core.registers[3][21] ),
    .C(net1445),
    .X(_04827_));
 sky130_fd_sc_hd__o221a_1 _09915_ (.A1(\core.registers[2][21] ),
    .A2(net1331),
    .B1(_04826_),
    .B2(net1434),
    .C1(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__mux4_1 _09916_ (.A0(\core.registers[0][21] ),
    .A1(\core.registers[1][21] ),
    .A2(\core.registers[4][21] ),
    .A3(\core.registers[5][21] ),
    .S0(net1390),
    .S1(net1446),
    .X(_04829_));
 sky130_fd_sc_hd__mux2_1 _09917_ (.A0(_04828_),
    .A1(_04829_),
    .S(net1467),
    .X(_04830_));
 sky130_fd_sc_hd__mux2_1 _09918_ (.A0(_04825_),
    .A1(_04830_),
    .S(net1460),
    .X(_04831_));
 sky130_fd_sc_hd__a221o_1 _09919_ (.A1(net1677),
    .A2(\core.registers[26][21] ),
    .B1(\core.registers[27][21] ),
    .B2(net1382),
    .C1(net1705),
    .X(_04832_));
 sky130_fd_sc_hd__mux2_1 _09920_ (.A0(\core.registers[24][21] ),
    .A1(\core.registers[25][21] ),
    .S(net1382),
    .X(_04833_));
 sky130_fd_sc_hd__o21ai_1 _09921_ (.A1(net1869),
    .A2(_04833_),
    .B1(_04832_),
    .Y(_04834_));
 sky130_fd_sc_hd__a221o_1 _09922_ (.A1(net1677),
    .A2(\core.registers[10][21] ),
    .B1(\core.registers[11][21] ),
    .B2(net1381),
    .C1(net1704),
    .X(_04835_));
 sky130_fd_sc_hd__a21o_1 _09923_ (.A1(\core.registers[8][21] ),
    .A2(net1373),
    .B1(net1869),
    .X(_04836_));
 sky130_fd_sc_hd__a21o_1 _09924_ (.A1(\core.registers[9][21] ),
    .A2(net1381),
    .B1(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__a21oi_1 _09925_ (.A1(_04835_),
    .A2(_04837_),
    .B1(net1853),
    .Y(_04838_));
 sky130_fd_sc_hd__a211o_1 _09926_ (.A1(net1854),
    .A2(_04834_),
    .B1(_04838_),
    .C1(net1862),
    .X(_04839_));
 sky130_fd_sc_hd__mux2_1 _09927_ (.A0(\core.registers[12][21] ),
    .A1(\core.registers[13][21] ),
    .S(net1381),
    .X(_04840_));
 sky130_fd_sc_hd__mux2_1 _09928_ (.A0(\core.registers[14][21] ),
    .A1(\core.registers[15][21] ),
    .S(net1381),
    .X(_04841_));
 sky130_fd_sc_hd__mux2_1 _09929_ (.A0(_04840_),
    .A1(_04841_),
    .S(net1480),
    .X(_04842_));
 sky130_fd_sc_hd__a221o_1 _09930_ (.A1(net1678),
    .A2(\core.registers[30][21] ),
    .B1(\core.registers[31][21] ),
    .B2(net1382),
    .C1(net1704),
    .X(_04843_));
 sky130_fd_sc_hd__mux2_1 _09931_ (.A0(\core.registers[28][21] ),
    .A1(\core.registers[29][21] ),
    .S(net1382),
    .X(_04844_));
 sky130_fd_sc_hd__o21a_1 _09932_ (.A1(net1868),
    .A2(_04844_),
    .B1(_04843_),
    .X(_04845_));
 sky130_fd_sc_hd__mux2_1 _09933_ (.A0(_04842_),
    .A1(_04845_),
    .S(net1853),
    .X(_04846_));
 sky130_fd_sc_hd__a21oi_2 _09934_ (.A1(net1862),
    .A2(_04846_),
    .B1(net1484),
    .Y(_04847_));
 sky130_fd_sc_hd__o2bb2a_2 _09935_ (.A1_N(_04839_),
    .A2_N(_04847_),
    .B1(net1490),
    .B2(_04831_),
    .X(_04848_));
 sky130_fd_sc_hd__a22o_2 _09936_ (.A1(net1068),
    .A2(net1144),
    .B1(_04848_),
    .B2(net1065),
    .X(_04849_));
 sky130_fd_sc_hd__mux2_8 _09937_ (.A0(net463),
    .A1(_04849_),
    .S(net1278),
    .X(_04850_));
 sky130_fd_sc_hd__or2_1 _09938_ (.A(_04820_),
    .B(_04850_),
    .X(_04851_));
 sky130_fd_sc_hd__nand2_2 _09939_ (.A(_04820_),
    .B(_04850_),
    .Y(_04852_));
 sky130_fd_sc_hd__inv_2 _09940_ (.A(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__and2_4 _09941_ (.A(_04851_),
    .B(_04852_),
    .X(_04854_));
 sky130_fd_sc_hd__a22o_1 _09942_ (.A1(\core.pipe1_resultRegister[20] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[20] ),
    .X(_04855_));
 sky130_fd_sc_hd__mux2_8 _09943_ (.A0(net119),
    .A1(net154),
    .S(net1805),
    .X(_04856_));
 sky130_fd_sc_hd__o32a_1 _09944_ (.A1(net1673),
    .A2(net1651),
    .A3(_04856_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[20] ),
    .X(_04857_));
 sky130_fd_sc_hd__mux2_2 _09945_ (.A0(\core.pipe1_loadResult[20] ),
    .A1(_04857_),
    .S(net1757),
    .X(_04858_));
 sky130_fd_sc_hd__a21o_4 _09946_ (.A1(net1235),
    .A2(_04858_),
    .B1(net1237),
    .X(_04859_));
 sky130_fd_sc_hd__a21o_4 _09947_ (.A1(net1188),
    .A2(_04859_),
    .B1(_04855_),
    .X(_04860_));
 sky130_fd_sc_hd__or2_1 _09948_ (.A(\core.registers[1][20] ),
    .B(net1494),
    .X(_04861_));
 sky130_fd_sc_hd__or2_1 _09949_ (.A(\core.registers[6][20] ),
    .B(net1520),
    .X(_04862_));
 sky130_fd_sc_hd__or2_1 _09950_ (.A(\core.registers[17][20] ),
    .B(net1495),
    .X(_04863_));
 sky130_fd_sc_hd__or2_1 _09951_ (.A(\core.registers[28][20] ),
    .B(net1505),
    .X(_04864_));
 sky130_fd_sc_hd__o211a_1 _09952_ (.A1(\core.registers[29][20] ),
    .A2(net1493),
    .B1(_04864_),
    .C1(net1735),
    .X(_04865_));
 sky130_fd_sc_hd__a31o_1 _09953_ (.A1(net1838),
    .A2(net1719),
    .A3(\core.registers[30][20] ),
    .B1(net1748),
    .X(_04866_));
 sky130_fd_sc_hd__a31o_1 _09954_ (.A1(net1838),
    .A2(\core.registers[31][20] ),
    .A3(net1505),
    .B1(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__mux2_1 _09955_ (.A0(\core.registers[8][20] ),
    .A1(\core.registers[9][20] ),
    .S(net1504),
    .X(_04868_));
 sky130_fd_sc_hd__mux2_1 _09956_ (.A0(\core.registers[10][20] ),
    .A1(\core.registers[11][20] ),
    .S(net1504),
    .X(_04869_));
 sky130_fd_sc_hd__mux2_1 _09957_ (.A0(\core.registers[24][20] ),
    .A1(\core.registers[25][20] ),
    .S(net1510),
    .X(_04870_));
 sky130_fd_sc_hd__a221o_1 _09958_ (.A1(net1719),
    .A2(\core.registers[26][20] ),
    .B1(\core.registers[27][20] ),
    .B2(net1509),
    .C1(net1735),
    .X(_04871_));
 sky130_fd_sc_hd__mux2_1 _09959_ (.A0(\core.registers[12][20] ),
    .A1(\core.registers[13][20] ),
    .S(net1504),
    .X(_04872_));
 sky130_fd_sc_hd__mux2_1 _09960_ (.A0(\core.registers[14][20] ),
    .A1(\core.registers[15][20] ),
    .S(net1504),
    .X(_04873_));
 sky130_fd_sc_hd__mux2_1 _09961_ (.A0(_04872_),
    .A1(_04873_),
    .S(net1611),
    .X(_04874_));
 sky130_fd_sc_hd__o221a_1 _09962_ (.A1(_04865_),
    .A2(_04867_),
    .B1(_04874_),
    .B2(net1823),
    .C1(net1832),
    .X(_04875_));
 sky130_fd_sc_hd__mux2_1 _09963_ (.A0(_04868_),
    .A1(_04869_),
    .S(net1611),
    .X(_04876_));
 sky130_fd_sc_hd__o21a_1 _09964_ (.A1(net1838),
    .A2(_04870_),
    .B1(_04871_),
    .X(_04877_));
 sky130_fd_sc_hd__mux2_1 _09965_ (.A0(_04876_),
    .A1(_04877_),
    .S(net1823),
    .X(_04878_));
 sky130_fd_sc_hd__a211o_2 _09966_ (.A1(net1744),
    .A2(_04878_),
    .B1(_04875_),
    .C1(net1631),
    .X(_04879_));
 sky130_fd_sc_hd__o211a_1 _09967_ (.A1(net1721),
    .A2(\core.registers[7][20] ),
    .B1(net1616),
    .C1(_04862_),
    .X(_04880_));
 sky130_fd_sc_hd__mux2_1 _09968_ (.A0(\core.registers[4][20] ),
    .A1(\core.registers[5][20] ),
    .S(net1515),
    .X(_04881_));
 sky130_fd_sc_hd__a211o_1 _09969_ (.A1(net1600),
    .A2(_04881_),
    .B1(_04880_),
    .C1(net1576),
    .X(_04882_));
 sky130_fd_sc_hd__o211a_1 _09970_ (.A1(\core.registers[0][20] ),
    .A2(net1515),
    .B1(_04861_),
    .C1(net1600),
    .X(_04883_));
 sky130_fd_sc_hd__mux2_1 _09971_ (.A0(\core.registers[2][20] ),
    .A1(\core.registers[3][20] ),
    .S(net1515),
    .X(_04884_));
 sky130_fd_sc_hd__a211o_1 _09972_ (.A1(net1614),
    .A2(_04884_),
    .B1(_04883_),
    .C1(net1586),
    .X(_04885_));
 sky130_fd_sc_hd__o211a_1 _09973_ (.A1(\core.registers[16][20] ),
    .A2(net1520),
    .B1(_04863_),
    .C1(net1601),
    .X(_04886_));
 sky130_fd_sc_hd__mux2_1 _09974_ (.A0(\core.registers[18][20] ),
    .A1(\core.registers[19][20] ),
    .S(net1516),
    .X(_04887_));
 sky130_fd_sc_hd__a211o_1 _09975_ (.A1(net1614),
    .A2(_04887_),
    .B1(_04886_),
    .C1(net1586),
    .X(_04888_));
 sky130_fd_sc_hd__mux2_1 _09976_ (.A0(\core.registers[22][20] ),
    .A1(\core.registers[23][20] ),
    .S(net1516),
    .X(_04889_));
 sky130_fd_sc_hd__mux2_1 _09977_ (.A0(\core.registers[20][20] ),
    .A1(\core.registers[21][20] ),
    .S(net1512),
    .X(_04890_));
 sky130_fd_sc_hd__mux2_1 _09978_ (.A0(_04889_),
    .A1(_04890_),
    .S(net1598),
    .X(_04891_));
 sky130_fd_sc_hd__o211a_1 _09979_ (.A1(net1575),
    .A2(_04891_),
    .B1(_04888_),
    .C1(net1571),
    .X(_04892_));
 sky130_fd_sc_hd__a311o_1 _09980_ (.A1(net1567),
    .A2(_04882_),
    .A3(_04885_),
    .B1(_04892_),
    .C1(net1635),
    .X(_04893_));
 sky130_fd_sc_hd__a21o_2 _09981_ (.A1(_04879_),
    .A2(_04893_),
    .B1(net1157),
    .X(_04894_));
 sky130_fd_sc_hd__o211ai_4 _09982_ (.A1(net1153),
    .A2(net1138),
    .B1(_04894_),
    .C1(net1263),
    .Y(_04895_));
 sky130_fd_sc_hd__o21a_1 _09983_ (.A1(net1192),
    .A2(_04895_),
    .B1(net1161),
    .X(_04896_));
 sky130_fd_sc_hd__a21oi_2 _09984_ (.A1(net1721),
    .A2(net1285),
    .B1(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__o22a_1 _09985_ (.A1(net1677),
    .A2(\core.registers[23][20] ),
    .B1(net1389),
    .B2(\core.registers[22][20] ),
    .X(_04898_));
 sky130_fd_sc_hd__or3_1 _09986_ (.A(net1677),
    .B(\core.registers[19][20] ),
    .C(net1444),
    .X(_04899_));
 sky130_fd_sc_hd__o221a_1 _09987_ (.A1(\core.registers[18][20] ),
    .A2(net1331),
    .B1(_04898_),
    .B2(net1431),
    .C1(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__mux4_1 _09988_ (.A0(\core.registers[16][20] ),
    .A1(\core.registers[17][20] ),
    .A2(\core.registers[20][20] ),
    .A3(\core.registers[21][20] ),
    .S0(net1385),
    .S1(net1442),
    .X(_04901_));
 sky130_fd_sc_hd__mux2_1 _09989_ (.A0(_04900_),
    .A1(_04901_),
    .S(net1465),
    .X(_04902_));
 sky130_fd_sc_hd__o22a_1 _09990_ (.A1(net1683),
    .A2(\core.registers[7][20] ),
    .B1(net1392),
    .B2(\core.registers[6][20] ),
    .X(_04903_));
 sky130_fd_sc_hd__or3_1 _09991_ (.A(net1682),
    .B(\core.registers[3][20] ),
    .C(net1445),
    .X(_04904_));
 sky130_fd_sc_hd__o221a_1 _09992_ (.A1(\core.registers[2][20] ),
    .A2(net1331),
    .B1(_04903_),
    .B2(net1434),
    .C1(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__mux4_1 _09993_ (.A0(\core.registers[0][20] ),
    .A1(\core.registers[1][20] ),
    .A2(\core.registers[4][20] ),
    .A3(\core.registers[5][20] ),
    .S0(net1389),
    .S1(net1445),
    .X(_04906_));
 sky130_fd_sc_hd__mux2_1 _09994_ (.A0(_04905_),
    .A1(_04906_),
    .S(net1467),
    .X(_04907_));
 sky130_fd_sc_hd__mux2_1 _09995_ (.A0(_04902_),
    .A1(_04907_),
    .S(net1460),
    .X(_04908_));
 sky130_fd_sc_hd__mux2_1 _09996_ (.A0(\core.registers[24][20] ),
    .A1(\core.registers[25][20] ),
    .S(net1383),
    .X(_04909_));
 sky130_fd_sc_hd__a221o_1 _09997_ (.A1(net1679),
    .A2(\core.registers[26][20] ),
    .B1(\core.registers[27][20] ),
    .B2(net1383),
    .C1(net1704),
    .X(_04910_));
 sky130_fd_sc_hd__o21ai_1 _09998_ (.A1(net1869),
    .A2(_04909_),
    .B1(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__a221o_1 _09999_ (.A1(net1678),
    .A2(\core.registers[10][20] ),
    .B1(\core.registers[11][20] ),
    .B2(net1379),
    .C1(net1704),
    .X(_04912_));
 sky130_fd_sc_hd__a21o_1 _10000_ (.A1(\core.registers[8][20] ),
    .A2(net1373),
    .B1(net1868),
    .X(_04913_));
 sky130_fd_sc_hd__a21o_1 _10001_ (.A1(\core.registers[9][20] ),
    .A2(net1379),
    .B1(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__a21oi_1 _10002_ (.A1(_04912_),
    .A2(_04914_),
    .B1(net1853),
    .Y(_04915_));
 sky130_fd_sc_hd__a211o_1 _10003_ (.A1(net1854),
    .A2(_04911_),
    .B1(_04915_),
    .C1(net1862),
    .X(_04916_));
 sky130_fd_sc_hd__mux2_1 _10004_ (.A0(\core.registers[12][20] ),
    .A1(\core.registers[13][20] ),
    .S(net1379),
    .X(_04917_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(\core.registers[14][20] ),
    .A1(\core.registers[15][20] ),
    .S(net1379),
    .X(_04918_));
 sky130_fd_sc_hd__mux2_1 _10006_ (.A0(_04917_),
    .A1(_04918_),
    .S(net1480),
    .X(_04919_));
 sky130_fd_sc_hd__a221o_1 _10007_ (.A1(net1678),
    .A2(\core.registers[30][20] ),
    .B1(\core.registers[31][20] ),
    .B2(net1380),
    .C1(net1704),
    .X(_04920_));
 sky130_fd_sc_hd__mux2_1 _10008_ (.A0(\core.registers[28][20] ),
    .A1(\core.registers[29][20] ),
    .S(net1380),
    .X(_04921_));
 sky130_fd_sc_hd__o21a_1 _10009_ (.A1(net1868),
    .A2(_04921_),
    .B1(_04920_),
    .X(_04922_));
 sky130_fd_sc_hd__mux2_1 _10010_ (.A0(_04919_),
    .A1(_04922_),
    .S(net1853),
    .X(_04923_));
 sky130_fd_sc_hd__a21oi_1 _10011_ (.A1(net1862),
    .A2(_04923_),
    .B1(net1484),
    .Y(_04924_));
 sky130_fd_sc_hd__o2bb2a_2 _10012_ (.A1_N(_04916_),
    .A2_N(_04924_),
    .B1(net1489),
    .B2(_04908_),
    .X(_04925_));
 sky130_fd_sc_hd__a22o_4 _10013_ (.A1(net1068),
    .A2(net1139),
    .B1(_04925_),
    .B2(net1065),
    .X(_04926_));
 sky130_fd_sc_hd__mux2_8 _10014_ (.A0(net462),
    .A1(_04926_),
    .S(net1278),
    .X(_04927_));
 sky130_fd_sc_hd__nand2b_2 _10015_ (.A_N(_04897_),
    .B(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2b_1 _10016_ (.A_N(_04820_),
    .B(_04850_),
    .Y(_04929_));
 sky130_fd_sc_hd__o21ai_2 _10017_ (.A1(_04854_),
    .A2(_04928_),
    .B1(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__inv_2 _10018_ (.A(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__a221o_1 _10019_ (.A1(\core.pipe1_resultRegister[12] ),
    .A2(_04498_),
    .B1(net1270),
    .B2(\core.pipe1_csrData[12] ),
    .C1(net1187),
    .X(_04932_));
 sky130_fd_sc_hd__nor2_2 _10020_ (.A(net1810),
    .B(_04490_),
    .Y(_04933_));
 sky130_fd_sc_hd__a21oi_1 _10021_ (.A1(_04525_),
    .A2(_04548_),
    .B1(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__a21o_4 _10022_ (.A1(_04525_),
    .A2(_04548_),
    .B1(_04933_),
    .X(_04935_));
 sky130_fd_sc_hd__o21ai_2 _10023_ (.A1(net1808),
    .A2(_04935_),
    .B1(net1236),
    .Y(_04936_));
 sky130_fd_sc_hd__and2_4 _10024_ (.A(_04571_),
    .B(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__mux2_8 _10025_ (.A0(net110),
    .A1(net145),
    .S(net1805),
    .X(_04938_));
 sky130_fd_sc_hd__o32a_1 _10026_ (.A1(net1674),
    .A2(net1653),
    .A3(_04938_),
    .B1(net1659),
    .B2(\coreWBInterface.readDataBuffered[12] ),
    .X(_04939_));
 sky130_fd_sc_hd__mux2_1 _10027_ (.A0(\core.pipe1_loadResult[12] ),
    .A1(_04939_),
    .S(net1759),
    .X(_04940_));
 sky130_fd_sc_hd__or3b_2 _10028_ (.A(net1807),
    .B(_04935_),
    .C_N(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__nor2_1 _10029_ (.A(net1806),
    .B(_04552_),
    .Y(_04942_));
 sky130_fd_sc_hd__or2_1 _10030_ (.A(net1806),
    .B(_04552_),
    .X(_04943_));
 sky130_fd_sc_hd__a211oi_4 _10031_ (.A1(_04524_),
    .A2(_04548_),
    .B1(_04557_),
    .C1(_04942_),
    .Y(_04944_));
 sky130_fd_sc_hd__nand2b_4 _10032_ (.A_N(_04944_),
    .B(net1237),
    .Y(_04945_));
 sky130_fd_sc_hd__nand2_1 _10033_ (.A(_04858_),
    .B(_04944_),
    .Y(_04946_));
 sky130_fd_sc_hd__a21o_1 _10034_ (.A1(_04945_),
    .A2(_04946_),
    .B1(_04551_),
    .X(_04947_));
 sky130_fd_sc_hd__a21oi_4 _10035_ (.A1(_04557_),
    .A2(net1236),
    .B1(_04571_),
    .Y(_04948_));
 sky130_fd_sc_hd__mux2_2 _10036_ (.A0(_04550_),
    .A1(_04934_),
    .S(net1808),
    .X(_04949_));
 sky130_fd_sc_hd__nand2b_4 _10037_ (.A_N(net1233),
    .B(net1237),
    .Y(_04950_));
 sky130_fd_sc_hd__mux2_8 _10038_ (.A0(net127),
    .A1(net163),
    .S(net1805),
    .X(_04951_));
 sky130_fd_sc_hd__o32a_1 _10039_ (.A1(net1675),
    .A2(net1661),
    .A3(_04951_),
    .B1(net1658),
    .B2(\coreWBInterface.readDataBuffered[28] ),
    .X(_04952_));
 sky130_fd_sc_hd__mux2_2 _10040_ (.A0(\core.pipe1_loadResult[28] ),
    .A1(_04952_),
    .S(net1758),
    .X(_04953_));
 sky130_fd_sc_hd__nand2_1 _10041_ (.A(net1233),
    .B(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__a21o_1 _10042_ (.A1(_04950_),
    .A2(_04954_),
    .B1(_04582_),
    .X(_04955_));
 sky130_fd_sc_hd__a32o_2 _10043_ (.A1(_04947_),
    .A2(_04948_),
    .A3(_04955_),
    .B1(_04941_),
    .B2(_04937_),
    .X(_04956_));
 sky130_fd_sc_hd__nand2_1 _10044_ (.A(net1190),
    .B(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__a22o_2 _10045_ (.A1(\core.pipe1_resultRegister[12] ),
    .A2(net1271),
    .B1(_04932_),
    .B2(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__mux2_1 _10046_ (.A0(\core.registers[14][12] ),
    .A1(\core.registers[15][12] ),
    .S(net1531),
    .X(_04959_));
 sky130_fd_sc_hd__mux2_1 _10047_ (.A0(\core.registers[12][12] ),
    .A1(\core.registers[13][12] ),
    .S(net1531),
    .X(_04960_));
 sky130_fd_sc_hd__mux2_1 _10048_ (.A0(_04959_),
    .A1(_04960_),
    .S(net1602),
    .X(_04961_));
 sky130_fd_sc_hd__mux2_1 _10049_ (.A0(\core.registers[28][12] ),
    .A1(\core.registers[29][12] ),
    .S(net1536),
    .X(_04962_));
 sky130_fd_sc_hd__a221o_1 _10050_ (.A1(net1727),
    .A2(\core.registers[30][12] ),
    .B1(\core.registers[31][12] ),
    .B2(net1536),
    .C1(net1743),
    .X(_04963_));
 sky130_fd_sc_hd__o21a_1 _10051_ (.A1(net1848),
    .A2(_04962_),
    .B1(_04963_),
    .X(_04964_));
 sky130_fd_sc_hd__mux2_1 _10052_ (.A0(\core.registers[8][12] ),
    .A1(\core.registers[9][12] ),
    .S(net1536),
    .X(_04965_));
 sky130_fd_sc_hd__mux2_1 _10053_ (.A0(\core.registers[10][12] ),
    .A1(\core.registers[11][12] ),
    .S(net1529),
    .X(_04966_));
 sky130_fd_sc_hd__mux2_1 _10054_ (.A0(_04965_),
    .A1(_04966_),
    .S(net1619),
    .X(_04967_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(\core.registers[24][12] ),
    .A1(\core.registers[25][12] ),
    .S(net1529),
    .X(_04968_));
 sky130_fd_sc_hd__a22o_1 _10056_ (.A1(net1723),
    .A2(\core.registers[26][12] ),
    .B1(\core.registers[27][12] ),
    .B2(net1529),
    .X(_04969_));
 sky130_fd_sc_hd__mux2_1 _10057_ (.A0(_04968_),
    .A1(_04969_),
    .S(net1842),
    .X(_04970_));
 sky130_fd_sc_hd__mux4_2 _10058_ (.A0(_04961_),
    .A1(_04964_),
    .A2(_04967_),
    .A3(_04970_),
    .S0(net1825),
    .S1(net1745),
    .X(_04971_));
 sky130_fd_sc_hd__and3_1 _10059_ (.A(net1852),
    .B(\core.registers[5][12] ),
    .C(net1662),
    .X(_04972_));
 sky130_fd_sc_hd__a21o_1 _10060_ (.A1(\core.registers[4][12] ),
    .A2(net1496),
    .B1(net1577),
    .X(_04973_));
 sky130_fd_sc_hd__o31a_1 _10061_ (.A1(\core.registers[1][12] ),
    .A2(net1588),
    .A3(net1496),
    .B1(net1602),
    .X(_04974_));
 sky130_fd_sc_hd__o221a_1 _10062_ (.A1(\core.registers[0][12] ),
    .A2(net1341),
    .B1(_04972_),
    .B2(_04973_),
    .C1(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__o22a_1 _10063_ (.A1(net1723),
    .A2(\core.registers[7][12] ),
    .B1(net1531),
    .B2(\core.registers[6][12] ),
    .X(_04976_));
 sky130_fd_sc_hd__o31a_1 _10064_ (.A1(net1723),
    .A2(\core.registers[3][12] ),
    .A3(net1588),
    .B1(net1618),
    .X(_04977_));
 sky130_fd_sc_hd__o221a_1 _10065_ (.A1(\core.registers[2][12] ),
    .A2(net1341),
    .B1(_04976_),
    .B2(net1577),
    .C1(_04977_),
    .X(_04978_));
 sky130_fd_sc_hd__and3_1 _10066_ (.A(net1852),
    .B(\core.registers[21][12] ),
    .C(net1662),
    .X(_04979_));
 sky130_fd_sc_hd__a21o_1 _10067_ (.A1(\core.registers[20][12] ),
    .A2(net1498),
    .B1(net1577),
    .X(_04980_));
 sky130_fd_sc_hd__o31a_1 _10068_ (.A1(\core.registers[17][12] ),
    .A2(net1588),
    .A3(net1498),
    .B1(net1602),
    .X(_04981_));
 sky130_fd_sc_hd__o221a_1 _10069_ (.A1(\core.registers[16][12] ),
    .A2(net1341),
    .B1(_04979_),
    .B2(_04980_),
    .C1(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__o22a_1 _10070_ (.A1(net1723),
    .A2(\core.registers[23][12] ),
    .B1(net1530),
    .B2(\core.registers[22][12] ),
    .X(_04983_));
 sky130_fd_sc_hd__o31a_1 _10071_ (.A1(net1723),
    .A2(\core.registers[19][12] ),
    .A3(net1588),
    .B1(net1618),
    .X(_04984_));
 sky130_fd_sc_hd__o221a_1 _10072_ (.A1(\core.registers[18][12] ),
    .A2(net1341),
    .B1(_04983_),
    .B2(net1577),
    .C1(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__o31a_1 _10073_ (.A1(net1568),
    .A2(_04982_),
    .A3(_04985_),
    .B1(net1632),
    .X(_04986_));
 sky130_fd_sc_hd__o31a_1 _10074_ (.A1(net1572),
    .A2(_04975_),
    .A3(_04978_),
    .B1(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__a211o_2 _10075_ (.A1(net1636),
    .A2(_04971_),
    .B1(_04987_),
    .C1(net1158),
    .X(_04988_));
 sky130_fd_sc_hd__o211a_2 _10076_ (.A1(net1154),
    .A2(net990),
    .B1(_04988_),
    .C1(net1264),
    .X(_04989_));
 sky130_fd_sc_hd__nand2_1 _10077_ (.A(_04484_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__o2bb2a_1 _10078_ (.A1_N(net1162),
    .A2_N(_04990_),
    .B1(net1881),
    .B2(net1282),
    .X(_04991_));
 sky130_fd_sc_hd__or2_1 _10079_ (.A(\core.registers[24][12] ),
    .B(net1400),
    .X(_04992_));
 sky130_fd_sc_hd__o21a_1 _10080_ (.A1(\core.registers[25][12] ),
    .A2(net1374),
    .B1(net1706),
    .X(_04993_));
 sky130_fd_sc_hd__a22o_1 _10081_ (.A1(net1686),
    .A2(\core.registers[26][12] ),
    .B1(\core.registers[27][12] ),
    .B2(net1400),
    .X(_04994_));
 sky130_fd_sc_hd__a221o_1 _10082_ (.A1(_04992_),
    .A2(_04993_),
    .B1(_04994_),
    .B2(net1870),
    .C1(net1716),
    .X(_04995_));
 sky130_fd_sc_hd__a221o_1 _10083_ (.A1(net1686),
    .A2(\core.registers[10][12] ),
    .B1(\core.registers[11][12] ),
    .B2(net1400),
    .C1(net1707),
    .X(_04996_));
 sky130_fd_sc_hd__a21o_1 _10084_ (.A1(\core.registers[8][12] ),
    .A2(net1377),
    .B1(net1872),
    .X(_04997_));
 sky130_fd_sc_hd__a21o_1 _10085_ (.A1(\core.registers[9][12] ),
    .A2(net1405),
    .B1(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__a21o_1 _10086_ (.A1(_04996_),
    .A2(_04998_),
    .B1(net1856),
    .X(_04999_));
 sky130_fd_sc_hd__a21o_1 _10087_ (.A1(_04995_),
    .A2(_04999_),
    .B1(net1867),
    .X(_05000_));
 sky130_fd_sc_hd__a221o_1 _10088_ (.A1(net1690),
    .A2(\core.registers[30][12] ),
    .B1(\core.registers[31][12] ),
    .B2(net1405),
    .C1(net1707),
    .X(_05001_));
 sky130_fd_sc_hd__mux2_1 _10089_ (.A0(\core.registers[28][12] ),
    .A1(\core.registers[29][12] ),
    .S(net1405),
    .X(_05002_));
 sky130_fd_sc_hd__o21a_1 _10090_ (.A1(net1872),
    .A2(_05002_),
    .B1(_05001_),
    .X(_05003_));
 sky130_fd_sc_hd__mux2_1 _10091_ (.A0(\core.registers[12][12] ),
    .A1(\core.registers[13][12] ),
    .S(net1401),
    .X(_05004_));
 sky130_fd_sc_hd__mux2_1 _10092_ (.A0(\core.registers[14][12] ),
    .A1(\core.registers[15][12] ),
    .S(net1401),
    .X(_05005_));
 sky130_fd_sc_hd__mux2_1 _10093_ (.A0(_05004_),
    .A1(_05005_),
    .S(net1483),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _10094_ (.A0(_05003_),
    .A1(_05006_),
    .S(net1716),
    .X(_05007_));
 sky130_fd_sc_hd__o21a_1 _10095_ (.A1(net1715),
    .A2(_05007_),
    .B1(net1492),
    .X(_05008_));
 sky130_fd_sc_hd__o22a_1 _10096_ (.A1(net1687),
    .A2(\core.registers[7][12] ),
    .B1(net1401),
    .B2(\core.registers[6][12] ),
    .X(_05009_));
 sky130_fd_sc_hd__or3_1 _10097_ (.A(net1687),
    .B(\core.registers[3][12] ),
    .C(net1448),
    .X(_05010_));
 sky130_fd_sc_hd__o221a_1 _10098_ (.A1(\core.registers[2][12] ),
    .A2(net1332),
    .B1(_05009_),
    .B2(net1436),
    .C1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__mux4_1 _10099_ (.A0(\core.registers[0][12] ),
    .A1(\core.registers[1][12] ),
    .A2(\core.registers[4][12] ),
    .A3(\core.registers[5][12] ),
    .S0(net1401),
    .S1(net1449),
    .X(_05012_));
 sky130_fd_sc_hd__mux2_1 _10100_ (.A0(_05011_),
    .A1(_05012_),
    .S(net1470),
    .X(_05013_));
 sky130_fd_sc_hd__or2_1 _10101_ (.A(net1464),
    .B(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__o22a_1 _10102_ (.A1(net1687),
    .A2(\core.registers[23][12] ),
    .B1(net1401),
    .B2(\core.registers[22][12] ),
    .X(_05015_));
 sky130_fd_sc_hd__or3_1 _10103_ (.A(net1687),
    .B(\core.registers[19][12] ),
    .C(net1448),
    .X(_05016_));
 sky130_fd_sc_hd__o221a_1 _10104_ (.A1(\core.registers[18][12] ),
    .A2(net1333),
    .B1(_05015_),
    .B2(net1436),
    .C1(_05016_),
    .X(_05017_));
 sky130_fd_sc_hd__mux4_1 _10105_ (.A0(\core.registers[16][12] ),
    .A1(\core.registers[17][12] ),
    .A2(\core.registers[20][12] ),
    .A3(\core.registers[21][12] ),
    .S0(net1401),
    .S1(net1448),
    .X(_05018_));
 sky130_fd_sc_hd__mux2_1 _10106_ (.A0(_05017_),
    .A1(_05018_),
    .S(net1469),
    .X(_05019_));
 sky130_fd_sc_hd__o21a_1 _10107_ (.A1(net1461),
    .A2(_05019_),
    .B1(net1488),
    .X(_05020_));
 sky130_fd_sc_hd__a22o_2 _10108_ (.A1(_05000_),
    .A2(_05008_),
    .B1(_05014_),
    .B2(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__a22o_2 _10109_ (.A1(net1069),
    .A2(net990),
    .B1(_05021_),
    .B2(net1065),
    .X(_05022_));
 sky130_fd_sc_hd__mux2_2 _10110_ (.A0(net453),
    .A1(_05022_),
    .S(net1282),
    .X(_05023_));
 sky130_fd_sc_hd__or2_4 _10111_ (.A(_04991_),
    .B(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__nand2_2 _10112_ (.A(_04991_),
    .B(_05023_),
    .Y(_05025_));
 sky130_fd_sc_hd__nand2_4 _10113_ (.A(_05024_),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__a221o_1 _10114_ (.A1(\core.pipe1_resultRegister[13] ),
    .A2(_04498_),
    .B1(net1268),
    .B2(\core.pipe1_csrData[13] ),
    .C1(net1187),
    .X(_05027_));
 sky130_fd_sc_hd__mux2_8 _10115_ (.A0(net111),
    .A1(net146),
    .S(net1805),
    .X(_05028_));
 sky130_fd_sc_hd__o32a_1 _10116_ (.A1(net1674),
    .A2(net1653),
    .A3(_05028_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[13] ),
    .X(_05029_));
 sky130_fd_sc_hd__mux2_1 _10117_ (.A0(\core.pipe1_loadResult[13] ),
    .A1(_05029_),
    .S(net1758),
    .X(_05030_));
 sky130_fd_sc_hd__or3b_2 _10118_ (.A(net1807),
    .B(_04935_),
    .C_N(_05030_),
    .X(_05031_));
 sky130_fd_sc_hd__nand2_1 _10119_ (.A(_04781_),
    .B(_04944_),
    .Y(_05032_));
 sky130_fd_sc_hd__a21o_1 _10120_ (.A1(_04945_),
    .A2(_05032_),
    .B1(_04551_),
    .X(_05033_));
 sky130_fd_sc_hd__mux2_8 _10121_ (.A0(net128),
    .A1(net164),
    .S(net1805),
    .X(_05034_));
 sky130_fd_sc_hd__o32a_1 _10122_ (.A1(net1674),
    .A2(net1661),
    .A3(_05034_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[29] ),
    .X(_05035_));
 sky130_fd_sc_hd__mux2_2 _10123_ (.A0(\core.pipe1_loadResult[29] ),
    .A1(_05035_),
    .S(net1757),
    .X(_05036_));
 sky130_fd_sc_hd__nand2_1 _10124_ (.A(net1233),
    .B(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__a21o_1 _10125_ (.A1(_04950_),
    .A2(_05037_),
    .B1(_04582_),
    .X(_05038_));
 sky130_fd_sc_hd__a32o_1 _10126_ (.A1(_04948_),
    .A2(_05033_),
    .A3(_05038_),
    .B1(_05031_),
    .B2(_04937_),
    .X(_05039_));
 sky130_fd_sc_hd__nand2_2 _10127_ (.A(net1189),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__a22o_4 _10128_ (.A1(\core.pipe1_resultRegister[13] ),
    .A2(net1271),
    .B1(_05027_),
    .B2(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__mux2_1 _10129_ (.A0(\core.registers[28][13] ),
    .A1(\core.registers[29][13] ),
    .S(net1539),
    .X(_05042_));
 sky130_fd_sc_hd__a221o_1 _10130_ (.A1(net1729),
    .A2(\core.registers[30][13] ),
    .B1(\core.registers[31][13] ),
    .B2(net1539),
    .C1(net1739),
    .X(_05043_));
 sky130_fd_sc_hd__mux2_1 _10131_ (.A0(\core.registers[12][13] ),
    .A1(\core.registers[13][13] ),
    .S(net1547),
    .X(_05044_));
 sky130_fd_sc_hd__mux2_1 _10132_ (.A0(\core.registers[14][13] ),
    .A1(\core.registers[15][13] ),
    .S(net1547),
    .X(_05045_));
 sky130_fd_sc_hd__mux2_1 _10133_ (.A0(\core.registers[8][13] ),
    .A1(\core.registers[9][13] ),
    .S(net1540),
    .X(_05046_));
 sky130_fd_sc_hd__mux2_1 _10134_ (.A0(\core.registers[10][13] ),
    .A1(\core.registers[11][13] ),
    .S(net1540),
    .X(_05047_));
 sky130_fd_sc_hd__mux2_1 _10135_ (.A0(_05046_),
    .A1(_05047_),
    .S(net1621),
    .X(_05048_));
 sky130_fd_sc_hd__mux2_1 _10136_ (.A0(\core.registers[24][13] ),
    .A1(\core.registers[25][13] ),
    .S(net1543),
    .X(_05049_));
 sky130_fd_sc_hd__and3_1 _10137_ (.A(net1844),
    .B(\core.registers[27][13] ),
    .C(net1543),
    .X(_05050_));
 sky130_fd_sc_hd__a211o_1 _10138_ (.A1(\core.registers[26][13] ),
    .A2(_04608_),
    .B1(_05050_),
    .C1(net1750),
    .X(_05051_));
 sky130_fd_sc_hd__a21o_1 _10139_ (.A1(net1739),
    .A2(_05049_),
    .B1(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__o21a_1 _10140_ (.A1(net1844),
    .A2(_05042_),
    .B1(_05043_),
    .X(_05053_));
 sky130_fd_sc_hd__mux2_1 _10141_ (.A0(_05044_),
    .A1(_05045_),
    .S(net1626),
    .X(_05054_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(_05053_),
    .A1(_05054_),
    .S(net1750),
    .X(_05055_));
 sky130_fd_sc_hd__o211a_1 _10143_ (.A1(net1829),
    .A2(_05048_),
    .B1(_05052_),
    .C1(net1746),
    .X(_05056_));
 sky130_fd_sc_hd__a211o_2 _10144_ (.A1(net1836),
    .A2(_05055_),
    .B1(_05056_),
    .C1(net1633),
    .X(_05057_));
 sky130_fd_sc_hd__or2_1 _10145_ (.A(\core.registers[22][13] ),
    .B(net1557),
    .X(_05058_));
 sky130_fd_sc_hd__or2_1 _10146_ (.A(\core.registers[6][13] ),
    .B(net1544),
    .X(_05059_));
 sky130_fd_sc_hd__o211a_1 _10147_ (.A1(net1730),
    .A2(\core.registers[7][13] ),
    .B1(net1623),
    .C1(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__mux2_1 _10148_ (.A0(\core.registers[4][13] ),
    .A1(\core.registers[5][13] ),
    .S(net1544),
    .X(_05061_));
 sky130_fd_sc_hd__a211o_1 _10149_ (.A1(net1606),
    .A2(_05061_),
    .B1(_05060_),
    .C1(net1580),
    .X(_05062_));
 sky130_fd_sc_hd__mux2_1 _10150_ (.A0(\core.registers[0][13] ),
    .A1(\core.registers[1][13] ),
    .S(net1544),
    .X(_05063_));
 sky130_fd_sc_hd__mux2_1 _10151_ (.A0(\core.registers[2][13] ),
    .A1(\core.registers[3][13] ),
    .S(net1545),
    .X(_05064_));
 sky130_fd_sc_hd__mux2_1 _10152_ (.A0(_05063_),
    .A1(_05064_),
    .S(net1623),
    .X(_05065_));
 sky130_fd_sc_hd__o211a_1 _10153_ (.A1(net1591),
    .A2(_05065_),
    .B1(_05062_),
    .C1(net1569),
    .X(_05066_));
 sky130_fd_sc_hd__mux2_1 _10154_ (.A0(\core.registers[16][13] ),
    .A1(\core.registers[17][13] ),
    .S(net1559),
    .X(_05067_));
 sky130_fd_sc_hd__mux2_1 _10155_ (.A0(\core.registers[18][13] ),
    .A1(\core.registers[19][13] ),
    .S(net1557),
    .X(_05068_));
 sky130_fd_sc_hd__mux2_1 _10156_ (.A0(_05067_),
    .A1(_05068_),
    .S(net1629),
    .X(_05069_));
 sky130_fd_sc_hd__o211a_1 _10157_ (.A1(net1733),
    .A2(\core.registers[23][13] ),
    .B1(net1629),
    .C1(_05058_),
    .X(_05070_));
 sky130_fd_sc_hd__mux2_1 _10158_ (.A0(\core.registers[20][13] ),
    .A1(\core.registers[21][13] ),
    .S(net1557),
    .X(_05071_));
 sky130_fd_sc_hd__a211o_1 _10159_ (.A1(net1609),
    .A2(_05071_),
    .B1(_05070_),
    .C1(net1583),
    .X(_05072_));
 sky130_fd_sc_hd__o211a_1 _10160_ (.A1(net1594),
    .A2(_05069_),
    .B1(_05072_),
    .C1(net1573),
    .X(_05073_));
 sky130_fd_sc_hd__o31a_1 _10161_ (.A1(net1637),
    .A2(_05066_),
    .A3(_05073_),
    .B1(_05057_),
    .X(_05074_));
 sky130_fd_sc_hd__o21a_1 _10162_ (.A1(net1159),
    .A2(_05074_),
    .B1(net1265),
    .X(_05075_));
 sky130_fd_sc_hd__o21ai_4 _10163_ (.A1(net1155),
    .A2(net985),
    .B1(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__o21ai_1 _10164_ (.A1(net1193),
    .A2(_05076_),
    .B1(net1162),
    .Y(_05077_));
 sky130_fd_sc_hd__o21a_2 _10165_ (.A1(net1880),
    .A2(net1279),
    .B1(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__mux2_1 _10166_ (.A0(\core.registers[28][13] ),
    .A1(\core.registers[29][13] ),
    .S(net1408),
    .X(_05079_));
 sky130_fd_sc_hd__a221o_1 _10167_ (.A1(net1692),
    .A2(\core.registers[30][13] ),
    .B1(\core.registers[31][13] ),
    .B2(net1408),
    .C1(net1710),
    .X(_05080_));
 sky130_fd_sc_hd__o21a_1 _10168_ (.A1(net1874),
    .A2(_05079_),
    .B1(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__mux2_1 _10169_ (.A0(\core.registers[14][13] ),
    .A1(\core.registers[15][13] ),
    .S(net1415),
    .X(_05082_));
 sky130_fd_sc_hd__mux2_1 _10170_ (.A0(\core.registers[12][13] ),
    .A1(\core.registers[13][13] ),
    .S(net1415),
    .X(_05083_));
 sky130_fd_sc_hd__mux2_1 _10171_ (.A0(_05082_),
    .A1(_05083_),
    .S(net1474),
    .X(_05084_));
 sky130_fd_sc_hd__mux2_1 _10172_ (.A0(_05081_),
    .A1(_05084_),
    .S(net1717),
    .X(_05085_));
 sky130_fd_sc_hd__a22o_1 _10173_ (.A1(net1692),
    .A2(\core.registers[26][13] ),
    .B1(\core.registers[27][13] ),
    .B2(net1412),
    .X(_05086_));
 sky130_fd_sc_hd__mux2_1 _10174_ (.A0(\core.registers[24][13] ),
    .A1(\core.registers[25][13] ),
    .S(net1412),
    .X(_05087_));
 sky130_fd_sc_hd__mux2_1 _10175_ (.A0(_05086_),
    .A1(_05087_),
    .S(net1710),
    .X(_05088_));
 sky130_fd_sc_hd__or2_1 _10176_ (.A(\core.registers[9][13] ),
    .B(net1377),
    .X(_05089_));
 sky130_fd_sc_hd__o21a_1 _10177_ (.A1(\core.registers[8][13] ),
    .A2(net1409),
    .B1(net1708),
    .X(_05090_));
 sky130_fd_sc_hd__a22o_1 _10178_ (.A1(net1692),
    .A2(\core.registers[10][13] ),
    .B1(\core.registers[11][13] ),
    .B2(net1409),
    .X(_05091_));
 sky130_fd_sc_hd__a221o_1 _10179_ (.A1(_05089_),
    .A2(_05090_),
    .B1(_05091_),
    .B2(net1873),
    .C1(net1856),
    .X(_05092_));
 sky130_fd_sc_hd__o21a_1 _10180_ (.A1(net1717),
    .A2(_05088_),
    .B1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__mux2_2 _10181_ (.A0(_05085_),
    .A1(_05093_),
    .S(net1715),
    .X(_05094_));
 sky130_fd_sc_hd__o22a_1 _10182_ (.A1(net1701),
    .A2(\core.registers[23][13] ),
    .B1(net1423),
    .B2(\core.registers[22][13] ),
    .X(_05095_));
 sky130_fd_sc_hd__or3_1 _10183_ (.A(net1701),
    .B(\core.registers[19][13] ),
    .C(net1459),
    .X(_05096_));
 sky130_fd_sc_hd__o221a_1 _10184_ (.A1(\core.registers[18][13] ),
    .A2(net1337),
    .B1(_05095_),
    .B2(net1440),
    .C1(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__mux4_1 _10185_ (.A0(\core.registers[16][13] ),
    .A1(\core.registers[17][13] ),
    .A2(\core.registers[20][13] ),
    .A3(\core.registers[21][13] ),
    .S0(net1423),
    .S1(net1459),
    .X(_05098_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(_05097_),
    .A1(_05098_),
    .S(net1475),
    .X(_05099_));
 sky130_fd_sc_hd__o22a_1 _10187_ (.A1(net1694),
    .A2(\core.registers[7][13] ),
    .B1(net1413),
    .B2(\core.registers[6][13] ),
    .X(_05100_));
 sky130_fd_sc_hd__or3_1 _10188_ (.A(net1694),
    .B(\core.registers[3][13] ),
    .C(net1454),
    .X(_05101_));
 sky130_fd_sc_hd__o221a_1 _10189_ (.A1(\core.registers[2][13] ),
    .A2(net1338),
    .B1(_05100_),
    .B2(net1439),
    .C1(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__mux4_1 _10190_ (.A0(\core.registers[0][13] ),
    .A1(\core.registers[1][13] ),
    .A2(\core.registers[4][13] ),
    .A3(\core.registers[5][13] ),
    .S0(net1413),
    .S1(net1454),
    .X(_05103_));
 sky130_fd_sc_hd__mux2_1 _10191_ (.A0(_05102_),
    .A1(_05103_),
    .S(net1473),
    .X(_05104_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(_05099_),
    .A1(_05104_),
    .S(net1462),
    .X(_05105_));
 sky130_fd_sc_hd__mux2_2 _10193_ (.A0(_05094_),
    .A1(_05105_),
    .S(net1487),
    .X(_05106_));
 sky130_fd_sc_hd__a22o_4 _10194_ (.A1(net1070),
    .A2(net985),
    .B1(_05106_),
    .B2(net1066),
    .X(_05107_));
 sky130_fd_sc_hd__mux2_4 _10195_ (.A0(net454),
    .A1(_05107_),
    .S(net1282),
    .X(_05108_));
 sky130_fd_sc_hd__or2_4 _10196_ (.A(_05078_),
    .B(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__nand2_4 _10197_ (.A(_05078_),
    .B(_05108_),
    .Y(_05110_));
 sky130_fd_sc_hd__nand2_8 _10198_ (.A(_05109_),
    .B(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__a221o_1 _10199_ (.A1(\core.pipe1_resultRegister[15] ),
    .A2(_04498_),
    .B1(net1268),
    .B2(\core.pipe1_csrData[15] ),
    .C1(net1187),
    .X(_05112_));
 sky130_fd_sc_hd__a21o_1 _10200_ (.A1(_04571_),
    .A2(_04935_),
    .B1(_04593_),
    .X(_05113_));
 sky130_fd_sc_hd__and2_1 _10201_ (.A(_04936_),
    .B(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__a21boi_1 _10202_ (.A1(_04589_),
    .A2(_04944_),
    .B1_N(_04945_),
    .Y(_05115_));
 sky130_fd_sc_hd__nand2_1 _10203_ (.A(_04566_),
    .B(net1233),
    .Y(_05116_));
 sky130_fd_sc_hd__a21o_1 _10204_ (.A1(_04950_),
    .A2(_05116_),
    .B1(_04582_),
    .X(_05117_));
 sky130_fd_sc_hd__o211a_1 _10205_ (.A1(_04551_),
    .A2(_05115_),
    .B1(_05117_),
    .C1(_04948_),
    .X(_05118_));
 sky130_fd_sc_hd__o21ai_2 _10206_ (.A1(_05114_),
    .A2(_05118_),
    .B1(net1189),
    .Y(_05119_));
 sky130_fd_sc_hd__a22o_1 _10207_ (.A1(\core.pipe1_resultRegister[15] ),
    .A2(net1271),
    .B1(_05112_),
    .B2(_05119_),
    .X(_05120_));
 sky130_fd_sc_hd__mux2_1 _10208_ (.A0(\core.registers[8][15] ),
    .A1(\core.registers[9][15] ),
    .S(net1539),
    .X(_05121_));
 sky130_fd_sc_hd__mux2_1 _10209_ (.A0(\core.registers[10][15] ),
    .A1(\core.registers[11][15] ),
    .S(net1539),
    .X(_05122_));
 sky130_fd_sc_hd__mux2_1 _10210_ (.A0(_05121_),
    .A1(_05122_),
    .S(net1621),
    .X(_05123_));
 sky130_fd_sc_hd__mux2_1 _10211_ (.A0(\core.registers[24][15] ),
    .A1(\core.registers[25][15] ),
    .S(net1539),
    .X(_05124_));
 sky130_fd_sc_hd__and3_1 _10212_ (.A(net1844),
    .B(\core.registers[27][15] ),
    .C(net1539),
    .X(_05125_));
 sky130_fd_sc_hd__a211o_1 _10213_ (.A1(\core.registers[26][15] ),
    .A2(_04608_),
    .B1(_05125_),
    .C1(net1750),
    .X(_05126_));
 sky130_fd_sc_hd__a21o_1 _10214_ (.A1(net1739),
    .A2(_05124_),
    .B1(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__mux2_1 _10215_ (.A0(\core.registers[12][15] ),
    .A1(\core.registers[13][15] ),
    .S(net1539),
    .X(_05128_));
 sky130_fd_sc_hd__mux2_1 _10216_ (.A0(\core.registers[14][15] ),
    .A1(\core.registers[15][15] ),
    .S(net1540),
    .X(_05129_));
 sky130_fd_sc_hd__mux2_1 _10217_ (.A0(\core.registers[28][15] ),
    .A1(\core.registers[29][15] ),
    .S(net1539),
    .X(_05130_));
 sky130_fd_sc_hd__a221o_1 _10218_ (.A1(net1729),
    .A2(\core.registers[30][15] ),
    .B1(\core.registers[31][15] ),
    .B2(net1539),
    .C1(net1739),
    .X(_05131_));
 sky130_fd_sc_hd__o21a_1 _10219_ (.A1(net1844),
    .A2(_05130_),
    .B1(_05131_),
    .X(_05132_));
 sky130_fd_sc_hd__mux2_1 _10220_ (.A0(_05128_),
    .A1(_05129_),
    .S(net1621),
    .X(_05133_));
 sky130_fd_sc_hd__mux2_1 _10221_ (.A0(_05132_),
    .A1(_05133_),
    .S(net1750),
    .X(_05134_));
 sky130_fd_sc_hd__o211a_1 _10222_ (.A1(net1827),
    .A2(_05123_),
    .B1(_05127_),
    .C1(net1747),
    .X(_05135_));
 sky130_fd_sc_hd__a211o_1 _10223_ (.A1(net1836),
    .A2(_05134_),
    .B1(_05135_),
    .C1(net1633),
    .X(_05136_));
 sky130_fd_sc_hd__or2_1 _10224_ (.A(\core.registers[22][15] ),
    .B(net1540),
    .X(_05137_));
 sky130_fd_sc_hd__or2_1 _10225_ (.A(\core.registers[6][15] ),
    .B(net1541),
    .X(_05138_));
 sky130_fd_sc_hd__o211a_1 _10226_ (.A1(net1728),
    .A2(\core.registers[7][15] ),
    .B1(net1621),
    .C1(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__mux2_1 _10227_ (.A0(\core.registers[4][15] ),
    .A1(\core.registers[5][15] ),
    .S(net1541),
    .X(_05140_));
 sky130_fd_sc_hd__a211o_1 _10228_ (.A1(net1605),
    .A2(_05140_),
    .B1(_05139_),
    .C1(net1584),
    .X(_05141_));
 sky130_fd_sc_hd__mux2_1 _10229_ (.A0(\core.registers[0][15] ),
    .A1(\core.registers[1][15] ),
    .S(net1541),
    .X(_05142_));
 sky130_fd_sc_hd__mux2_1 _10230_ (.A0(\core.registers[2][15] ),
    .A1(\core.registers[3][15] ),
    .S(net1542),
    .X(_05143_));
 sky130_fd_sc_hd__mux2_1 _10231_ (.A0(_05142_),
    .A1(_05143_),
    .S(net1621),
    .X(_05144_));
 sky130_fd_sc_hd__o211a_1 _10232_ (.A1(net1595),
    .A2(_05144_),
    .B1(_05141_),
    .C1(net1569),
    .X(_05145_));
 sky130_fd_sc_hd__mux2_1 _10233_ (.A0(\core.registers[16][15] ),
    .A1(\core.registers[17][15] ),
    .S(net1541),
    .X(_05146_));
 sky130_fd_sc_hd__mux2_1 _10234_ (.A0(\core.registers[18][15] ),
    .A1(\core.registers[19][15] ),
    .S(net1541),
    .X(_05147_));
 sky130_fd_sc_hd__mux2_1 _10235_ (.A0(_05146_),
    .A1(_05147_),
    .S(net1621),
    .X(_05148_));
 sky130_fd_sc_hd__o211a_1 _10236_ (.A1(net1729),
    .A2(\core.registers[23][15] ),
    .B1(net1621),
    .C1(_05137_),
    .X(_05149_));
 sky130_fd_sc_hd__mux2_1 _10237_ (.A0(\core.registers[20][15] ),
    .A1(\core.registers[21][15] ),
    .S(net1540),
    .X(_05150_));
 sky130_fd_sc_hd__a211o_1 _10238_ (.A1(net1606),
    .A2(_05150_),
    .B1(_05149_),
    .C1(net1580),
    .X(_05151_));
 sky130_fd_sc_hd__o211a_1 _10239_ (.A1(net1591),
    .A2(_05148_),
    .B1(_05151_),
    .C1(net1573),
    .X(_05152_));
 sky130_fd_sc_hd__o31a_1 _10240_ (.A1(net1637),
    .A2(_05145_),
    .A3(_05152_),
    .B1(_05136_),
    .X(_05153_));
 sky130_fd_sc_hd__o21a_1 _10241_ (.A1(net1159),
    .A2(_05153_),
    .B1(net1265),
    .X(_05154_));
 sky130_fd_sc_hd__o21ai_4 _10242_ (.A1(net1155),
    .A2(net982),
    .B1(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__o21a_1 _10243_ (.A1(net1193),
    .A2(_05155_),
    .B1(net1162),
    .X(_05156_));
 sky130_fd_sc_hd__a21oi_4 _10244_ (.A1(net1688),
    .A2(net1286),
    .B1(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__mux2_1 _10245_ (.A0(\core.registers[28][15] ),
    .A1(\core.registers[29][15] ),
    .S(net1408),
    .X(_05158_));
 sky130_fd_sc_hd__a221o_1 _10246_ (.A1(net1692),
    .A2(\core.registers[30][15] ),
    .B1(\core.registers[31][15] ),
    .B2(net1408),
    .C1(net1710),
    .X(_05159_));
 sky130_fd_sc_hd__o21a_1 _10247_ (.A1(net1874),
    .A2(_05158_),
    .B1(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__mux2_1 _10248_ (.A0(\core.registers[14][15] ),
    .A1(\core.registers[15][15] ),
    .S(net1409),
    .X(_05161_));
 sky130_fd_sc_hd__mux2_1 _10249_ (.A0(\core.registers[12][15] ),
    .A1(\core.registers[13][15] ),
    .S(net1408),
    .X(_05162_));
 sky130_fd_sc_hd__mux2_1 _10250_ (.A0(_05161_),
    .A1(_05162_),
    .S(net1472),
    .X(_05163_));
 sky130_fd_sc_hd__mux2_1 _10251_ (.A0(_05160_),
    .A1(_05163_),
    .S(net1717),
    .X(_05164_));
 sky130_fd_sc_hd__a22o_1 _10252_ (.A1(net1692),
    .A2(\core.registers[26][15] ),
    .B1(\core.registers[27][15] ),
    .B2(net1408),
    .X(_05165_));
 sky130_fd_sc_hd__mux2_1 _10253_ (.A0(\core.registers[24][15] ),
    .A1(\core.registers[25][15] ),
    .S(net1408),
    .X(_05166_));
 sky130_fd_sc_hd__mux2_1 _10254_ (.A0(_05165_),
    .A1(_05166_),
    .S(net1710),
    .X(_05167_));
 sky130_fd_sc_hd__or2_1 _10255_ (.A(\core.registers[9][15] ),
    .B(net1376),
    .X(_05168_));
 sky130_fd_sc_hd__o21a_1 _10256_ (.A1(\core.registers[8][15] ),
    .A2(net1408),
    .B1(net1710),
    .X(_05169_));
 sky130_fd_sc_hd__a22o_1 _10257_ (.A1(net1692),
    .A2(\core.registers[10][15] ),
    .B1(\core.registers[11][15] ),
    .B2(net1408),
    .X(_05170_));
 sky130_fd_sc_hd__a221o_1 _10258_ (.A1(_05168_),
    .A2(_05169_),
    .B1(_05170_),
    .B2(net1874),
    .C1(net1857),
    .X(_05171_));
 sky130_fd_sc_hd__o21a_1 _10259_ (.A1(net1717),
    .A2(_05167_),
    .B1(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__mux2_1 _10260_ (.A0(_05164_),
    .A1(_05172_),
    .S(net1715),
    .X(_05173_));
 sky130_fd_sc_hd__o22a_1 _10261_ (.A1(net1692),
    .A2(\core.registers[23][15] ),
    .B1(net1409),
    .B2(\core.registers[22][15] ),
    .X(_05174_));
 sky130_fd_sc_hd__or3_1 _10262_ (.A(net1692),
    .B(\core.registers[19][15] ),
    .C(net1453),
    .X(_05175_));
 sky130_fd_sc_hd__o221a_1 _10263_ (.A1(\core.registers[18][15] ),
    .A2(net1338),
    .B1(_05174_),
    .B2(net1439),
    .C1(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__mux4_1 _10264_ (.A0(\core.registers[16][15] ),
    .A1(\core.registers[17][15] ),
    .A2(\core.registers[20][15] ),
    .A3(\core.registers[21][15] ),
    .S0(net1410),
    .S1(net1453),
    .X(_05177_));
 sky130_fd_sc_hd__mux2_1 _10265_ (.A0(_05176_),
    .A1(_05177_),
    .S(net1472),
    .X(_05178_));
 sky130_fd_sc_hd__o22a_1 _10266_ (.A1(net1693),
    .A2(\core.registers[7][15] ),
    .B1(net1410),
    .B2(\core.registers[6][15] ),
    .X(_05179_));
 sky130_fd_sc_hd__or3_1 _10267_ (.A(net1693),
    .B(\core.registers[3][15] ),
    .C(net1453),
    .X(_05180_));
 sky130_fd_sc_hd__o221a_1 _10268_ (.A1(\core.registers[2][15] ),
    .A2(net1334),
    .B1(_05179_),
    .B2(net1439),
    .C1(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__mux4_1 _10269_ (.A0(\core.registers[0][15] ),
    .A1(\core.registers[1][15] ),
    .A2(\core.registers[4][15] ),
    .A3(\core.registers[5][15] ),
    .S0(net1410),
    .S1(net1453),
    .X(_05182_));
 sky130_fd_sc_hd__mux2_1 _10270_ (.A0(_05181_),
    .A1(_05182_),
    .S(net1472),
    .X(_05183_));
 sky130_fd_sc_hd__mux2_1 _10271_ (.A0(_05178_),
    .A1(_05183_),
    .S(net1462),
    .X(_05184_));
 sky130_fd_sc_hd__mux2_4 _10272_ (.A0(_05173_),
    .A1(_05184_),
    .S(net1487),
    .X(_05185_));
 sky130_fd_sc_hd__a22o_4 _10273_ (.A1(net1070),
    .A2(net982),
    .B1(_05185_),
    .B2(net1066),
    .X(_05186_));
 sky130_fd_sc_hd__mux2_4 _10274_ (.A0(net456),
    .A1(_05186_),
    .S(net1279),
    .X(_05187_));
 sky130_fd_sc_hd__nand2_4 _10275_ (.A(_05157_),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__inv_2 _10276_ (.A(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__or2_4 _10277_ (.A(_05157_),
    .B(_05187_),
    .X(_05190_));
 sky130_fd_sc_hd__nand2_8 _10278_ (.A(_05188_),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__clkinv_2 _10279_ (.A(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__a221o_1 _10280_ (.A1(\core.pipe1_resultRegister[14] ),
    .A2(_04498_),
    .B1(net1270),
    .B2(\core.pipe1_csrData[14] ),
    .C1(net1187),
    .X(_05193_));
 sky130_fd_sc_hd__mux2_8 _10281_ (.A0(net112),
    .A1(net147),
    .S(net1805),
    .X(_05194_));
 sky130_fd_sc_hd__o32a_1 _10282_ (.A1(net1675),
    .A2(net1653),
    .A3(_05194_),
    .B1(net1658),
    .B2(\coreWBInterface.readDataBuffered[14] ),
    .X(_05195_));
 sky130_fd_sc_hd__mux2_1 _10283_ (.A0(\core.pipe1_loadResult[14] ),
    .A1(_05195_),
    .S(net1758),
    .X(_05196_));
 sky130_fd_sc_hd__or3b_2 _10284_ (.A(net1808),
    .B(_04935_),
    .C_N(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__nand2_1 _10285_ (.A(_04701_),
    .B(_04944_),
    .Y(_05198_));
 sky130_fd_sc_hd__a21o_1 _10286_ (.A1(_04945_),
    .A2(_05198_),
    .B1(_04551_),
    .X(_05199_));
 sky130_fd_sc_hd__mux2_8 _10287_ (.A0(net130),
    .A1(net165),
    .S(net1805),
    .X(_05200_));
 sky130_fd_sc_hd__o32a_1 _10288_ (.A1(net1675),
    .A2(net1660),
    .A3(_05200_),
    .B1(net1658),
    .B2(\coreWBInterface.readDataBuffered[30] ),
    .X(_05201_));
 sky130_fd_sc_hd__mux2_2 _10289_ (.A0(\core.pipe1_loadResult[30] ),
    .A1(_05201_),
    .S(net1759),
    .X(_05202_));
 sky130_fd_sc_hd__nand2_1 _10290_ (.A(net1233),
    .B(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__a21o_1 _10291_ (.A1(_04950_),
    .A2(_05203_),
    .B1(_04582_),
    .X(_05204_));
 sky130_fd_sc_hd__a32o_2 _10292_ (.A1(_04948_),
    .A2(_05199_),
    .A3(_05204_),
    .B1(_05197_),
    .B2(_04937_),
    .X(_05205_));
 sky130_fd_sc_hd__nand2_1 _10293_ (.A(net1190),
    .B(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__a22o_2 _10294_ (.A1(\core.pipe1_resultRegister[14] ),
    .A2(net1271),
    .B1(_05193_),
    .B2(_05206_),
    .X(_05207_));
 sky130_fd_sc_hd__mux2_1 _10295_ (.A0(\core.registers[8][14] ),
    .A1(\core.registers[9][14] ),
    .S(net1535),
    .X(_05208_));
 sky130_fd_sc_hd__mux2_1 _10296_ (.A0(\core.registers[10][14] ),
    .A1(\core.registers[11][14] ),
    .S(net1535),
    .X(_05209_));
 sky130_fd_sc_hd__mux2_1 _10297_ (.A0(_05208_),
    .A1(_05209_),
    .S(net1620),
    .X(_05210_));
 sky130_fd_sc_hd__mux2_1 _10298_ (.A0(\core.registers[24][14] ),
    .A1(\core.registers[25][14] ),
    .S(net1538),
    .X(_05211_));
 sky130_fd_sc_hd__and3_1 _10299_ (.A(net1848),
    .B(\core.registers[27][14] ),
    .C(net1535),
    .X(_05212_));
 sky130_fd_sc_hd__a211o_1 _10300_ (.A1(\core.registers[26][14] ),
    .A2(_04608_),
    .B1(_05212_),
    .C1(net1752),
    .X(_05213_));
 sky130_fd_sc_hd__a21o_1 _10301_ (.A1(net1743),
    .A2(_05211_),
    .B1(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__mux2_1 _10302_ (.A0(\core.registers[12][14] ),
    .A1(\core.registers[13][14] ),
    .S(net1538),
    .X(_05215_));
 sky130_fd_sc_hd__mux2_1 _10303_ (.A0(\core.registers[14][14] ),
    .A1(\core.registers[15][14] ),
    .S(net1538),
    .X(_05216_));
 sky130_fd_sc_hd__mux2_1 _10304_ (.A0(\core.registers[28][14] ),
    .A1(\core.registers[29][14] ),
    .S(net1536),
    .X(_05217_));
 sky130_fd_sc_hd__a221o_1 _10305_ (.A1(net1727),
    .A2(\core.registers[30][14] ),
    .B1(\core.registers[31][14] ),
    .B2(net1536),
    .C1(net1743),
    .X(_05218_));
 sky130_fd_sc_hd__o21a_1 _10306_ (.A1(net1848),
    .A2(_05217_),
    .B1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__mux2_1 _10307_ (.A0(_05215_),
    .A1(_05216_),
    .S(net1620),
    .X(_05220_));
 sky130_fd_sc_hd__mux2_1 _10308_ (.A0(_05219_),
    .A1(_05220_),
    .S(net1752),
    .X(_05221_));
 sky130_fd_sc_hd__o211a_1 _10309_ (.A1(net1829),
    .A2(_05210_),
    .B1(_05214_),
    .C1(net1746),
    .X(_05222_));
 sky130_fd_sc_hd__a211o_1 _10310_ (.A1(net1836),
    .A2(_05221_),
    .B1(_05222_),
    .C1(net1633),
    .X(_05223_));
 sky130_fd_sc_hd__or2_1 _10311_ (.A(\core.registers[22][14] ),
    .B(net1536),
    .X(_05224_));
 sky130_fd_sc_hd__or2_1 _10312_ (.A(\core.registers[6][14] ),
    .B(net1537),
    .X(_05225_));
 sky130_fd_sc_hd__o211a_1 _10313_ (.A1(net1726),
    .A2(\core.registers[7][14] ),
    .B1(net1620),
    .C1(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__mux2_1 _10314_ (.A0(\core.registers[4][14] ),
    .A1(\core.registers[5][14] ),
    .S(net1537),
    .X(_05227_));
 sky130_fd_sc_hd__a211o_1 _10315_ (.A1(net1605),
    .A2(_05227_),
    .B1(_05226_),
    .C1(net1579),
    .X(_05228_));
 sky130_fd_sc_hd__mux2_1 _10316_ (.A0(\core.registers[0][14] ),
    .A1(\core.registers[1][14] ),
    .S(net1546),
    .X(_05229_));
 sky130_fd_sc_hd__mux2_1 _10317_ (.A0(\core.registers[2][14] ),
    .A1(\core.registers[3][14] ),
    .S(net1537),
    .X(_05230_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(_05229_),
    .A1(_05230_),
    .S(net1620),
    .X(_05231_));
 sky130_fd_sc_hd__o211a_1 _10319_ (.A1(net1590),
    .A2(_05231_),
    .B1(_05228_),
    .C1(net1569),
    .X(_05232_));
 sky130_fd_sc_hd__mux2_1 _10320_ (.A0(\core.registers[16][14] ),
    .A1(\core.registers[17][14] ),
    .S(net1537),
    .X(_05233_));
 sky130_fd_sc_hd__mux2_1 _10321_ (.A0(\core.registers[18][14] ),
    .A1(\core.registers[19][14] ),
    .S(net1537),
    .X(_05234_));
 sky130_fd_sc_hd__mux2_1 _10322_ (.A0(_05233_),
    .A1(_05234_),
    .S(net1622),
    .X(_05235_));
 sky130_fd_sc_hd__o211a_1 _10323_ (.A1(net1727),
    .A2(\core.registers[23][14] ),
    .B1(net1620),
    .C1(_05224_),
    .X(_05236_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(\core.registers[20][14] ),
    .A1(\core.registers[21][14] ),
    .S(net1537),
    .X(_05237_));
 sky130_fd_sc_hd__a211o_1 _10325_ (.A1(net1605),
    .A2(_05237_),
    .B1(_05236_),
    .C1(net1579),
    .X(_05238_));
 sky130_fd_sc_hd__o211a_1 _10326_ (.A1(net1590),
    .A2(_05235_),
    .B1(_05238_),
    .C1(net1573),
    .X(_05239_));
 sky130_fd_sc_hd__o31a_1 _10327_ (.A1(net1637),
    .A2(_05232_),
    .A3(_05239_),
    .B1(_05223_),
    .X(_05240_));
 sky130_fd_sc_hd__o21a_1 _10328_ (.A1(net1159),
    .A2(_05240_),
    .B1(net1266),
    .X(_05241_));
 sky130_fd_sc_hd__o21ai_4 _10329_ (.A1(net1156),
    .A2(net978),
    .B1(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__o21a_1 _10330_ (.A1(net1193),
    .A2(_05242_),
    .B1(net1162),
    .X(_05243_));
 sky130_fd_sc_hd__a21oi_4 _10331_ (.A1(_04423_),
    .A2(net1286),
    .B1(_05243_),
    .Y(_05244_));
 sky130_fd_sc_hd__or2_1 _10332_ (.A(\core.registers[24][14] ),
    .B(net1407),
    .X(_05245_));
 sky130_fd_sc_hd__o21a_1 _10333_ (.A1(\core.registers[25][14] ),
    .A2(net1377),
    .B1(net1708),
    .X(_05246_));
 sky130_fd_sc_hd__a22o_1 _10334_ (.A1(net1690),
    .A2(\core.registers[26][14] ),
    .B1(\core.registers[27][14] ),
    .B2(net1407),
    .X(_05247_));
 sky130_fd_sc_hd__a221o_1 _10335_ (.A1(_05245_),
    .A2(_05246_),
    .B1(_05247_),
    .B2(net1873),
    .C1(net1716),
    .X(_05248_));
 sky130_fd_sc_hd__a221o_1 _10336_ (.A1(net1690),
    .A2(\core.registers[10][14] ),
    .B1(\core.registers[11][14] ),
    .B2(net1404),
    .C1(net1708),
    .X(_05249_));
 sky130_fd_sc_hd__a21o_1 _10337_ (.A1(\core.registers[8][14] ),
    .A2(net1377),
    .B1(net1873),
    .X(_05250_));
 sky130_fd_sc_hd__a21o_1 _10338_ (.A1(\core.registers[9][14] ),
    .A2(net1404),
    .B1(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__a21o_1 _10339_ (.A1(_05249_),
    .A2(_05251_),
    .B1(net1856),
    .X(_05252_));
 sky130_fd_sc_hd__a21o_1 _10340_ (.A1(_05248_),
    .A2(_05252_),
    .B1(net1866),
    .X(_05253_));
 sky130_fd_sc_hd__a221o_1 _10341_ (.A1(net1690),
    .A2(\core.registers[30][14] ),
    .B1(\core.registers[31][14] ),
    .B2(net1405),
    .C1(net1707),
    .X(_05254_));
 sky130_fd_sc_hd__mux2_1 _10342_ (.A0(\core.registers[28][14] ),
    .A1(\core.registers[29][14] ),
    .S(net1405),
    .X(_05255_));
 sky130_fd_sc_hd__o21a_1 _10343_ (.A1(net1872),
    .A2(_05255_),
    .B1(_05254_),
    .X(_05256_));
 sky130_fd_sc_hd__mux2_1 _10344_ (.A0(\core.registers[12][14] ),
    .A1(\core.registers[13][14] ),
    .S(net1404),
    .X(_05257_));
 sky130_fd_sc_hd__mux2_1 _10345_ (.A0(\core.registers[14][14] ),
    .A1(\core.registers[15][14] ),
    .S(net1407),
    .X(_05258_));
 sky130_fd_sc_hd__mux2_1 _10346_ (.A0(_05257_),
    .A1(_05258_),
    .S(net1483),
    .X(_05259_));
 sky130_fd_sc_hd__mux2_1 _10347_ (.A0(_05256_),
    .A1(_05259_),
    .S(net1716),
    .X(_05260_));
 sky130_fd_sc_hd__o21a_1 _10348_ (.A1(net1715),
    .A2(_05260_),
    .B1(net1492),
    .X(_05261_));
 sky130_fd_sc_hd__o22a_1 _10349_ (.A1(net1689),
    .A2(\core.registers[7][14] ),
    .B1(net1406),
    .B2(\core.registers[6][14] ),
    .X(_05262_));
 sky130_fd_sc_hd__or3_1 _10350_ (.A(net1689),
    .B(\core.registers[3][14] ),
    .C(net1452),
    .X(_05263_));
 sky130_fd_sc_hd__o221a_1 _10351_ (.A1(\core.registers[2][14] ),
    .A2(net1333),
    .B1(_05262_),
    .B2(net1438),
    .C1(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__mux4_1 _10352_ (.A0(\core.registers[0][14] ),
    .A1(\core.registers[1][14] ),
    .A2(\core.registers[4][14] ),
    .A3(\core.registers[5][14] ),
    .S0(net1414),
    .S1(net1452),
    .X(_05265_));
 sky130_fd_sc_hd__mux2_1 _10353_ (.A0(_05264_),
    .A1(_05265_),
    .S(net1472),
    .X(_05266_));
 sky130_fd_sc_hd__or2_1 _10354_ (.A(net1464),
    .B(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__o22a_1 _10355_ (.A1(net1690),
    .A2(\core.registers[23][14] ),
    .B1(net1405),
    .B2(\core.registers[22][14] ),
    .X(_05268_));
 sky130_fd_sc_hd__or3_1 _10356_ (.A(net1690),
    .B(\core.registers[19][14] ),
    .C(net1451),
    .X(_05269_));
 sky130_fd_sc_hd__o221a_1 _10357_ (.A1(\core.registers[18][14] ),
    .A2(net1334),
    .B1(_05268_),
    .B2(net1438),
    .C1(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__mux4_1 _10358_ (.A0(\core.registers[16][14] ),
    .A1(\core.registers[17][14] ),
    .A2(\core.registers[20][14] ),
    .A3(\core.registers[21][14] ),
    .S0(net1406),
    .S1(net1451),
    .X(_05271_));
 sky130_fd_sc_hd__mux2_1 _10359_ (.A0(_05270_),
    .A1(_05271_),
    .S(net1472),
    .X(_05272_));
 sky130_fd_sc_hd__o21a_1 _10360_ (.A1(net1462),
    .A2(_05272_),
    .B1(net1488),
    .X(_05273_));
 sky130_fd_sc_hd__a22o_2 _10361_ (.A1(_05253_),
    .A2(_05261_),
    .B1(_05267_),
    .B2(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__a22o_4 _10362_ (.A1(net1071),
    .A2(net978),
    .B1(_05274_),
    .B2(net1066),
    .X(_05275_));
 sky130_fd_sc_hd__mux2_4 _10363_ (.A0(net455),
    .A1(_05275_),
    .S(net1279),
    .X(_05276_));
 sky130_fd_sc_hd__or2_4 _10364_ (.A(_05244_),
    .B(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__nand2_4 _10365_ (.A(_05244_),
    .B(_05276_),
    .Y(_05278_));
 sky130_fd_sc_hd__nand2_8 _10366_ (.A(_05277_),
    .B(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__inv_2 _10367_ (.A(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__and4_2 _10368_ (.A(_05026_),
    .B(_05111_),
    .C(_05191_),
    .D(_05279_),
    .X(_05281_));
 sky130_fd_sc_hd__a221o_1 _10369_ (.A1(\core.pipe1_resultRegister[11] ),
    .A2(_04498_),
    .B1(net1270),
    .B2(\core.pipe1_csrData[11] ),
    .C1(net1187),
    .X(_05282_));
 sky130_fd_sc_hd__mux2_8 _10370_ (.A0(net109),
    .A1(net144),
    .S(net1805),
    .X(_05283_));
 sky130_fd_sc_hd__o32a_1 _10371_ (.A1(net1674),
    .A2(net1653),
    .A3(_05283_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[11] ),
    .X(_05284_));
 sky130_fd_sc_hd__mux2_1 _10372_ (.A0(\core.pipe1_loadResult[11] ),
    .A1(_05284_),
    .S(net1758),
    .X(_05285_));
 sky130_fd_sc_hd__or3b_1 _10373_ (.A(net1807),
    .B(_04935_),
    .C_N(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__mux2_8 _10374_ (.A0(net117),
    .A1(net153),
    .S(net1805),
    .X(_05287_));
 sky130_fd_sc_hd__o32a_1 _10375_ (.A1(net1673),
    .A2(net1651),
    .A3(_05287_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[19] ),
    .X(_05288_));
 sky130_fd_sc_hd__mux2_2 _10376_ (.A0(\core.pipe1_loadResult[19] ),
    .A1(_05288_),
    .S(net1758),
    .X(_05289_));
 sky130_fd_sc_hd__nand2_1 _10377_ (.A(_04944_),
    .B(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__a21o_1 _10378_ (.A1(_04945_),
    .A2(_05290_),
    .B1(_04551_),
    .X(_05291_));
 sky130_fd_sc_hd__mux2_8 _10379_ (.A0(net126),
    .A1(net161),
    .S(net1805),
    .X(_05292_));
 sky130_fd_sc_hd__o32a_1 _10380_ (.A1(net1673),
    .A2(net1660),
    .A3(_05292_),
    .B1(net1658),
    .B2(\coreWBInterface.readDataBuffered[27] ),
    .X(_05293_));
 sky130_fd_sc_hd__mux2_2 _10381_ (.A0(\core.pipe1_loadResult[27] ),
    .A1(_05293_),
    .S(net1757),
    .X(_05294_));
 sky130_fd_sc_hd__nand2_1 _10382_ (.A(_04949_),
    .B(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__a21o_1 _10383_ (.A1(_04950_),
    .A2(_05295_),
    .B1(_04582_),
    .X(_05296_));
 sky130_fd_sc_hd__a32o_2 _10384_ (.A1(_04948_),
    .A2(_05291_),
    .A3(_05296_),
    .B1(_05286_),
    .B2(_04937_),
    .X(_05297_));
 sky130_fd_sc_hd__nand2_1 _10385_ (.A(net1190),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__a22o_2 _10386_ (.A1(\core.pipe1_resultRegister[11] ),
    .A2(net1271),
    .B1(_05282_),
    .B2(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__or2_1 _10387_ (.A(\core.registers[24][11] ),
    .B(net1400),
    .X(_05300_));
 sky130_fd_sc_hd__o21a_1 _10388_ (.A1(\core.registers[25][11] ),
    .A2(net1377),
    .B1(net1707),
    .X(_05301_));
 sky130_fd_sc_hd__a22o_1 _10389_ (.A1(net1686),
    .A2(\core.registers[26][11] ),
    .B1(\core.registers[27][11] ),
    .B2(net1400),
    .X(_05302_));
 sky130_fd_sc_hd__a221o_1 _10390_ (.A1(_05300_),
    .A2(_05301_),
    .B1(_05302_),
    .B2(net1872),
    .C1(net1716),
    .X(_05303_));
 sky130_fd_sc_hd__a221o_1 _10391_ (.A1(net1686),
    .A2(\core.registers[10][11] ),
    .B1(\core.registers[11][11] ),
    .B2(net1399),
    .C1(net1706),
    .X(_05304_));
 sky130_fd_sc_hd__a21o_1 _10392_ (.A1(\core.registers[8][11] ),
    .A2(net1374),
    .B1(net1870),
    .X(_05305_));
 sky130_fd_sc_hd__a21o_1 _10393_ (.A1(\core.registers[9][11] ),
    .A2(net1400),
    .B1(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__a21o_1 _10394_ (.A1(_05304_),
    .A2(_05306_),
    .B1(net1861),
    .X(_05307_));
 sky130_fd_sc_hd__a21o_1 _10395_ (.A1(_05303_),
    .A2(_05307_),
    .B1(net1863),
    .X(_05308_));
 sky130_fd_sc_hd__a221o_1 _10396_ (.A1(net1686),
    .A2(\core.registers[30][11] ),
    .B1(\core.registers[31][11] ),
    .B2(net1399),
    .C1(net1706),
    .X(_05309_));
 sky130_fd_sc_hd__mux2_1 _10397_ (.A0(\core.registers[28][11] ),
    .A1(\core.registers[29][11] ),
    .S(net1399),
    .X(_05310_));
 sky130_fd_sc_hd__o21a_1 _10398_ (.A1(net1871),
    .A2(_05310_),
    .B1(_05309_),
    .X(_05311_));
 sky130_fd_sc_hd__mux2_1 _10399_ (.A0(\core.registers[12][11] ),
    .A1(\core.registers[13][11] ),
    .S(net1400),
    .X(_05312_));
 sky130_fd_sc_hd__mux2_1 _10400_ (.A0(\core.registers[14][11] ),
    .A1(\core.registers[15][11] ),
    .S(net1400),
    .X(_05313_));
 sky130_fd_sc_hd__mux2_1 _10401_ (.A0(_05312_),
    .A1(_05313_),
    .S(net1483),
    .X(_05314_));
 sky130_fd_sc_hd__mux2_1 _10402_ (.A0(_05311_),
    .A1(_05314_),
    .S(net1716),
    .X(_05315_));
 sky130_fd_sc_hd__o21a_1 _10403_ (.A1(net1715),
    .A2(_05315_),
    .B1(net1490),
    .X(_05316_));
 sky130_fd_sc_hd__o22a_1 _10404_ (.A1(net1687),
    .A2(\core.registers[7][11] ),
    .B1(net1403),
    .B2(\core.registers[6][11] ),
    .X(_05317_));
 sky130_fd_sc_hd__or3_1 _10405_ (.A(net1687),
    .B(\core.registers[3][11] ),
    .C(net1449),
    .X(_05318_));
 sky130_fd_sc_hd__o221a_1 _10406_ (.A1(\core.registers[2][11] ),
    .A2(net1332),
    .B1(_05317_),
    .B2(net1436),
    .C1(_05318_),
    .X(_05319_));
 sky130_fd_sc_hd__mux4_1 _10407_ (.A0(\core.registers[0][11] ),
    .A1(\core.registers[1][11] ),
    .A2(\core.registers[4][11] ),
    .A3(\core.registers[5][11] ),
    .S0(net1403),
    .S1(net1449),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_1 _10408_ (.A0(_05319_),
    .A1(_05320_),
    .S(net1469),
    .X(_05321_));
 sky130_fd_sc_hd__or2_1 _10409_ (.A(net1464),
    .B(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__o22a_1 _10410_ (.A1(net1689),
    .A2(\core.registers[23][11] ),
    .B1(net1406),
    .B2(\core.registers[22][11] ),
    .X(_05323_));
 sky130_fd_sc_hd__or3_1 _10411_ (.A(net1689),
    .B(\core.registers[19][11] ),
    .C(net1451),
    .X(_05324_));
 sky130_fd_sc_hd__o221a_1 _10412_ (.A1(\core.registers[18][11] ),
    .A2(net1332),
    .B1(_05323_),
    .B2(net1436),
    .C1(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__mux4_1 _10413_ (.A0(\core.registers[16][11] ),
    .A1(\core.registers[17][11] ),
    .A2(\core.registers[20][11] ),
    .A3(\core.registers[21][11] ),
    .S0(net1401),
    .S1(net1448),
    .X(_05326_));
 sky130_fd_sc_hd__mux2_1 _10414_ (.A0(_05325_),
    .A1(_05326_),
    .S(net1470),
    .X(_05327_));
 sky130_fd_sc_hd__o21a_1 _10415_ (.A1(net1461),
    .A2(_05327_),
    .B1(net1486),
    .X(_05328_));
 sky130_fd_sc_hd__a22o_2 _10416_ (.A1(_05308_),
    .A2(_05316_),
    .B1(_05322_),
    .B2(_05328_),
    .X(_05329_));
 sky130_fd_sc_hd__a22o_4 _10417_ (.A1(net1069),
    .A2(net973),
    .B1(_05329_),
    .B2(net1065),
    .X(_05330_));
 sky130_fd_sc_hd__mux2_8 _10418_ (.A0(net452),
    .A1(_05330_),
    .S(net1282),
    .X(_05331_));
 sky130_fd_sc_hd__mux2_1 _10419_ (.A0(\core.registers[14][11] ),
    .A1(\core.registers[15][11] ),
    .S(net1529),
    .X(_05332_));
 sky130_fd_sc_hd__mux2_1 _10420_ (.A0(\core.registers[12][11] ),
    .A1(\core.registers[13][11] ),
    .S(net1529),
    .X(_05333_));
 sky130_fd_sc_hd__mux2_1 _10421_ (.A0(_05332_),
    .A1(_05333_),
    .S(net1602),
    .X(_05334_));
 sky130_fd_sc_hd__mux2_1 _10422_ (.A0(\core.registers[28][11] ),
    .A1(\core.registers[29][11] ),
    .S(net1528),
    .X(_05335_));
 sky130_fd_sc_hd__a221o_1 _10423_ (.A1(net1723),
    .A2(\core.registers[30][11] ),
    .B1(\core.registers[31][11] ),
    .B2(net1528),
    .C1(net1737),
    .X(_05336_));
 sky130_fd_sc_hd__o21a_1 _10424_ (.A1(net1841),
    .A2(_05335_),
    .B1(_05336_),
    .X(_05337_));
 sky130_fd_sc_hd__mux2_1 _10425_ (.A0(\core.registers[8][11] ),
    .A1(\core.registers[9][11] ),
    .S(net1531),
    .X(_05338_));
 sky130_fd_sc_hd__mux2_1 _10426_ (.A0(\core.registers[10][11] ),
    .A1(\core.registers[11][11] ),
    .S(net1528),
    .X(_05339_));
 sky130_fd_sc_hd__mux2_1 _10427_ (.A0(_05338_),
    .A1(_05339_),
    .S(net1619),
    .X(_05340_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(\core.registers[24][11] ),
    .A1(\core.registers[25][11] ),
    .S(net1529),
    .X(_05341_));
 sky130_fd_sc_hd__a22o_1 _10429_ (.A1(net1723),
    .A2(\core.registers[26][11] ),
    .B1(\core.registers[27][11] ),
    .B2(net1529),
    .X(_05342_));
 sky130_fd_sc_hd__mux2_1 _10430_ (.A0(_05341_),
    .A1(_05342_),
    .S(net1841),
    .X(_05343_));
 sky130_fd_sc_hd__mux4_2 _10431_ (.A0(_05334_),
    .A1(_05337_),
    .A2(_05340_),
    .A3(_05343_),
    .S0(net1825),
    .S1(net1745),
    .X(_05344_));
 sky130_fd_sc_hd__and3_1 _10432_ (.A(net1852),
    .B(\core.registers[5][11] ),
    .C(net1662),
    .X(_05345_));
 sky130_fd_sc_hd__a21o_1 _10433_ (.A1(\core.registers[4][11] ),
    .A2(net1497),
    .B1(net1578),
    .X(_05346_));
 sky130_fd_sc_hd__o31a_1 _10434_ (.A1(\core.registers[1][11] ),
    .A2(net1588),
    .A3(net1497),
    .B1(net1604),
    .X(_05347_));
 sky130_fd_sc_hd__o221a_1 _10435_ (.A1(\core.registers[0][11] ),
    .A2(net1341),
    .B1(_05345_),
    .B2(_05346_),
    .C1(_05347_),
    .X(_05348_));
 sky130_fd_sc_hd__o22a_1 _10436_ (.A1(net1724),
    .A2(\core.registers[7][11] ),
    .B1(net1533),
    .B2(\core.registers[6][11] ),
    .X(_05349_));
 sky130_fd_sc_hd__o31a_1 _10437_ (.A1(net1724),
    .A2(\core.registers[3][11] ),
    .A3(net1589),
    .B1(net1619),
    .X(_05350_));
 sky130_fd_sc_hd__o221a_1 _10438_ (.A1(\core.registers[2][11] ),
    .A2(net1341),
    .B1(_05349_),
    .B2(net1578),
    .C1(_05350_),
    .X(_05351_));
 sky130_fd_sc_hd__and3_1 _10439_ (.A(net1852),
    .B(\core.registers[21][11] ),
    .C(net1662),
    .X(_05352_));
 sky130_fd_sc_hd__a21o_1 _10440_ (.A1(\core.registers[20][11] ),
    .A2(net1496),
    .B1(net1577),
    .X(_05353_));
 sky130_fd_sc_hd__o31a_1 _10441_ (.A1(\core.registers[17][11] ),
    .A2(net1589),
    .A3(net1496),
    .B1(net1602),
    .X(_05354_));
 sky130_fd_sc_hd__o221a_1 _10442_ (.A1(\core.registers[16][11] ),
    .A2(net1341),
    .B1(_05352_),
    .B2(_05353_),
    .C1(_05354_),
    .X(_05355_));
 sky130_fd_sc_hd__o22a_1 _10443_ (.A1(net1726),
    .A2(\core.registers[23][11] ),
    .B1(net1537),
    .B2(\core.registers[22][11] ),
    .X(_05356_));
 sky130_fd_sc_hd__o31a_1 _10444_ (.A1(net1726),
    .A2(\core.registers[19][11] ),
    .A3(net1590),
    .B1(net1620),
    .X(_05357_));
 sky130_fd_sc_hd__o221a_1 _10445_ (.A1(\core.registers[18][11] ),
    .A2(net1341),
    .B1(_05356_),
    .B2(net1579),
    .C1(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__o31a_1 _10446_ (.A1(net1568),
    .A2(_05355_),
    .A3(_05358_),
    .B1(net1632),
    .X(_05359_));
 sky130_fd_sc_hd__o31a_1 _10447_ (.A1(net1572),
    .A2(_05348_),
    .A3(_05351_),
    .B1(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__a211o_1 _10448_ (.A1(net1636),
    .A2(_05344_),
    .B1(_05360_),
    .C1(net1158),
    .X(_05361_));
 sky130_fd_sc_hd__o211a_2 _10449_ (.A1(net1154),
    .A2(net973),
    .B1(_05361_),
    .C1(net1264),
    .X(_05362_));
 sky130_fd_sc_hd__or2_1 _10450_ (.A(net1815),
    .B(_04484_),
    .X(_05363_));
 sky130_fd_sc_hd__o211a_4 _10451_ (.A1(net1194),
    .A2(_05362_),
    .B1(_05363_),
    .C1(net1282),
    .X(_05364_));
 sky130_fd_sc_hd__nor2_1 _10452_ (.A(_05331_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__inv_2 _10453_ (.A(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__nand2_1 _10454_ (.A(_05331_),
    .B(_05364_),
    .Y(_05367_));
 sky130_fd_sc_hd__xor2_4 _10455_ (.A(_05331_),
    .B(_05364_),
    .X(_05368_));
 sky130_fd_sc_hd__nand2_1 _10456_ (.A(_05366_),
    .B(_05367_),
    .Y(_05369_));
 sky130_fd_sc_hd__a221oi_4 _10457_ (.A1(\core.pipe1_resultRegister[10] ),
    .A2(_04498_),
    .B1(net1270),
    .B2(\core.pipe1_csrData[10] ),
    .C1(net1187),
    .Y(_05370_));
 sky130_fd_sc_hd__mux2_8 _10458_ (.A0(net108),
    .A1(net143),
    .S(net1805),
    .X(_05371_));
 sky130_fd_sc_hd__o32a_1 _10459_ (.A1(net1674),
    .A2(net1654),
    .A3(_05371_),
    .B1(net1659),
    .B2(\coreWBInterface.readDataBuffered[10] ),
    .X(_05372_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(\core.pipe1_loadResult[10] ),
    .A1(_05372_),
    .S(net1759),
    .X(_05373_));
 sky130_fd_sc_hd__or3b_1 _10461_ (.A(net1806),
    .B(_04935_),
    .C_N(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__mux2_8 _10462_ (.A0(net116),
    .A1(net152),
    .S(net1805),
    .X(_05375_));
 sky130_fd_sc_hd__o32a_1 _10463_ (.A1(net1676),
    .A2(_04583_),
    .A3(_05375_),
    .B1(net1659),
    .B2(\coreWBInterface.readDataBuffered[18] ),
    .X(_05376_));
 sky130_fd_sc_hd__mux2_1 _10464_ (.A0(\core.pipe1_loadResult[18] ),
    .A1(_05376_),
    .S(net1759),
    .X(_05377_));
 sky130_fd_sc_hd__nand2_1 _10465_ (.A(_04944_),
    .B(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__a21o_1 _10466_ (.A1(_04945_),
    .A2(_05378_),
    .B1(_04551_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_8 _10467_ (.A0(net125),
    .A1(net160),
    .S(net1805),
    .X(_05380_));
 sky130_fd_sc_hd__o32a_1 _10468_ (.A1(net1673),
    .A2(net1660),
    .A3(_05380_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[26] ),
    .X(_05381_));
 sky130_fd_sc_hd__mux2_4 _10469_ (.A0(\core.pipe1_loadResult[26] ),
    .A1(_05381_),
    .S(net1757),
    .X(_05382_));
 sky130_fd_sc_hd__nand2_1 _10470_ (.A(net1233),
    .B(_05382_),
    .Y(_05383_));
 sky130_fd_sc_hd__a21o_1 _10471_ (.A1(_04950_),
    .A2(_05383_),
    .B1(_04582_),
    .X(_05384_));
 sky130_fd_sc_hd__a32o_2 _10472_ (.A1(_04948_),
    .A2(_05379_),
    .A3(_05384_),
    .B1(_05374_),
    .B2(_04937_),
    .X(_05385_));
 sky130_fd_sc_hd__a21oi_2 _10473_ (.A1(net1191),
    .A2(_05385_),
    .B1(_05370_),
    .Y(_05386_));
 sky130_fd_sc_hd__a21o_4 _10474_ (.A1(\core.pipe1_resultRegister[10] ),
    .A2(net1271),
    .B1(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__a211o_4 _10475_ (.A1(\core.pipe1_resultRegister[10] ),
    .A2(net1271),
    .B1(net1155),
    .C1(_05386_),
    .X(_05388_));
 sky130_fd_sc_hd__mux2_1 _10476_ (.A0(\core.registers[14][10] ),
    .A1(\core.registers[15][10] ),
    .S(net1535),
    .X(_05389_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(\core.registers[12][10] ),
    .A1(\core.registers[13][10] ),
    .S(net1535),
    .X(_05390_));
 sky130_fd_sc_hd__mux2_1 _10478_ (.A0(_05389_),
    .A1(_05390_),
    .S(net1605),
    .X(_05391_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(\core.registers[28][10] ),
    .A1(\core.registers[29][10] ),
    .S(net1536),
    .X(_05392_));
 sky130_fd_sc_hd__a221o_1 _10480_ (.A1(net1727),
    .A2(\core.registers[30][10] ),
    .B1(\core.registers[31][10] ),
    .B2(net1536),
    .C1(net1743),
    .X(_05393_));
 sky130_fd_sc_hd__o21a_1 _10481_ (.A1(net1848),
    .A2(_05392_),
    .B1(_05393_),
    .X(_05394_));
 sky130_fd_sc_hd__mux2_1 _10482_ (.A0(\core.registers[8][10] ),
    .A1(\core.registers[9][10] ),
    .S(net1535),
    .X(_05395_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(\core.registers[10][10] ),
    .A1(\core.registers[11][10] ),
    .S(net1535),
    .X(_05396_));
 sky130_fd_sc_hd__mux2_1 _10484_ (.A0(_05395_),
    .A1(_05396_),
    .S(net1620),
    .X(_05397_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(\core.registers[24][10] ),
    .A1(\core.registers[25][10] ),
    .S(net1536),
    .X(_05398_));
 sky130_fd_sc_hd__a22o_1 _10486_ (.A1(net1727),
    .A2(\core.registers[26][10] ),
    .B1(\core.registers[27][10] ),
    .B2(net1536),
    .X(_05399_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(_05398_),
    .A1(_05399_),
    .S(net1848),
    .X(_05400_));
 sky130_fd_sc_hd__mux4_2 _10488_ (.A0(_05391_),
    .A1(_05394_),
    .A2(_05397_),
    .A3(_05400_),
    .S0(net1829),
    .S1(net1746),
    .X(_05401_));
 sky130_fd_sc_hd__and3_1 _10489_ (.A(net1852),
    .B(\core.registers[5][10] ),
    .C(net1662),
    .X(_05402_));
 sky130_fd_sc_hd__a21o_1 _10490_ (.A1(\core.registers[4][10] ),
    .A2(net1500),
    .B1(net1579),
    .X(_05403_));
 sky130_fd_sc_hd__o31a_1 _10491_ (.A1(\core.registers[1][10] ),
    .A2(net1590),
    .A3(net1500),
    .B1(net1606),
    .X(_05404_));
 sky130_fd_sc_hd__o221a_1 _10492_ (.A1(\core.registers[0][10] ),
    .A2(net1341),
    .B1(_05402_),
    .B2(_05403_),
    .C1(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__o22a_1 _10493_ (.A1(net1726),
    .A2(\core.registers[7][10] ),
    .B1(net1546),
    .B2(\core.registers[6][10] ),
    .X(_05406_));
 sky130_fd_sc_hd__o31a_1 _10494_ (.A1(net1726),
    .A2(\core.registers[3][10] ),
    .A3(net1591),
    .B1(net1623),
    .X(_05407_));
 sky130_fd_sc_hd__o221a_1 _10495_ (.A1(\core.registers[2][10] ),
    .A2(net1339),
    .B1(_05406_),
    .B2(net1579),
    .C1(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__and3_1 _10496_ (.A(net1852),
    .B(\core.registers[21][10] ),
    .C(net1662),
    .X(_05409_));
 sky130_fd_sc_hd__a21o_1 _10497_ (.A1(\core.registers[20][10] ),
    .A2(net1498),
    .B1(net1579),
    .X(_05410_));
 sky130_fd_sc_hd__o31a_1 _10498_ (.A1(\core.registers[17][10] ),
    .A2(net1590),
    .A3(net1500),
    .B1(net1605),
    .X(_05411_));
 sky130_fd_sc_hd__o221a_1 _10499_ (.A1(\core.registers[16][10] ),
    .A2(net1339),
    .B1(_05409_),
    .B2(_05410_),
    .C1(_05411_),
    .X(_05412_));
 sky130_fd_sc_hd__o22a_1 _10500_ (.A1(net1726),
    .A2(\core.registers[23][10] ),
    .B1(net1537),
    .B2(\core.registers[22][10] ),
    .X(_05413_));
 sky130_fd_sc_hd__o31a_1 _10501_ (.A1(net1726),
    .A2(\core.registers[19][10] ),
    .A3(net1590),
    .B1(net1622),
    .X(_05414_));
 sky130_fd_sc_hd__o221a_1 _10502_ (.A1(\core.registers[18][10] ),
    .A2(net1341),
    .B1(_05413_),
    .B2(net1579),
    .C1(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__o31a_1 _10503_ (.A1(net1569),
    .A2(_05412_),
    .A3(_05415_),
    .B1(net1633),
    .X(_05416_));
 sky130_fd_sc_hd__o31a_1 _10504_ (.A1(net1573),
    .A2(_05405_),
    .A3(_05408_),
    .B1(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__a211o_4 _10505_ (.A1(net1637),
    .A2(_05401_),
    .B1(_05417_),
    .C1(net1159),
    .X(_05418_));
 sky130_fd_sc_hd__a31o_4 _10506_ (.A1(net1266),
    .A2(_05388_),
    .A3(_05418_),
    .B1(net1194),
    .X(_05419_));
 sky130_fd_sc_hd__o21a_2 _10507_ (.A1(net1817),
    .A2(_04484_),
    .B1(net1282),
    .X(_05420_));
 sky130_fd_sc_hd__nand2_4 _10508_ (.A(_05419_),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__nor2_2 _10509_ (.A(net451),
    .B(net1281),
    .Y(_05422_));
 sky130_fd_sc_hd__mux2_1 _10510_ (.A0(\core.registers[28][10] ),
    .A1(\core.registers[29][10] ),
    .S(net1405),
    .X(_05423_));
 sky130_fd_sc_hd__a221o_1 _10511_ (.A1(net1690),
    .A2(\core.registers[30][10] ),
    .B1(\core.registers[31][10] ),
    .B2(net1405),
    .C1(net1707),
    .X(_05424_));
 sky130_fd_sc_hd__o21a_1 _10512_ (.A1(net1872),
    .A2(_05423_),
    .B1(_05424_),
    .X(_05425_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(\core.registers[14][10] ),
    .A1(\core.registers[15][10] ),
    .S(net1404),
    .X(_05426_));
 sky130_fd_sc_hd__mux2_1 _10514_ (.A0(\core.registers[12][10] ),
    .A1(\core.registers[13][10] ),
    .S(net1404),
    .X(_05427_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(_05426_),
    .A1(_05427_),
    .S(net1472),
    .X(_05428_));
 sky130_fd_sc_hd__mux2_1 _10516_ (.A0(_05425_),
    .A1(_05428_),
    .S(net1716),
    .X(_05429_));
 sky130_fd_sc_hd__a22o_1 _10517_ (.A1(net1690),
    .A2(\core.registers[26][10] ),
    .B1(\core.registers[27][10] ),
    .B2(net1405),
    .X(_05430_));
 sky130_fd_sc_hd__mux2_1 _10518_ (.A0(\core.registers[24][10] ),
    .A1(\core.registers[25][10] ),
    .S(net1405),
    .X(_05431_));
 sky130_fd_sc_hd__mux2_1 _10519_ (.A0(_05430_),
    .A1(_05431_),
    .S(net1707),
    .X(_05432_));
 sky130_fd_sc_hd__or2_1 _10520_ (.A(\core.registers[9][10] ),
    .B(net1377),
    .X(_05433_));
 sky130_fd_sc_hd__o21a_1 _10521_ (.A1(\core.registers[8][10] ),
    .A2(net1404),
    .B1(net1707),
    .X(_05434_));
 sky130_fd_sc_hd__a22o_1 _10522_ (.A1(net1690),
    .A2(\core.registers[10][10] ),
    .B1(\core.registers[11][10] ),
    .B2(net1404),
    .X(_05435_));
 sky130_fd_sc_hd__a221o_1 _10523_ (.A1(_05433_),
    .A2(_05434_),
    .B1(_05435_),
    .B2(net1872),
    .C1(net1856),
    .X(_05436_));
 sky130_fd_sc_hd__o21a_1 _10524_ (.A1(net1716),
    .A2(_05432_),
    .B1(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__mux2_2 _10525_ (.A0(_05429_),
    .A1(_05437_),
    .S(_04420_),
    .X(_05438_));
 sky130_fd_sc_hd__o22a_1 _10526_ (.A1(net1689),
    .A2(\core.registers[23][10] ),
    .B1(net1406),
    .B2(\core.registers[22][10] ),
    .X(_05439_));
 sky130_fd_sc_hd__or3_1 _10527_ (.A(net1689),
    .B(\core.registers[19][10] ),
    .C(net1451),
    .X(_05440_));
 sky130_fd_sc_hd__o221a_1 _10528_ (.A1(\core.registers[18][10] ),
    .A2(net1334),
    .B1(_05439_),
    .B2(net1438),
    .C1(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__mux4_1 _10529_ (.A0(\core.registers[16][10] ),
    .A1(\core.registers[17][10] ),
    .A2(\core.registers[20][10] ),
    .A3(\core.registers[21][10] ),
    .S0(net1406),
    .S1(net1452),
    .X(_05442_));
 sky130_fd_sc_hd__mux2_1 _10530_ (.A0(_05441_),
    .A1(_05442_),
    .S(net1472),
    .X(_05443_));
 sky130_fd_sc_hd__o22a_1 _10531_ (.A1(net1694),
    .A2(\core.registers[7][10] ),
    .B1(net1414),
    .B2(\core.registers[6][10] ),
    .X(_05444_));
 sky130_fd_sc_hd__or3_1 _10532_ (.A(net1689),
    .B(\core.registers[3][10] ),
    .C(net1452),
    .X(_05445_));
 sky130_fd_sc_hd__o221a_1 _10533_ (.A1(\core.registers[2][10] ),
    .A2(net1334),
    .B1(_05444_),
    .B2(net1438),
    .C1(_05445_),
    .X(_05446_));
 sky130_fd_sc_hd__mux4_1 _10534_ (.A0(\core.registers[0][10] ),
    .A1(\core.registers[1][10] ),
    .A2(\core.registers[4][10] ),
    .A3(\core.registers[5][10] ),
    .S0(net1414),
    .S1(net1451),
    .X(_05447_));
 sky130_fd_sc_hd__mux2_1 _10535_ (.A0(_05446_),
    .A1(_05447_),
    .S(net1473),
    .X(_05448_));
 sky130_fd_sc_hd__mux2_1 _10536_ (.A0(_05443_),
    .A1(_05448_),
    .S(net1462),
    .X(_05449_));
 sky130_fd_sc_hd__mux2_2 _10537_ (.A0(_05438_),
    .A1(_05449_),
    .S(net1488),
    .X(_05450_));
 sky130_fd_sc_hd__a22o_4 _10538_ (.A1(net1071),
    .A2(_05387_),
    .B1(_05450_),
    .B2(net1066),
    .X(_05451_));
 sky130_fd_sc_hd__o21ba_4 _10539_ (.A1(net1289),
    .A2(_05451_),
    .B1_N(_05422_),
    .X(_05452_));
 sky130_fd_sc_hd__and3_1 _10540_ (.A(_05419_),
    .B(_05420_),
    .C(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__a21o_2 _10541_ (.A1(_05419_),
    .A2(_05420_),
    .B1(_05452_),
    .X(_05454_));
 sky130_fd_sc_hd__xnor2_4 _10542_ (.A(_05421_),
    .B(_05452_),
    .Y(_05455_));
 sky130_fd_sc_hd__a221o_1 _10543_ (.A1(\core.pipe1_resultRegister[9] ),
    .A2(_04498_),
    .B1(net1270),
    .B2(\core.pipe1_csrData[9] ),
    .C1(net1187),
    .X(_05456_));
 sky130_fd_sc_hd__or2_1 _10544_ (.A(\core.pipe1_loadResult[9] ),
    .B(net1759),
    .X(_05457_));
 sky130_fd_sc_hd__mux2_8 _10545_ (.A0(net170),
    .A1(net142),
    .S(net1805),
    .X(_05458_));
 sky130_fd_sc_hd__o32a_1 _10546_ (.A1(net1676),
    .A2(net1654),
    .A3(_05458_),
    .B1(net1659),
    .B2(\coreWBInterface.readDataBuffered[9] ),
    .X(_05459_));
 sky130_fd_sc_hd__o21ai_1 _10547_ (.A1(net1814),
    .A2(_05459_),
    .B1(_05457_),
    .Y(_05460_));
 sky130_fd_sc_hd__a2111o_2 _10548_ (.A1(_04524_),
    .A2(_04548_),
    .B1(_04933_),
    .C1(_05460_),
    .D1(net1809),
    .X(_05461_));
 sky130_fd_sc_hd__inv_2 _10549_ (.A(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__mux2_8 _10550_ (.A0(net115),
    .A1(net150),
    .S(net1805),
    .X(_05463_));
 sky130_fd_sc_hd__o32a_1 _10551_ (.A1(net1674),
    .A2(net1652),
    .A3(_05463_),
    .B1(net1658),
    .B2(\coreWBInterface.readDataBuffered[17] ),
    .X(_05464_));
 sky130_fd_sc_hd__mux2_4 _10552_ (.A0(\core.pipe1_loadResult[17] ),
    .A1(_05464_),
    .S(net1758),
    .X(_05465_));
 sky130_fd_sc_hd__nand4_2 _10553_ (.A(_04549_),
    .B(_04558_),
    .C(_04943_),
    .D(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__a21o_1 _10554_ (.A1(_04945_),
    .A2(_05466_),
    .B1(_04551_),
    .X(_05467_));
 sky130_fd_sc_hd__mux2_8 _10555_ (.A0(net124),
    .A1(net159),
    .S(net1805),
    .X(_05468_));
 sky130_fd_sc_hd__o32a_1 _10556_ (.A1(net1673),
    .A2(net1660),
    .A3(_05468_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[25] ),
    .X(_05469_));
 sky130_fd_sc_hd__mux2_4 _10557_ (.A0(\core.pipe1_loadResult[25] ),
    .A1(_05469_),
    .S(net1757),
    .X(_05470_));
 sky130_fd_sc_hd__nand2_1 _10558_ (.A(net1233),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__a21o_1 _10559_ (.A1(_04950_),
    .A2(_05471_),
    .B1(_04582_),
    .X(_05472_));
 sky130_fd_sc_hd__a32o_2 _10560_ (.A1(_04948_),
    .A2(_05467_),
    .A3(_05472_),
    .B1(_05461_),
    .B2(_04937_),
    .X(_05473_));
 sky130_fd_sc_hd__nand2_1 _10561_ (.A(net1191),
    .B(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__a22o_2 _10562_ (.A1(\core.pipe1_resultRegister[9] ),
    .A2(net1271),
    .B1(_05456_),
    .B2(_05474_),
    .X(_05475_));
 sky130_fd_sc_hd__mux2_1 _10563_ (.A0(\core.registers[8][9] ),
    .A1(\core.registers[9][9] ),
    .S(net1525),
    .X(_05476_));
 sky130_fd_sc_hd__a221o_1 _10564_ (.A1(net1722),
    .A2(\core.registers[10][9] ),
    .B1(\core.registers[11][9] ),
    .B2(net1525),
    .C1(net1603),
    .X(_05477_));
 sky130_fd_sc_hd__o21a_1 _10565_ (.A1(net1617),
    .A2(_05476_),
    .B1(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__or2_1 _10566_ (.A(\core.registers[13][9] ),
    .B(net1496),
    .X(_05479_));
 sky130_fd_sc_hd__o211a_1 _10567_ (.A1(\core.registers[12][9] ),
    .A2(net1526),
    .B1(_05479_),
    .C1(net1737),
    .X(_05480_));
 sky130_fd_sc_hd__a31o_1 _10568_ (.A1(net1842),
    .A2(net1724),
    .A3(\core.registers[14][9] ),
    .B1(net1745),
    .X(_05481_));
 sky130_fd_sc_hd__a31o_1 _10569_ (.A1(net1842),
    .A2(\core.registers[15][9] ),
    .A3(net1525),
    .B1(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__o221a_1 _10570_ (.A1(net1833),
    .A2(_05478_),
    .B1(_05480_),
    .B2(_05482_),
    .C1(net1749),
    .X(_05483_));
 sky130_fd_sc_hd__or2_1 _10571_ (.A(\core.registers[25][9] ),
    .B(net1497),
    .X(_05484_));
 sky130_fd_sc_hd__o211a_1 _10572_ (.A1(\core.registers[24][9] ),
    .A2(net1532),
    .B1(_05484_),
    .C1(net1737),
    .X(_05485_));
 sky130_fd_sc_hd__a31o_1 _10573_ (.A1(net1842),
    .A2(net1724),
    .A3(\core.registers[26][9] ),
    .B1(net1833),
    .X(_05486_));
 sky130_fd_sc_hd__a311o_1 _10574_ (.A1(net1842),
    .A2(\core.registers[27][9] ),
    .A3(net1532),
    .B1(_05485_),
    .C1(_05486_),
    .X(_05487_));
 sky130_fd_sc_hd__or2_1 _10575_ (.A(\core.registers[29][9] ),
    .B(net1497),
    .X(_05488_));
 sky130_fd_sc_hd__o211a_1 _10576_ (.A1(\core.registers[28][9] ),
    .A2(net1532),
    .B1(_05488_),
    .C1(net1738),
    .X(_05489_));
 sky130_fd_sc_hd__a31o_1 _10577_ (.A1(net1840),
    .A2(net1725),
    .A3(\core.registers[30][9] ),
    .B1(net1745),
    .X(_05490_));
 sky130_fd_sc_hd__a311o_1 _10578_ (.A1(net1840),
    .A2(\core.registers[31][9] ),
    .A3(net1532),
    .B1(_05489_),
    .C1(_05490_),
    .X(_05491_));
 sky130_fd_sc_hd__a31o_1 _10579_ (.A1(net1830),
    .A2(_05487_),
    .A3(_05491_),
    .B1(net1632),
    .X(_05492_));
 sky130_fd_sc_hd__mux2_1 _10580_ (.A0(\core.registers[0][9] ),
    .A1(\core.registers[1][9] ),
    .S(net1532),
    .X(_05493_));
 sky130_fd_sc_hd__o221a_1 _10581_ (.A1(net1724),
    .A2(\core.registers[3][9] ),
    .B1(net1533),
    .B2(\core.registers[2][9] ),
    .C1(net1619),
    .X(_05494_));
 sky130_fd_sc_hd__a211o_1 _10582_ (.A1(net1604),
    .A2(_05493_),
    .B1(_05494_),
    .C1(net1588),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(\core.registers[4][9] ),
    .A1(\core.registers[5][9] ),
    .S(net1532),
    .X(_05496_));
 sky130_fd_sc_hd__mux2_1 _10584_ (.A0(\core.registers[6][9] ),
    .A1(\core.registers[7][9] ),
    .S(net1533),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(_05496_),
    .A1(_05497_),
    .S(net1619),
    .X(_05498_));
 sky130_fd_sc_hd__o211a_1 _10586_ (.A1(net1577),
    .A2(_05498_),
    .B1(_05495_),
    .C1(net1568),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _10587_ (.A0(\core.registers[16][9] ),
    .A1(\core.registers[17][9] ),
    .S(net1532),
    .X(_05500_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(\core.registers[18][9] ),
    .A1(\core.registers[19][9] ),
    .S(net1526),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_1 _10589_ (.A0(_05500_),
    .A1(_05501_),
    .S(net1617),
    .X(_05502_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(\core.registers[20][9] ),
    .A1(\core.registers[21][9] ),
    .S(net1532),
    .X(_05503_));
 sky130_fd_sc_hd__o221a_1 _10591_ (.A1(net1722),
    .A2(\core.registers[23][9] ),
    .B1(net1525),
    .B2(\core.registers[22][9] ),
    .C1(net1617),
    .X(_05504_));
 sky130_fd_sc_hd__a211o_1 _10592_ (.A1(net1603),
    .A2(_05503_),
    .B1(_05504_),
    .C1(net1577),
    .X(_05505_));
 sky130_fd_sc_hd__o211a_1 _10593_ (.A1(net1588),
    .A2(_05502_),
    .B1(_05505_),
    .C1(net1572),
    .X(_05506_));
 sky130_fd_sc_hd__o32a_1 _10594_ (.A1(net1636),
    .A2(_05499_),
    .A3(_05506_),
    .B1(_05483_),
    .B2(_05492_),
    .X(_05507_));
 sky130_fd_sc_hd__o21a_4 _10595_ (.A1(net1158),
    .A2(_05507_),
    .B1(net1264),
    .X(_05508_));
 sky130_fd_sc_hd__o211a_1 _10596_ (.A1(net1156),
    .A2(net965),
    .B1(_05508_),
    .C1(_04482_),
    .X(_05509_));
 sky130_fd_sc_hd__a21o_1 _10597_ (.A1(\core.pipe0_currentInstruction[29] ),
    .A2(net1241),
    .B1(_04478_),
    .X(_05510_));
 sky130_fd_sc_hd__a21oi_2 _10598_ (.A1(_04414_),
    .A2(_04478_),
    .B1(net1289),
    .Y(_05511_));
 sky130_fd_sc_hd__o21ai_4 _10599_ (.A1(_05509_),
    .A2(_05510_),
    .B1(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__nor2_2 _10600_ (.A(net481),
    .B(net1281),
    .Y(_05513_));
 sky130_fd_sc_hd__a21o_1 _10601_ (.A1(\core.registers[20][9] ),
    .A2(net1375),
    .B1(net1433),
    .X(_05514_));
 sky130_fd_sc_hd__a21o_1 _10602_ (.A1(\core.registers[21][9] ),
    .A2(net1402),
    .B1(_05514_),
    .X(_05515_));
 sky130_fd_sc_hd__or2_1 _10603_ (.A(\core.registers[16][9] ),
    .B(net1332),
    .X(_05516_));
 sky130_fd_sc_hd__o31a_1 _10604_ (.A1(\core.registers[17][9] ),
    .A2(net1449),
    .A3(net1375),
    .B1(net1469),
    .X(_05517_));
 sky130_fd_sc_hd__o22a_1 _10605_ (.A1(net1685),
    .A2(\core.registers[23][9] ),
    .B1(net1396),
    .B2(\core.registers[22][9] ),
    .X(_05518_));
 sky130_fd_sc_hd__o31a_1 _10606_ (.A1(net1685),
    .A2(\core.registers[19][9] ),
    .A3(net1449),
    .B1(net1481),
    .X(_05519_));
 sky130_fd_sc_hd__o221a_1 _10607_ (.A1(\core.registers[18][9] ),
    .A2(net1332),
    .B1(_05518_),
    .B2(net1436),
    .C1(_05519_),
    .X(_05520_));
 sky130_fd_sc_hd__a311o_1 _10608_ (.A1(_05515_),
    .A2(_05516_),
    .A3(_05517_),
    .B1(_05520_),
    .C1(net1461),
    .X(_05521_));
 sky130_fd_sc_hd__a21o_1 _10609_ (.A1(\core.registers[4][9] ),
    .A2(net1375),
    .B1(net1437),
    .X(_05522_));
 sky130_fd_sc_hd__a21o_1 _10610_ (.A1(\core.registers[5][9] ),
    .A2(net1402),
    .B1(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__or3_1 _10611_ (.A(\core.registers[1][9] ),
    .B(net1450),
    .C(net1375),
    .X(_05524_));
 sky130_fd_sc_hd__o211a_1 _10612_ (.A1(\core.registers[0][9] ),
    .A2(net1332),
    .B1(_05524_),
    .C1(net1471),
    .X(_05525_));
 sky130_fd_sc_hd__o22a_1 _10613_ (.A1(net1688),
    .A2(\core.registers[7][9] ),
    .B1(net1402),
    .B2(\core.registers[6][9] ),
    .X(_05526_));
 sky130_fd_sc_hd__o31a_1 _10614_ (.A1(net1688),
    .A2(\core.registers[3][9] ),
    .A3(net1449),
    .B1(net1482),
    .X(_05527_));
 sky130_fd_sc_hd__o221a_1 _10615_ (.A1(\core.registers[2][9] ),
    .A2(net1332),
    .B1(_05526_),
    .B2(net1435),
    .C1(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__a211o_1 _10616_ (.A1(_05523_),
    .A2(_05525_),
    .B1(_05528_),
    .C1(net1464),
    .X(_05529_));
 sky130_fd_sc_hd__a21o_1 _10617_ (.A1(_05521_),
    .A2(_05529_),
    .B1(net1490),
    .X(_05530_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(\core.registers[8][9] ),
    .A1(\core.registers[9][9] ),
    .S(net1396),
    .X(_05531_));
 sky130_fd_sc_hd__mux2_1 _10619_ (.A0(\core.registers[10][9] ),
    .A1(\core.registers[11][9] ),
    .S(net1396),
    .X(_05532_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(_05531_),
    .A1(_05532_),
    .S(net1481),
    .X(_05533_));
 sky130_fd_sc_hd__mux2_1 _10621_ (.A0(\core.registers[12][9] ),
    .A1(\core.registers[13][9] ),
    .S(net1397),
    .X(_05534_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(\core.registers[14][9] ),
    .A1(\core.registers[15][9] ),
    .S(net1396),
    .X(_05535_));
 sky130_fd_sc_hd__mux2_1 _10623_ (.A0(_05534_),
    .A1(_05535_),
    .S(net1481),
    .X(_05536_));
 sky130_fd_sc_hd__o22a_1 _10624_ (.A1(net1863),
    .A2(_05533_),
    .B1(_05536_),
    .B2(net1436),
    .X(_05537_));
 sky130_fd_sc_hd__mux2_1 _10625_ (.A0(\core.registers[28][9] ),
    .A1(\core.registers[29][9] ),
    .S(net1402),
    .X(_05538_));
 sky130_fd_sc_hd__a221o_1 _10626_ (.A1(net1688),
    .A2(\core.registers[30][9] ),
    .B1(\core.registers[31][9] ),
    .B2(net1402),
    .C1(net1471),
    .X(_05539_));
 sky130_fd_sc_hd__o211a_1 _10627_ (.A1(net1482),
    .A2(_05538_),
    .B1(_05539_),
    .C1(net1863),
    .X(_05540_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(\core.registers[24][9] ),
    .A1(\core.registers[25][9] ),
    .S(net1402),
    .X(_05541_));
 sky130_fd_sc_hd__or2_1 _10629_ (.A(net1482),
    .B(_05541_),
    .X(_05542_));
 sky130_fd_sc_hd__a221o_1 _10630_ (.A1(net1688),
    .A2(\core.registers[26][9] ),
    .B1(\core.registers[27][9] ),
    .B2(net1402),
    .C1(net1471),
    .X(_05543_));
 sky130_fd_sc_hd__a31o_1 _10631_ (.A1(net1715),
    .A2(_05542_),
    .A3(_05543_),
    .B1(net1461),
    .X(_05544_));
 sky130_fd_sc_hd__o22a_1 _10632_ (.A1(net1464),
    .A2(_05537_),
    .B1(_05540_),
    .B2(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__o21a_2 _10633_ (.A1(net1486),
    .A2(_05545_),
    .B1(_05530_),
    .X(_05546_));
 sky130_fd_sc_hd__a22o_2 _10634_ (.A1(net1069),
    .A2(net965),
    .B1(_05546_),
    .B2(net1067),
    .X(_05547_));
 sky130_fd_sc_hd__o21bai_4 _10635_ (.A1(net1289),
    .A2(_05547_),
    .B1_N(_05513_),
    .Y(_05548_));
 sky130_fd_sc_hd__inv_2 _10636_ (.A(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__nor2_2 _10637_ (.A(_05512_),
    .B(_05548_),
    .Y(_05550_));
 sky130_fd_sc_hd__xor2_4 _10638_ (.A(_05512_),
    .B(_05548_),
    .X(_05551_));
 sky130_fd_sc_hd__nor3_4 _10639_ (.A(_05368_),
    .B(_05455_),
    .C(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__and2b_1 _10640_ (.A_N(_05364_),
    .B(_05331_),
    .X(_05553_));
 sky130_fd_sc_hd__nand2_1 _10641_ (.A(_05421_),
    .B(_05452_),
    .Y(_05554_));
 sky130_fd_sc_hd__nand2b_2 _10642_ (.A_N(_05548_),
    .B(_05512_),
    .Y(_05555_));
 sky130_fd_sc_hd__o21ai_1 _10643_ (.A1(_05455_),
    .A2(_05555_),
    .B1(_05554_),
    .Y(_05556_));
 sky130_fd_sc_hd__a21o_1 _10644_ (.A1(_05369_),
    .A2(_05556_),
    .B1(_05553_),
    .X(_05557_));
 sky130_fd_sc_hd__or2_1 _10645_ (.A(_05552_),
    .B(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__a221o_1 _10646_ (.A1(net1731),
    .A2(\core.registers[26][7] ),
    .B1(\core.registers[27][7] ),
    .B2(net1551),
    .C1(net1740),
    .X(_05559_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(\core.registers[24][7] ),
    .A1(\core.registers[25][7] ),
    .S(net1551),
    .X(_05560_));
 sky130_fd_sc_hd__o21ai_1 _10648_ (.A1(net1845),
    .A2(_05560_),
    .B1(_05559_),
    .Y(_05561_));
 sky130_fd_sc_hd__a221o_1 _10649_ (.A1(net1732),
    .A2(\core.registers[30][7] ),
    .B1(\core.registers[31][7] ),
    .B2(net1548),
    .C1(net1740),
    .X(_05562_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(\core.registers[28][7] ),
    .A1(\core.registers[29][7] ),
    .S(net1548),
    .X(_05563_));
 sky130_fd_sc_hd__o21a_1 _10651_ (.A1(net1845),
    .A2(_05563_),
    .B1(_05562_),
    .X(_05564_));
 sky130_fd_sc_hd__mux2_1 _10652_ (.A0(\core.registers[12][7] ),
    .A1(\core.registers[13][7] ),
    .S(net1548),
    .X(_05565_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(\core.registers[14][7] ),
    .A1(\core.registers[15][7] ),
    .S(net1548),
    .X(_05566_));
 sky130_fd_sc_hd__mux2_1 _10654_ (.A0(_05565_),
    .A1(_05566_),
    .S(net1626),
    .X(_05567_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(_05564_),
    .A1(_05567_),
    .S(net1750),
    .X(_05568_));
 sky130_fd_sc_hd__or2_1 _10656_ (.A(\core.registers[1][7] ),
    .B(net1501),
    .X(_05569_));
 sky130_fd_sc_hd__or2_1 _10657_ (.A(\core.registers[6][7] ),
    .B(net1561),
    .X(_05570_));
 sky130_fd_sc_hd__or2_1 _10658_ (.A(\core.registers[22][7] ),
    .B(net1552),
    .X(_05571_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(\core.registers[8][7] ),
    .A1(\core.registers[9][7] ),
    .S(net1551),
    .X(_05572_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(\core.registers[10][7] ),
    .A1(\core.registers[11][7] ),
    .S(net1551),
    .X(_05573_));
 sky130_fd_sc_hd__mux2_1 _10661_ (.A0(_05572_),
    .A1(_05573_),
    .S(net1624),
    .X(_05574_));
 sky130_fd_sc_hd__or2_1 _10662_ (.A(net1826),
    .B(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__a21oi_1 _10663_ (.A1(net1826),
    .A2(_05561_),
    .B1(net1834),
    .Y(_05576_));
 sky130_fd_sc_hd__a221o_2 _10664_ (.A1(net1834),
    .A2(_05568_),
    .B1(_05575_),
    .B2(_05576_),
    .C1(net1634),
    .X(_05577_));
 sky130_fd_sc_hd__o211a_1 _10665_ (.A1(net1734),
    .A2(\core.registers[7][7] ),
    .B1(net1627),
    .C1(_05570_),
    .X(_05578_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\core.registers[4][7] ),
    .A1(\core.registers[5][7] ),
    .S(net1554),
    .X(_05579_));
 sky130_fd_sc_hd__a211o_1 _10667_ (.A1(net1610),
    .A2(_05579_),
    .B1(_05578_),
    .C1(net1581),
    .X(_05580_));
 sky130_fd_sc_hd__o211a_1 _10668_ (.A1(\core.registers[0][7] ),
    .A2(net1561),
    .B1(_05569_),
    .C1(net1607),
    .X(_05581_));
 sky130_fd_sc_hd__mux2_1 _10669_ (.A0(\core.registers[2][7] ),
    .A1(\core.registers[3][7] ),
    .S(net1554),
    .X(_05582_));
 sky130_fd_sc_hd__a211o_1 _10670_ (.A1(net1624),
    .A2(_05582_),
    .B1(_05581_),
    .C1(net1592),
    .X(_05583_));
 sky130_fd_sc_hd__mux2_1 _10671_ (.A0(\core.registers[16][7] ),
    .A1(\core.registers[17][7] ),
    .S(net1554),
    .X(_05584_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(\core.registers[18][7] ),
    .A1(\core.registers[19][7] ),
    .S(net1554),
    .X(_05585_));
 sky130_fd_sc_hd__mux2_1 _10673_ (.A0(_05584_),
    .A1(_05585_),
    .S(net1624),
    .X(_05586_));
 sky130_fd_sc_hd__o211a_1 _10674_ (.A1(net1731),
    .A2(\core.registers[23][7] ),
    .B1(net1624),
    .C1(_05571_),
    .X(_05587_));
 sky130_fd_sc_hd__mux2_1 _10675_ (.A0(\core.registers[20][7] ),
    .A1(\core.registers[21][7] ),
    .S(net1552),
    .X(_05588_));
 sky130_fd_sc_hd__a211o_1 _10676_ (.A1(net1610),
    .A2(_05588_),
    .B1(_05587_),
    .C1(net1581),
    .X(_05589_));
 sky130_fd_sc_hd__o211a_1 _10677_ (.A1(net1592),
    .A2(_05586_),
    .B1(_05589_),
    .C1(net1574),
    .X(_05590_));
 sky130_fd_sc_hd__a311o_1 _10678_ (.A1(net1570),
    .A2(_05580_),
    .A3(_05583_),
    .B1(_05590_),
    .C1(net1638),
    .X(_05591_));
 sky130_fd_sc_hd__a21o_2 _10679_ (.A1(_05577_),
    .A2(_05591_),
    .B1(net1160),
    .X(_05592_));
 sky130_fd_sc_hd__a22o_1 _10680_ (.A1(\core.pipe1_resultRegister[7] ),
    .A2(net1240),
    .B1(net1268),
    .B2(\core.pipe1_csrData[7] ),
    .X(_05593_));
 sky130_fd_sc_hd__a21o_1 _10681_ (.A1(net1189),
    .A2(_04591_),
    .B1(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__o211a_4 _10682_ (.A1(net1155),
    .A2(net1135),
    .B1(_05592_),
    .C1(net1265),
    .X(_05595_));
 sky130_fd_sc_hd__or2_1 _10683_ (.A(\core.pipe0_currentInstruction[27] ),
    .B(_04484_),
    .X(_05596_));
 sky130_fd_sc_hd__o211a_2 _10684_ (.A1(net1194),
    .A2(_05595_),
    .B1(_05596_),
    .C1(net1283),
    .X(_05597_));
 sky130_fd_sc_hd__nor2_1 _10685_ (.A(net479),
    .B(net1283),
    .Y(_05598_));
 sky130_fd_sc_hd__o22a_1 _10686_ (.A1(net1698),
    .A2(\core.registers[23][7] ),
    .B1(net1421),
    .B2(\core.registers[22][7] ),
    .X(_05599_));
 sky130_fd_sc_hd__or3_1 _10687_ (.A(net1698),
    .B(\core.registers[19][7] ),
    .C(net1455),
    .X(_05600_));
 sky130_fd_sc_hd__o221a_1 _10688_ (.A1(\core.registers[18][7] ),
    .A2(net1335),
    .B1(_05599_),
    .B2(net1441),
    .C1(_05600_),
    .X(_05601_));
 sky130_fd_sc_hd__mux4_1 _10689_ (.A0(\core.registers[16][7] ),
    .A1(\core.registers[17][7] ),
    .A2(\core.registers[20][7] ),
    .A3(\core.registers[21][7] ),
    .S0(net1420),
    .S1(net1455),
    .X(_05602_));
 sky130_fd_sc_hd__mux2_1 _10690_ (.A0(_05601_),
    .A1(_05602_),
    .S(net1476),
    .X(_05603_));
 sky130_fd_sc_hd__o22a_1 _10691_ (.A1(net1697),
    .A2(\core.registers[7][7] ),
    .B1(net1427),
    .B2(\core.registers[6][7] ),
    .X(_05604_));
 sky130_fd_sc_hd__or3_1 _10692_ (.A(net1698),
    .B(\core.registers[3][7] ),
    .C(net1455),
    .X(_05605_));
 sky130_fd_sc_hd__o221a_1 _10693_ (.A1(\core.registers[2][7] ),
    .A2(net1335),
    .B1(_05604_),
    .B2(net1441),
    .C1(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__mux4_1 _10694_ (.A0(\core.registers[0][7] ),
    .A1(\core.registers[1][7] ),
    .A2(\core.registers[4][7] ),
    .A3(\core.registers[5][7] ),
    .S0(net1420),
    .S1(net1455),
    .X(_05607_));
 sky130_fd_sc_hd__mux2_1 _10695_ (.A0(_05606_),
    .A1(_05607_),
    .S(net1474),
    .X(_05608_));
 sky130_fd_sc_hd__mux2_2 _10696_ (.A0(_05603_),
    .A1(_05608_),
    .S(net1463),
    .X(_05609_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(\core.registers[10][7] ),
    .A1(\core.registers[11][7] ),
    .S(net1419),
    .X(_05610_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(\core.registers[8][7] ),
    .A1(\core.registers[9][7] ),
    .S(net1419),
    .X(_05611_));
 sky130_fd_sc_hd__mux2_1 _10699_ (.A0(_05610_),
    .A1(_05611_),
    .S(net1474),
    .X(_05612_));
 sky130_fd_sc_hd__nor2_1 _10700_ (.A(net1858),
    .B(_05612_),
    .Y(_05613_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(\core.registers[24][7] ),
    .A1(\core.registers[25][7] ),
    .S(net1419),
    .X(_05614_));
 sky130_fd_sc_hd__a221o_1 _10702_ (.A1(net1698),
    .A2(\core.registers[26][7] ),
    .B1(\core.registers[27][7] ),
    .B2(net1419),
    .C1(net1709),
    .X(_05615_));
 sky130_fd_sc_hd__o21ai_1 _10703_ (.A1(net1875),
    .A2(_05614_),
    .B1(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__a211o_1 _10704_ (.A1(net1859),
    .A2(_05616_),
    .B1(_05613_),
    .C1(net1864),
    .X(_05617_));
 sky130_fd_sc_hd__or2_1 _10705_ (.A(\core.registers[13][7] ),
    .B(net1376),
    .X(_05618_));
 sky130_fd_sc_hd__o21a_1 _10706_ (.A1(\core.registers[12][7] ),
    .A2(net1416),
    .B1(net1709),
    .X(_05619_));
 sky130_fd_sc_hd__a22o_1 _10707_ (.A1(net1695),
    .A2(\core.registers[14][7] ),
    .B1(\core.registers[15][7] ),
    .B2(net1416),
    .X(_05620_));
 sky130_fd_sc_hd__a221o_1 _10708_ (.A1(_05618_),
    .A2(_05619_),
    .B1(_05620_),
    .B2(net1876),
    .C1(net1858),
    .X(_05621_));
 sky130_fd_sc_hd__a221o_1 _10709_ (.A1(net1695),
    .A2(\core.registers[30][7] ),
    .B1(\core.registers[31][7] ),
    .B2(net1416),
    .C1(net1709),
    .X(_05622_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(\core.registers[28][7] ),
    .A1(\core.registers[29][7] ),
    .S(net1416),
    .X(_05623_));
 sky130_fd_sc_hd__o21a_1 _10711_ (.A1(net1875),
    .A2(_05623_),
    .B1(_05622_),
    .X(_05624_));
 sky130_fd_sc_hd__o211a_1 _10712_ (.A1(net1717),
    .A2(_05624_),
    .B1(_05621_),
    .C1(net1864),
    .X(_05625_));
 sky130_fd_sc_hd__nor2_1 _10713_ (.A(net1487),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__o2bb2a_4 _10714_ (.A1_N(_05617_),
    .A2_N(_05626_),
    .B1(net1491),
    .B2(_05609_),
    .X(_05627_));
 sky130_fd_sc_hd__a22o_4 _10715_ (.A1(net1070),
    .A2(net1135),
    .B1(_05627_),
    .B2(net1066),
    .X(_05628_));
 sky130_fd_sc_hd__o21ba_4 _10716_ (.A1(net1288),
    .A2(_05628_),
    .B1_N(_05598_),
    .X(_05629_));
 sky130_fd_sc_hd__and2_4 _10717_ (.A(_05597_),
    .B(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__nor2_4 _10718_ (.A(_05597_),
    .B(_05629_),
    .Y(_05631_));
 sky130_fd_sc_hd__inv_2 _10719_ (.A(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__nor2_8 _10720_ (.A(_05630_),
    .B(_05631_),
    .Y(_05633_));
 sky130_fd_sc_hd__a22o_1 _10721_ (.A1(\core.pipe1_resultRegister[6] ),
    .A2(net1239),
    .B1(net1268),
    .B2(\core.pipe1_csrData[6] ),
    .X(_05634_));
 sky130_fd_sc_hd__a21o_1 _10722_ (.A1(net1807),
    .A2(_05198_),
    .B1(net1811),
    .X(_05635_));
 sky130_fd_sc_hd__o211ai_2 _10723_ (.A1(_04558_),
    .A2(_05203_),
    .B1(_05635_),
    .C1(_05197_),
    .Y(_05636_));
 sky130_fd_sc_hd__mux2_8 _10724_ (.A0(net167),
    .A1(net138),
    .S(net1805),
    .X(_05637_));
 sky130_fd_sc_hd__o32ai_4 _10725_ (.A1(net1675),
    .A2(net1655),
    .A3(_05637_),
    .B1(net1659),
    .B2(\coreWBInterface.readDataBuffered[6] ),
    .Y(_05638_));
 sky130_fd_sc_hd__nor2_1 _10726_ (.A(net1812),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__a211o_1 _10727_ (.A1(\core.pipe1_loadResult[6] ),
    .A2(net1812),
    .B1(_04572_),
    .C1(_05639_),
    .X(_05640_));
 sky130_fd_sc_hd__a31o_4 _10728_ (.A1(net1189),
    .A2(_05636_),
    .A3(_05640_),
    .B1(_05634_),
    .X(_05641_));
 sky130_fd_sc_hd__a221o_1 _10729_ (.A1(net1731),
    .A2(\core.registers[26][6] ),
    .B1(\core.registers[27][6] ),
    .B2(net1553),
    .C1(net1740),
    .X(_05642_));
 sky130_fd_sc_hd__mux2_1 _10730_ (.A0(\core.registers[24][6] ),
    .A1(\core.registers[25][6] ),
    .S(net1553),
    .X(_05643_));
 sky130_fd_sc_hd__o21ai_1 _10731_ (.A1(net1845),
    .A2(_05643_),
    .B1(_05642_),
    .Y(_05644_));
 sky130_fd_sc_hd__a221o_1 _10732_ (.A1(net1732),
    .A2(\core.registers[30][6] ),
    .B1(\core.registers[31][6] ),
    .B2(net1550),
    .C1(net1740),
    .X(_05645_));
 sky130_fd_sc_hd__mux2_1 _10733_ (.A0(\core.registers[28][6] ),
    .A1(\core.registers[29][6] ),
    .S(net1550),
    .X(_05646_));
 sky130_fd_sc_hd__o21a_1 _10734_ (.A1(net1845),
    .A2(_05646_),
    .B1(_05645_),
    .X(_05647_));
 sky130_fd_sc_hd__mux2_1 _10735_ (.A0(\core.registers[12][6] ),
    .A1(\core.registers[13][6] ),
    .S(net1550),
    .X(_05648_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(\core.registers[14][6] ),
    .A1(\core.registers[15][6] ),
    .S(net1550),
    .X(_05649_));
 sky130_fd_sc_hd__mux2_1 _10737_ (.A0(_05648_),
    .A1(_05649_),
    .S(net1626),
    .X(_05650_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(_05647_),
    .A1(_05650_),
    .S(net1751),
    .X(_05651_));
 sky130_fd_sc_hd__or2_1 _10739_ (.A(\core.registers[6][6] ),
    .B(net1563),
    .X(_05652_));
 sky130_fd_sc_hd__or2_1 _10740_ (.A(\core.registers[22][6] ),
    .B(net1554),
    .X(_05653_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(\core.registers[8][6] ),
    .A1(\core.registers[9][6] ),
    .S(net1552),
    .X(_05654_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(\core.registers[10][6] ),
    .A1(\core.registers[11][6] ),
    .S(net1551),
    .X(_05655_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(_05654_),
    .A1(_05655_),
    .S(net1624),
    .X(_05656_));
 sky130_fd_sc_hd__or2_1 _10744_ (.A(net1826),
    .B(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__a21oi_1 _10745_ (.A1(net1826),
    .A2(_05644_),
    .B1(net1834),
    .Y(_05658_));
 sky130_fd_sc_hd__a221o_4 _10746_ (.A1(net1834),
    .A2(_05651_),
    .B1(_05657_),
    .B2(_05658_),
    .C1(net1634),
    .X(_05659_));
 sky130_fd_sc_hd__o211a_1 _10747_ (.A1(net1734),
    .A2(\core.registers[7][6] ),
    .B1(net1627),
    .C1(_05652_),
    .X(_05660_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(\core.registers[4][6] ),
    .A1(\core.registers[5][6] ),
    .S(net1563),
    .X(_05661_));
 sky130_fd_sc_hd__a211o_1 _10749_ (.A1(net1607),
    .A2(_05661_),
    .B1(_05660_),
    .C1(net1582),
    .X(_05662_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(\core.registers[0][6] ),
    .A1(\core.registers[1][6] ),
    .S(net1564),
    .X(_05663_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(\core.registers[2][6] ),
    .A1(\core.registers[3][6] ),
    .S(net1564),
    .X(_05664_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(_05663_),
    .A1(_05664_),
    .S(net1628),
    .X(_05665_));
 sky130_fd_sc_hd__o211a_2 _10753_ (.A1(net1592),
    .A2(_05665_),
    .B1(_05662_),
    .C1(net1570),
    .X(_05666_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(\core.registers[16][6] ),
    .A1(\core.registers[17][6] ),
    .S(net1554),
    .X(_05667_));
 sky130_fd_sc_hd__mux2_1 _10755_ (.A0(\core.registers[18][6] ),
    .A1(\core.registers[19][6] ),
    .S(net1554),
    .X(_05668_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(_05667_),
    .A1(_05668_),
    .S(net1625),
    .X(_05669_));
 sky130_fd_sc_hd__o211a_1 _10757_ (.A1(net1731),
    .A2(\core.registers[23][6] ),
    .B1(net1625),
    .C1(_05653_),
    .X(_05670_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\core.registers[20][6] ),
    .A1(\core.registers[21][6] ),
    .S(net1554),
    .X(_05671_));
 sky130_fd_sc_hd__a211o_1 _10759_ (.A1(net1610),
    .A2(_05671_),
    .B1(_05670_),
    .C1(net1581),
    .X(_05672_));
 sky130_fd_sc_hd__o211a_2 _10760_ (.A1(net1592),
    .A2(_05669_),
    .B1(_05672_),
    .C1(net1574),
    .X(_05673_));
 sky130_fd_sc_hd__o31a_4 _10761_ (.A1(net1638),
    .A2(_05666_),
    .A3(_05673_),
    .B1(_05659_),
    .X(_05674_));
 sky130_fd_sc_hd__o21a_1 _10762_ (.A1(net1155),
    .A2(net1064),
    .B1(net1265),
    .X(_05675_));
 sky130_fd_sc_hd__o21ai_4 _10763_ (.A1(net1159),
    .A2(_05674_),
    .B1(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__nand2_1 _10764_ (.A(_04484_),
    .B(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__o211a_1 _10765_ (.A1(\core.pipe0_currentInstruction[26] ),
    .A2(_04484_),
    .B1(_05677_),
    .C1(net1283),
    .X(_05678_));
 sky130_fd_sc_hd__nor2_1 _10766_ (.A(net478),
    .B(net1283),
    .Y(_05679_));
 sky130_fd_sc_hd__o22a_1 _10767_ (.A1(net1697),
    .A2(\core.registers[23][6] ),
    .B1(net1421),
    .B2(\core.registers[22][6] ),
    .X(_05680_));
 sky130_fd_sc_hd__or3_1 _10768_ (.A(net1697),
    .B(\core.registers[19][6] ),
    .C(net1455),
    .X(_05681_));
 sky130_fd_sc_hd__o221a_1 _10769_ (.A1(\core.registers[18][6] ),
    .A2(net1335),
    .B1(_05680_),
    .B2(net1441),
    .C1(_05681_),
    .X(_05682_));
 sky130_fd_sc_hd__mux4_1 _10770_ (.A0(\core.registers[16][6] ),
    .A1(\core.registers[17][6] ),
    .A2(\core.registers[20][6] ),
    .A3(\core.registers[21][6] ),
    .S0(net1420),
    .S1(net1455),
    .X(_05683_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(_05682_),
    .A1(_05683_),
    .S(net1474),
    .X(_05684_));
 sky130_fd_sc_hd__o22a_1 _10772_ (.A1(net1700),
    .A2(\core.registers[7][6] ),
    .B1(net1428),
    .B2(\core.registers[6][6] ),
    .X(_05685_));
 sky130_fd_sc_hd__or3_1 _10773_ (.A(net1700),
    .B(\core.registers[3][6] ),
    .C(net1458),
    .X(_05686_));
 sky130_fd_sc_hd__o221a_1 _10774_ (.A1(\core.registers[2][6] ),
    .A2(net1336),
    .B1(_05685_),
    .B2(net1440),
    .C1(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__mux4_1 _10775_ (.A0(\core.registers[0][6] ),
    .A1(\core.registers[1][6] ),
    .A2(\core.registers[4][6] ),
    .A3(\core.registers[5][6] ),
    .S0(net1428),
    .S1(net1457),
    .X(_05688_));
 sky130_fd_sc_hd__mux2_2 _10776_ (.A0(_05687_),
    .A1(_05688_),
    .S(net1475),
    .X(_05689_));
 sky130_fd_sc_hd__mux2_2 _10777_ (.A0(_05684_),
    .A1(_05689_),
    .S(net1463),
    .X(_05690_));
 sky130_fd_sc_hd__mux2_1 _10778_ (.A0(\core.registers[10][6] ),
    .A1(\core.registers[11][6] ),
    .S(net1419),
    .X(_05691_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\core.registers[8][6] ),
    .A1(\core.registers[9][6] ),
    .S(net1419),
    .X(_05692_));
 sky130_fd_sc_hd__mux2_1 _10780_ (.A0(_05691_),
    .A1(_05692_),
    .S(net1474),
    .X(_05693_));
 sky130_fd_sc_hd__nor2_1 _10781_ (.A(net1858),
    .B(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__mux2_1 _10782_ (.A0(\core.registers[24][6] ),
    .A1(\core.registers[25][6] ),
    .S(net1420),
    .X(_05695_));
 sky130_fd_sc_hd__a221o_1 _10783_ (.A1(net1698),
    .A2(\core.registers[26][6] ),
    .B1(\core.registers[27][6] ),
    .B2(net1420),
    .C1(net1709),
    .X(_05696_));
 sky130_fd_sc_hd__o21ai_1 _10784_ (.A1(net1875),
    .A2(_05695_),
    .B1(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__a211o_1 _10785_ (.A1(net1858),
    .A2(_05697_),
    .B1(_05694_),
    .C1(net1864),
    .X(_05698_));
 sky130_fd_sc_hd__or2_1 _10786_ (.A(\core.registers[13][6] ),
    .B(net1376),
    .X(_05699_));
 sky130_fd_sc_hd__o21a_1 _10787_ (.A1(\core.registers[12][6] ),
    .A2(net1418),
    .B1(net1709),
    .X(_05700_));
 sky130_fd_sc_hd__a22o_1 _10788_ (.A1(net1695),
    .A2(\core.registers[14][6] ),
    .B1(\core.registers[15][6] ),
    .B2(net1418),
    .X(_05701_));
 sky130_fd_sc_hd__a221o_1 _10789_ (.A1(_05699_),
    .A2(_05700_),
    .B1(_05701_),
    .B2(net1875),
    .C1(net1858),
    .X(_05702_));
 sky130_fd_sc_hd__mux2_1 _10790_ (.A0(\core.registers[28][6] ),
    .A1(\core.registers[29][6] ),
    .S(net1418),
    .X(_05703_));
 sky130_fd_sc_hd__a221o_1 _10791_ (.A1(net1695),
    .A2(\core.registers[30][6] ),
    .B1(\core.registers[31][6] ),
    .B2(net1418),
    .C1(net1709),
    .X(_05704_));
 sky130_fd_sc_hd__o21a_1 _10792_ (.A1(net1876),
    .A2(_05703_),
    .B1(_05704_),
    .X(_05705_));
 sky130_fd_sc_hd__o211a_1 _10793_ (.A1(net1717),
    .A2(_05705_),
    .B1(_05702_),
    .C1(net1864),
    .X(_05706_));
 sky130_fd_sc_hd__nor2_1 _10794_ (.A(net1487),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__o2bb2a_4 _10795_ (.A1_N(_05698_),
    .A2_N(_05707_),
    .B1(net1491),
    .B2(_05690_),
    .X(_05708_));
 sky130_fd_sc_hd__a22o_4 _10796_ (.A1(net1070),
    .A2(net1064),
    .B1(_05708_),
    .B2(net1066),
    .X(_05709_));
 sky130_fd_sc_hd__o21ba_2 _10797_ (.A1(net1288),
    .A2(_05709_),
    .B1_N(_05679_),
    .X(_05710_));
 sky130_fd_sc_hd__and2_1 _10798_ (.A(_05678_),
    .B(_05710_),
    .X(_05711_));
 sky130_fd_sc_hd__or2_4 _10799_ (.A(_05678_),
    .B(_05710_),
    .X(_05712_));
 sky130_fd_sc_hd__and2b_4 _10800_ (.A_N(_05711_),
    .B(_05712_),
    .X(_05713_));
 sky130_fd_sc_hd__inv_2 _10801_ (.A(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__nand2b_2 _10802_ (.A_N(_05597_),
    .B(_05629_),
    .Y(_05715_));
 sky130_fd_sc_hd__nand2b_2 _10803_ (.A_N(_05678_),
    .B(_05710_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21ai_4 _10804_ (.A1(_05633_),
    .A2(_05716_),
    .B1(_05715_),
    .Y(_05717_));
 sky130_fd_sc_hd__o21bai_2 _10805_ (.A1(_05633_),
    .A2(_05713_),
    .B1_N(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__a22o_1 _10806_ (.A1(\core.pipe1_resultRegister[5] ),
    .A2(net1239),
    .B1(net1269),
    .B2(\core.pipe1_csrData[5] ),
    .X(_05719_));
 sky130_fd_sc_hd__a21o_1 _10807_ (.A1(net1807),
    .A2(_05032_),
    .B1(net1811),
    .X(_05720_));
 sky130_fd_sc_hd__o211ai_2 _10808_ (.A1(_04558_),
    .A2(_05037_),
    .B1(_05720_),
    .C1(_05031_),
    .Y(_05721_));
 sky130_fd_sc_hd__mux2_8 _10809_ (.A0(net162),
    .A1(net137),
    .S(net1805),
    .X(_05722_));
 sky130_fd_sc_hd__o32ai_4 _10810_ (.A1(net1675),
    .A2(net1655),
    .A3(_05722_),
    .B1(net1658),
    .B2(\coreWBInterface.readDataBuffered[5] ),
    .Y(_05723_));
 sky130_fd_sc_hd__nor2_1 _10811_ (.A(net1812),
    .B(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__a211o_1 _10812_ (.A1(\core.pipe1_loadResult[5] ),
    .A2(net1812),
    .B1(_04572_),
    .C1(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__a31o_4 _10813_ (.A1(net1189),
    .A2(_05721_),
    .A3(_05725_),
    .B1(_05719_),
    .X(_05726_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(\core.registers[8][5] ),
    .A1(\core.registers[9][5] ),
    .S(net1560),
    .X(_05727_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(\core.registers[10][5] ),
    .A1(\core.registers[11][5] ),
    .S(net1560),
    .X(_05728_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(\core.registers[24][5] ),
    .A1(\core.registers[25][5] ),
    .S(net1560),
    .X(_05729_));
 sky130_fd_sc_hd__a221o_1 _10817_ (.A1(net1733),
    .A2(\core.registers[26][5] ),
    .B1(\core.registers[27][5] ),
    .B2(net1560),
    .C1(net1742),
    .X(_05730_));
 sky130_fd_sc_hd__or2_1 _10818_ (.A(\core.registers[29][5] ),
    .B(net1501),
    .X(_05731_));
 sky130_fd_sc_hd__o211a_1 _10819_ (.A1(\core.registers[28][5] ),
    .A2(net1558),
    .B1(_05731_),
    .C1(net1742),
    .X(_05732_));
 sky130_fd_sc_hd__a31o_1 _10820_ (.A1(net1846),
    .A2(net1733),
    .A3(\core.registers[30][5] ),
    .B1(net1751),
    .X(_05733_));
 sky130_fd_sc_hd__a31o_1 _10821_ (.A1(net1847),
    .A2(\core.registers[31][5] ),
    .A3(net1558),
    .B1(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__or2_1 _10822_ (.A(\core.registers[1][5] ),
    .B(net1501),
    .X(_05735_));
 sky130_fd_sc_hd__or2_1 _10823_ (.A(\core.registers[6][5] ),
    .B(net1561),
    .X(_05736_));
 sky130_fd_sc_hd__or2_1 _10824_ (.A(\core.registers[17][5] ),
    .B(net1502),
    .X(_05737_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(\core.registers[12][5] ),
    .A1(\core.registers[13][5] ),
    .S(net1559),
    .X(_05738_));
 sky130_fd_sc_hd__mux2_1 _10826_ (.A0(\core.registers[14][5] ),
    .A1(\core.registers[15][5] ),
    .S(net1558),
    .X(_05739_));
 sky130_fd_sc_hd__mux2_1 _10827_ (.A0(_05738_),
    .A1(_05739_),
    .S(net1629),
    .X(_05740_));
 sky130_fd_sc_hd__o221a_1 _10828_ (.A1(_05732_),
    .A2(_05734_),
    .B1(_05740_),
    .B2(net1828),
    .C1(net1835),
    .X(_05741_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(_05727_),
    .A1(_05728_),
    .S(net1627),
    .X(_05742_));
 sky130_fd_sc_hd__o21a_1 _10830_ (.A1(net1846),
    .A2(_05729_),
    .B1(_05730_),
    .X(_05743_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(_05742_),
    .A1(_05743_),
    .S(net1828),
    .X(_05744_));
 sky130_fd_sc_hd__a211o_1 _10832_ (.A1(net1746),
    .A2(_05744_),
    .B1(_05741_),
    .C1(net1634),
    .X(_05745_));
 sky130_fd_sc_hd__o211a_1 _10833_ (.A1(net1733),
    .A2(\core.registers[7][5] ),
    .B1(net1627),
    .C1(_05736_),
    .X(_05746_));
 sky130_fd_sc_hd__mux2_1 _10834_ (.A0(\core.registers[4][5] ),
    .A1(\core.registers[5][5] ),
    .S(net1560),
    .X(_05747_));
 sky130_fd_sc_hd__a211o_1 _10835_ (.A1(net1607),
    .A2(_05747_),
    .B1(_05746_),
    .C1(net1581),
    .X(_05748_));
 sky130_fd_sc_hd__o211a_1 _10836_ (.A1(\core.registers[0][5] ),
    .A2(net1564),
    .B1(_05735_),
    .C1(net1607),
    .X(_05749_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(\core.registers[2][5] ),
    .A1(\core.registers[3][5] ),
    .S(net1562),
    .X(_05750_));
 sky130_fd_sc_hd__a211o_1 _10838_ (.A1(net1627),
    .A2(_05750_),
    .B1(_05749_),
    .C1(net1592),
    .X(_05751_));
 sky130_fd_sc_hd__o211a_1 _10839_ (.A1(\core.registers[16][5] ),
    .A2(net1561),
    .B1(_05737_),
    .C1(net1607),
    .X(_05752_));
 sky130_fd_sc_hd__mux2_1 _10840_ (.A0(\core.registers[18][5] ),
    .A1(\core.registers[19][5] ),
    .S(net1561),
    .X(_05753_));
 sky130_fd_sc_hd__a211o_1 _10841_ (.A1(net1627),
    .A2(_05753_),
    .B1(_05752_),
    .C1(net1593),
    .X(_05754_));
 sky130_fd_sc_hd__mux2_1 _10842_ (.A0(\core.registers[22][5] ),
    .A1(\core.registers[23][5] ),
    .S(net1565),
    .X(_05755_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(\core.registers[20][5] ),
    .A1(\core.registers[21][5] ),
    .S(net1561),
    .X(_05756_));
 sky130_fd_sc_hd__mux2_1 _10844_ (.A0(_05755_),
    .A1(_05756_),
    .S(net1607),
    .X(_05757_));
 sky130_fd_sc_hd__o211a_1 _10845_ (.A1(net1582),
    .A2(_05757_),
    .B1(_05754_),
    .C1(net1574),
    .X(_05758_));
 sky130_fd_sc_hd__a311o_1 _10846_ (.A1(net1570),
    .A2(_05748_),
    .A3(_05751_),
    .B1(_05758_),
    .C1(net1638),
    .X(_05759_));
 sky130_fd_sc_hd__a21o_2 _10847_ (.A1(_05745_),
    .A2(_05759_),
    .B1(net1160),
    .X(_05760_));
 sky130_fd_sc_hd__o211a_4 _10848_ (.A1(net1155),
    .A2(net1059),
    .B1(_05760_),
    .C1(net1265),
    .X(_05761_));
 sky130_fd_sc_hd__or2_1 _10849_ (.A(\core.pipe0_currentInstruction[25] ),
    .B(_04484_),
    .X(_05762_));
 sky130_fd_sc_hd__o211a_2 _10850_ (.A1(net1194),
    .A2(_05761_),
    .B1(_05762_),
    .C1(net1283),
    .X(_05763_));
 sky130_fd_sc_hd__nor2_1 _10851_ (.A(net477),
    .B(net1284),
    .Y(_05764_));
 sky130_fd_sc_hd__o22a_1 _10852_ (.A1(net1699),
    .A2(\core.registers[23][5] ),
    .B1(net1427),
    .B2(\core.registers[22][5] ),
    .X(_05765_));
 sky130_fd_sc_hd__or3_1 _10853_ (.A(net1700),
    .B(\core.registers[19][5] ),
    .C(net1457),
    .X(_05766_));
 sky130_fd_sc_hd__o221a_1 _10854_ (.A1(\core.registers[18][5] ),
    .A2(net1336),
    .B1(_05765_),
    .B2(net1440),
    .C1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__mux4_1 _10855_ (.A0(\core.registers[16][5] ),
    .A1(\core.registers[17][5] ),
    .A2(\core.registers[20][5] ),
    .A3(\core.registers[21][5] ),
    .S0(net1427),
    .S1(net1457),
    .X(_05768_));
 sky130_fd_sc_hd__mux2_1 _10856_ (.A0(_05767_),
    .A1(_05768_),
    .S(net1476),
    .X(_05769_));
 sky130_fd_sc_hd__o22a_1 _10857_ (.A1(net1699),
    .A2(\core.registers[7][5] ),
    .B1(net1427),
    .B2(\core.registers[6][5] ),
    .X(_05770_));
 sky130_fd_sc_hd__or3_1 _10858_ (.A(net1699),
    .B(\core.registers[3][5] ),
    .C(net1457),
    .X(_05771_));
 sky130_fd_sc_hd__o221a_1 _10859_ (.A1(\core.registers[2][5] ),
    .A2(net1335),
    .B1(_05770_),
    .B2(net1441),
    .C1(_05771_),
    .X(_05772_));
 sky130_fd_sc_hd__mux4_1 _10860_ (.A0(\core.registers[0][5] ),
    .A1(\core.registers[1][5] ),
    .A2(\core.registers[4][5] ),
    .A3(\core.registers[5][5] ),
    .S0(net1426),
    .S1(net1457),
    .X(_05773_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(_05772_),
    .A1(_05773_),
    .S(net1476),
    .X(_05774_));
 sky130_fd_sc_hd__mux2_1 _10862_ (.A0(_05769_),
    .A1(_05774_),
    .S(net1463),
    .X(_05775_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(\core.registers[10][5] ),
    .A1(\core.registers[11][5] ),
    .S(net1426),
    .X(_05776_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(\core.registers[8][5] ),
    .A1(\core.registers[9][5] ),
    .S(net1426),
    .X(_05777_));
 sky130_fd_sc_hd__mux2_1 _10865_ (.A0(_05776_),
    .A1(_05777_),
    .S(net1476),
    .X(_05778_));
 sky130_fd_sc_hd__nor2_1 _10866_ (.A(net1860),
    .B(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(\core.registers[24][5] ),
    .A1(\core.registers[25][5] ),
    .S(net1426),
    .X(_05780_));
 sky130_fd_sc_hd__a221o_1 _10868_ (.A1(net1699),
    .A2(\core.registers[26][5] ),
    .B1(\core.registers[27][5] ),
    .B2(net1426),
    .C1(net1712),
    .X(_05781_));
 sky130_fd_sc_hd__o21ai_1 _10869_ (.A1(net1877),
    .A2(_05780_),
    .B1(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__a211o_1 _10870_ (.A1(net1860),
    .A2(_05782_),
    .B1(_05779_),
    .C1(net1866),
    .X(_05783_));
 sky130_fd_sc_hd__or2_1 _10871_ (.A(\core.registers[13][5] ),
    .B(net1376),
    .X(_05784_));
 sky130_fd_sc_hd__o21a_1 _10872_ (.A1(\core.registers[12][5] ),
    .A2(net1424),
    .B1(net1711),
    .X(_05785_));
 sky130_fd_sc_hd__a22o_1 _10873_ (.A1(net1701),
    .A2(\core.registers[14][5] ),
    .B1(\core.registers[15][5] ),
    .B2(net1424),
    .X(_05786_));
 sky130_fd_sc_hd__a221o_1 _10874_ (.A1(_05784_),
    .A2(_05785_),
    .B1(_05786_),
    .B2(net1877),
    .C1(net1860),
    .X(_05787_));
 sky130_fd_sc_hd__a221o_1 _10875_ (.A1(net1701),
    .A2(\core.registers[30][5] ),
    .B1(\core.registers[31][5] ),
    .B2(net1424),
    .C1(net1711),
    .X(_05788_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(\core.registers[28][5] ),
    .A1(\core.registers[29][5] ),
    .S(net1424),
    .X(_05789_));
 sky130_fd_sc_hd__o21a_1 _10877_ (.A1(net1877),
    .A2(_05789_),
    .B1(_05788_),
    .X(_05790_));
 sky130_fd_sc_hd__o211a_1 _10878_ (.A1(net1718),
    .A2(_05790_),
    .B1(_05787_),
    .C1(net1866),
    .X(_05791_));
 sky130_fd_sc_hd__nor2_1 _10879_ (.A(net1487),
    .B(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__o2bb2a_2 _10880_ (.A1_N(_05783_),
    .A2_N(_05792_),
    .B1(net1491),
    .B2(_05775_),
    .X(_05793_));
 sky130_fd_sc_hd__a22o_4 _10881_ (.A1(net1070),
    .A2(net1059),
    .B1(_05793_),
    .B2(net1066),
    .X(_05794_));
 sky130_fd_sc_hd__o21ba_4 _10882_ (.A1(net1288),
    .A2(_05794_),
    .B1_N(_05764_),
    .X(_05795_));
 sky130_fd_sc_hd__and2_4 _10883_ (.A(_05763_),
    .B(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__nor2_4 _10884_ (.A(_05763_),
    .B(_05795_),
    .Y(_05797_));
 sky130_fd_sc_hd__nor2_8 _10885_ (.A(_05796_),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__inv_2 _10886_ (.A(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__a22o_1 _10887_ (.A1(\core.pipe1_resultRegister[4] ),
    .A2(net1239),
    .B1(net1269),
    .B2(\core.pipe1_csrData[4] ),
    .X(_05800_));
 sky130_fd_sc_hd__a21o_1 _10888_ (.A1(net1807),
    .A2(_04946_),
    .B1(net1811),
    .X(_05801_));
 sky130_fd_sc_hd__o211ai_2 _10889_ (.A1(_04558_),
    .A2(_04954_),
    .B1(_05801_),
    .C1(_04941_),
    .Y(_05802_));
 sky130_fd_sc_hd__mux2_8 _10890_ (.A0(net151),
    .A1(net136),
    .S(net1805),
    .X(_05803_));
 sky130_fd_sc_hd__o32ai_4 _10891_ (.A1(net1675),
    .A2(net1655),
    .A3(_05803_),
    .B1(net1658),
    .B2(\coreWBInterface.readDataBuffered[4] ),
    .Y(_05804_));
 sky130_fd_sc_hd__nor2_1 _10892_ (.A(net1812),
    .B(_05804_),
    .Y(_05805_));
 sky130_fd_sc_hd__a211o_1 _10893_ (.A1(\core.pipe1_loadResult[4] ),
    .A2(net1813),
    .B1(_04572_),
    .C1(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__a31o_4 _10894_ (.A1(net1189),
    .A2(_05802_),
    .A3(_05806_),
    .B1(_05800_),
    .X(_05807_));
 sky130_fd_sc_hd__and3_1 _10895_ (.A(net1850),
    .B(\core.registers[5][4] ),
    .C(net1664),
    .X(_05808_));
 sky130_fd_sc_hd__a21o_1 _10896_ (.A1(\core.registers[4][4] ),
    .A2(net1500),
    .B1(net1580),
    .X(_05809_));
 sky130_fd_sc_hd__o31a_1 _10897_ (.A1(\core.registers[1][4] ),
    .A2(net1591),
    .A3(net1500),
    .B1(net1606),
    .X(_05810_));
 sky130_fd_sc_hd__o221a_1 _10898_ (.A1(\core.registers[0][4] ),
    .A2(net1339),
    .B1(_05808_),
    .B2(_05809_),
    .C1(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__o22a_1 _10899_ (.A1(net1728),
    .A2(\core.registers[7][4] ),
    .B1(net1541),
    .B2(\core.registers[6][4] ),
    .X(_05812_));
 sky130_fd_sc_hd__o31a_1 _10900_ (.A1(net1726),
    .A2(\core.registers[3][4] ),
    .A3(net1590),
    .B1(net1620),
    .X(_05813_));
 sky130_fd_sc_hd__o221a_1 _10901_ (.A1(\core.registers[2][4] ),
    .A2(net1340),
    .B1(_05812_),
    .B2(net1580),
    .C1(_05813_),
    .X(_05814_));
 sky130_fd_sc_hd__and3_1 _10902_ (.A(net1850),
    .B(\core.registers[21][4] ),
    .C(net1664),
    .X(_05815_));
 sky130_fd_sc_hd__a21o_1 _10903_ (.A1(\core.registers[20][4] ),
    .A2(net1499),
    .B1(net1580),
    .X(_05816_));
 sky130_fd_sc_hd__o31a_1 _10904_ (.A1(\core.registers[17][4] ),
    .A2(net1591),
    .A3(net1499),
    .B1(net1606),
    .X(_05817_));
 sky130_fd_sc_hd__o221a_1 _10905_ (.A1(\core.registers[16][4] ),
    .A2(net1339),
    .B1(_05815_),
    .B2(_05816_),
    .C1(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__o22a_1 _10906_ (.A1(net1728),
    .A2(\core.registers[23][4] ),
    .B1(net1544),
    .B2(\core.registers[22][4] ),
    .X(_05819_));
 sky130_fd_sc_hd__o31a_1 _10907_ (.A1(net1728),
    .A2(\core.registers[19][4] ),
    .A3(net1591),
    .B1(net1623),
    .X(_05820_));
 sky130_fd_sc_hd__o221a_1 _10908_ (.A1(\core.registers[18][4] ),
    .A2(net1339),
    .B1(_05819_),
    .B2(net1580),
    .C1(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__o31a_1 _10909_ (.A1(net1569),
    .A2(_05818_),
    .A3(_05821_),
    .B1(net1633),
    .X(_05822_));
 sky130_fd_sc_hd__o31a_1 _10910_ (.A1(net1573),
    .A2(_05811_),
    .A3(_05814_),
    .B1(_05822_),
    .X(_05823_));
 sky130_fd_sc_hd__or2_1 _10911_ (.A(\core.registers[28][4] ),
    .B(net1557),
    .X(_05824_));
 sky130_fd_sc_hd__o211a_1 _10912_ (.A1(\core.registers[29][4] ),
    .A2(net1501),
    .B1(_05824_),
    .C1(net1739),
    .X(_05825_));
 sky130_fd_sc_hd__a31o_1 _10913_ (.A1(net1846),
    .A2(net1732),
    .A3(\core.registers[30][4] ),
    .B1(net1751),
    .X(_05826_));
 sky130_fd_sc_hd__a311o_1 _10914_ (.A1(net1846),
    .A2(\core.registers[31][4] ),
    .A3(net1557),
    .B1(_05825_),
    .C1(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__or2_1 _10915_ (.A(\core.registers[13][4] ),
    .B(net1502),
    .X(_05828_));
 sky130_fd_sc_hd__o211a_1 _10916_ (.A1(\core.registers[12][4] ),
    .A2(net1549),
    .B1(_05828_),
    .C1(net1739),
    .X(_05829_));
 sky130_fd_sc_hd__a31o_1 _10917_ (.A1(net1846),
    .A2(net1728),
    .A3(\core.registers[14][4] ),
    .B1(net1827),
    .X(_05830_));
 sky130_fd_sc_hd__a311o_1 _10918_ (.A1(net1846),
    .A2(\core.registers[15][4] ),
    .A3(net1542),
    .B1(_05829_),
    .C1(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__a21o_1 _10919_ (.A1(_05827_),
    .A2(_05831_),
    .B1(net1747),
    .X(_05832_));
 sky130_fd_sc_hd__and3_1 _10920_ (.A(net1850),
    .B(\core.registers[9][4] ),
    .C(net1663),
    .X(_05833_));
 sky130_fd_sc_hd__a21o_1 _10921_ (.A1(\core.registers[8][4] ),
    .A2(net1498),
    .B1(net1621),
    .X(_05834_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(\core.registers[10][4] ),
    .A1(\core.registers[11][4] ),
    .S(net1542),
    .X(_05835_));
 sky130_fd_sc_hd__o221a_1 _10923_ (.A1(_05833_),
    .A2(_05834_),
    .B1(_05835_),
    .B2(net1606),
    .C1(net1751),
    .X(_05836_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(\core.registers[24][4] ),
    .A1(\core.registers[25][4] ),
    .S(net1544),
    .X(_05837_));
 sky130_fd_sc_hd__a221o_1 _10925_ (.A1(net1728),
    .A2(\core.registers[26][4] ),
    .B1(\core.registers[27][4] ),
    .B2(net1544),
    .C1(net1739),
    .X(_05838_));
 sky130_fd_sc_hd__o211a_1 _10926_ (.A1(net1846),
    .A2(_05837_),
    .B1(_05838_),
    .C1(net1827),
    .X(_05839_));
 sky130_fd_sc_hd__o311a_1 _10927_ (.A1(net1835),
    .A2(_05836_),
    .A3(_05839_),
    .B1(net1637),
    .C1(_05832_),
    .X(_05840_));
 sky130_fd_sc_hd__or3_4 _10928_ (.A(net1159),
    .B(_05823_),
    .C(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__o211ai_4 _10929_ (.A1(net1156),
    .A2(net1053),
    .B1(_05841_),
    .C1(net1266),
    .Y(_05842_));
 sky130_fd_sc_hd__nor2_1 _10930_ (.A(\core.pipe0_currentInstruction[11] ),
    .B(_04468_),
    .Y(_05843_));
 sky130_fd_sc_hd__a211o_2 _10931_ (.A1(_04468_),
    .A2(_05842_),
    .B1(_05843_),
    .C1(_04481_),
    .X(_05844_));
 sky130_fd_sc_hd__nand2_2 _10932_ (.A(net1829),
    .B(_04481_),
    .Y(_05845_));
 sky130_fd_sc_hd__a21oi_4 _10933_ (.A1(_05844_),
    .A2(_05845_),
    .B1(net1287),
    .Y(_05846_));
 sky130_fd_sc_hd__a21o_4 _10934_ (.A1(_05844_),
    .A2(_05845_),
    .B1(net1287),
    .X(_05847_));
 sky130_fd_sc_hd__nor2_1 _10935_ (.A(net476),
    .B(net1284),
    .Y(_05848_));
 sky130_fd_sc_hd__o22a_1 _10936_ (.A1(net1694),
    .A2(\core.registers[23][4] ),
    .B1(net1413),
    .B2(\core.registers[22][4] ),
    .X(_05849_));
 sky130_fd_sc_hd__or3_1 _10937_ (.A(net1694),
    .B(\core.registers[19][4] ),
    .C(net1453),
    .X(_05850_));
 sky130_fd_sc_hd__o221a_1 _10938_ (.A1(\core.registers[18][4] ),
    .A2(net1334),
    .B1(_05849_),
    .B2(net1438),
    .C1(_05850_),
    .X(_05851_));
 sky130_fd_sc_hd__mux4_1 _10939_ (.A0(\core.registers[16][4] ),
    .A1(\core.registers[17][4] ),
    .A2(\core.registers[20][4] ),
    .A3(\core.registers[21][4] ),
    .S0(net1413),
    .S1(net1453),
    .X(_05852_));
 sky130_fd_sc_hd__mux2_1 _10940_ (.A0(_05851_),
    .A1(_05852_),
    .S(net1473),
    .X(_05853_));
 sky130_fd_sc_hd__o22a_1 _10941_ (.A1(net1693),
    .A2(\core.registers[7][4] ),
    .B1(net1410),
    .B2(\core.registers[6][4] ),
    .X(_05854_));
 sky130_fd_sc_hd__or3_1 _10942_ (.A(net1689),
    .B(\core.registers[3][4] ),
    .C(net1451),
    .X(_05855_));
 sky130_fd_sc_hd__o221a_1 _10943_ (.A1(\core.registers[2][4] ),
    .A2(net1334),
    .B1(_05854_),
    .B2(net1438),
    .C1(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__mux4_1 _10944_ (.A0(\core.registers[0][4] ),
    .A1(\core.registers[1][4] ),
    .A2(\core.registers[4][4] ),
    .A3(\core.registers[5][4] ),
    .S0(net1414),
    .S1(net1452),
    .X(_05857_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(_05856_),
    .A1(_05857_),
    .S(net1473),
    .X(_05858_));
 sky130_fd_sc_hd__mux2_1 _10946_ (.A0(_05853_),
    .A1(_05858_),
    .S(net1462),
    .X(_05859_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(\core.registers[10][4] ),
    .A1(\core.registers[11][4] ),
    .S(net1410),
    .X(_05860_));
 sky130_fd_sc_hd__mux2_1 _10948_ (.A0(\core.registers[8][4] ),
    .A1(\core.registers[9][4] ),
    .S(net1410),
    .X(_05861_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(_05860_),
    .A1(_05861_),
    .S(net1473),
    .X(_05862_));
 sky130_fd_sc_hd__nor2_1 _10950_ (.A(net1856),
    .B(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(\core.registers[24][4] ),
    .A1(\core.registers[25][4] ),
    .S(net1413),
    .X(_05864_));
 sky130_fd_sc_hd__a221o_1 _10952_ (.A1(net1693),
    .A2(\core.registers[26][4] ),
    .B1(\core.registers[27][4] ),
    .B2(net1413),
    .C1(net1711),
    .X(_05865_));
 sky130_fd_sc_hd__o21ai_1 _10953_ (.A1(net1874),
    .A2(_05864_),
    .B1(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__a211o_1 _10954_ (.A1(net1856),
    .A2(_05866_),
    .B1(_05863_),
    .C1(net1866),
    .X(_05867_));
 sky130_fd_sc_hd__a221o_1 _10955_ (.A1(net1696),
    .A2(\core.registers[30][4] ),
    .B1(\core.registers[31][4] ),
    .B2(net1417),
    .C1(net1711),
    .X(_05868_));
 sky130_fd_sc_hd__mux2_1 _10956_ (.A0(\core.registers[28][4] ),
    .A1(\core.registers[29][4] ),
    .S(net1423),
    .X(_05869_));
 sky130_fd_sc_hd__o21a_1 _10957_ (.A1(net1874),
    .A2(_05869_),
    .B1(_05868_),
    .X(_05870_));
 sky130_fd_sc_hd__or2_1 _10958_ (.A(\core.registers[12][4] ),
    .B(net1417),
    .X(_05871_));
 sky130_fd_sc_hd__o21a_1 _10959_ (.A1(\core.registers[13][4] ),
    .A2(net1376),
    .B1(net1711),
    .X(_05872_));
 sky130_fd_sc_hd__a22o_1 _10960_ (.A1(net1693),
    .A2(\core.registers[14][4] ),
    .B1(\core.registers[15][4] ),
    .B2(net1410),
    .X(_05873_));
 sky130_fd_sc_hd__a221o_1 _10961_ (.A1(_05871_),
    .A2(_05872_),
    .B1(_05873_),
    .B2(net1874),
    .C1(net1857),
    .X(_05874_));
 sky130_fd_sc_hd__o211a_1 _10962_ (.A1(net1718),
    .A2(_05870_),
    .B1(_05874_),
    .C1(net1865),
    .X(_05875_));
 sky130_fd_sc_hd__nor2_1 _10963_ (.A(net1487),
    .B(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__o2bb2a_2 _10964_ (.A1_N(_05867_),
    .A2_N(_05876_),
    .B1(net1491),
    .B2(_05859_),
    .X(_05877_));
 sky130_fd_sc_hd__a22o_4 _10965_ (.A1(net1070),
    .A2(_05807_),
    .B1(_05877_),
    .B2(net1066),
    .X(_05878_));
 sky130_fd_sc_hd__o21bai_4 _10966_ (.A1(net1288),
    .A2(_05878_),
    .B1_N(_05848_),
    .Y(_05879_));
 sky130_fd_sc_hd__inv_2 _10967_ (.A(_05879_),
    .Y(_05880_));
 sky130_fd_sc_hd__nor2_1 _10968_ (.A(net947),
    .B(_05879_),
    .Y(_05881_));
 sky130_fd_sc_hd__nand2_2 _10969_ (.A(net947),
    .B(_05879_),
    .Y(_05882_));
 sky130_fd_sc_hd__nand2b_4 _10970_ (.A_N(_05881_),
    .B(_05882_),
    .Y(_05883_));
 sky130_fd_sc_hd__a22o_1 _10971_ (.A1(\core.pipe1_resultRegister[3] ),
    .A2(net1239),
    .B1(net1269),
    .B2(\core.pipe1_csrData[3] ),
    .X(_05884_));
 sky130_fd_sc_hd__a21o_1 _10972_ (.A1(net1807),
    .A2(_05290_),
    .B1(net1811),
    .X(_05885_));
 sky130_fd_sc_hd__o211ai_1 _10973_ (.A1(_04558_),
    .A2(_05295_),
    .B1(_05885_),
    .C1(_05286_),
    .Y(_05886_));
 sky130_fd_sc_hd__mux2_8 _10974_ (.A0(net140),
    .A1(net135),
    .S(net1805),
    .X(_05887_));
 sky130_fd_sc_hd__o32ai_4 _10975_ (.A1(net1676),
    .A2(net1656),
    .A3(_05887_),
    .B1(net1658),
    .B2(\coreWBInterface.readDataBuffered[3] ),
    .Y(_05888_));
 sky130_fd_sc_hd__nor2_1 _10976_ (.A(net1812),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__a211o_1 _10977_ (.A1(\core.pipe1_loadResult[3] ),
    .A2(net1812),
    .B1(_04572_),
    .C1(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__a31o_2 _10978_ (.A1(net1189),
    .A2(_05886_),
    .A3(_05890_),
    .B1(_05884_),
    .X(_05891_));
 sky130_fd_sc_hd__and3_1 _10979_ (.A(net1850),
    .B(\core.registers[9][3] ),
    .C(net1663),
    .X(_05892_));
 sky130_fd_sc_hd__a21o_1 _10980_ (.A1(\core.registers[8][3] ),
    .A2(net1502),
    .B1(net1621),
    .X(_05893_));
 sky130_fd_sc_hd__mux2_1 _10981_ (.A0(\core.registers[10][3] ),
    .A1(\core.registers[11][3] ),
    .S(net1541),
    .X(_05894_));
 sky130_fd_sc_hd__o221a_1 _10982_ (.A1(_05892_),
    .A2(_05893_),
    .B1(_05894_),
    .B2(net1605),
    .C1(net1750),
    .X(_05895_));
 sky130_fd_sc_hd__mux2_1 _10983_ (.A0(\core.registers[24][3] ),
    .A1(\core.registers[25][3] ),
    .S(net1542),
    .X(_05896_));
 sky130_fd_sc_hd__a221o_1 _10984_ (.A1(net1732),
    .A2(\core.registers[26][3] ),
    .B1(\core.registers[27][3] ),
    .B2(net1549),
    .C1(net1739),
    .X(_05897_));
 sky130_fd_sc_hd__o211a_1 _10985_ (.A1(net1846),
    .A2(_05896_),
    .B1(_05897_),
    .C1(net1827),
    .X(_05898_));
 sky130_fd_sc_hd__or2_1 _10986_ (.A(\core.registers[28][3] ),
    .B(net1541),
    .X(_05899_));
 sky130_fd_sc_hd__o211a_1 _10987_ (.A1(\core.registers[29][3] ),
    .A2(net1499),
    .B1(_05899_),
    .C1(net1741),
    .X(_05900_));
 sky130_fd_sc_hd__a31o_1 _10988_ (.A1(net1844),
    .A2(net1728),
    .A3(\core.registers[30][3] ),
    .B1(net1750),
    .X(_05901_));
 sky130_fd_sc_hd__a311o_1 _10989_ (.A1(net1844),
    .A2(\core.registers[31][3] ),
    .A3(net1541),
    .B1(_05900_),
    .C1(_05901_),
    .X(_05902_));
 sky130_fd_sc_hd__or2_1 _10990_ (.A(\core.registers[13][3] ),
    .B(net1502),
    .X(_05903_));
 sky130_fd_sc_hd__o211a_1 _10991_ (.A1(\core.registers[12][3] ),
    .A2(net1539),
    .B1(_05903_),
    .C1(net1739),
    .X(_05904_));
 sky130_fd_sc_hd__a31o_1 _10992_ (.A1(net1844),
    .A2(net1729),
    .A3(\core.registers[14][3] ),
    .B1(net1827),
    .X(_05905_));
 sky130_fd_sc_hd__a311o_1 _10993_ (.A1(net1844),
    .A2(\core.registers[15][3] ),
    .A3(net1542),
    .B1(_05904_),
    .C1(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__a21o_1 _10994_ (.A1(_05902_),
    .A2(_05906_),
    .B1(net1746),
    .X(_05907_));
 sky130_fd_sc_hd__o311a_1 _10995_ (.A1(net1834),
    .A2(_05895_),
    .A3(_05898_),
    .B1(_05907_),
    .C1(net1637),
    .X(_05908_));
 sky130_fd_sc_hd__and3_1 _10996_ (.A(net1850),
    .B(\core.registers[5][3] ),
    .C(net1664),
    .X(_05909_));
 sky130_fd_sc_hd__a21o_1 _10997_ (.A1(\core.registers[4][3] ),
    .A2(net1499),
    .B1(net1580),
    .X(_05910_));
 sky130_fd_sc_hd__o31a_1 _10998_ (.A1(\core.registers[1][3] ),
    .A2(net1591),
    .A3(net1499),
    .B1(net1606),
    .X(_05911_));
 sky130_fd_sc_hd__o221a_1 _10999_ (.A1(\core.registers[0][3] ),
    .A2(net1340),
    .B1(_05909_),
    .B2(_05910_),
    .C1(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__o22a_1 _11000_ (.A1(net1727),
    .A2(\core.registers[7][3] ),
    .B1(net1538),
    .B2(\core.registers[6][3] ),
    .X(_05913_));
 sky130_fd_sc_hd__o31a_1 _11001_ (.A1(net1728),
    .A2(\core.registers[3][3] ),
    .A3(net1595),
    .B1(net1622),
    .X(_05914_));
 sky130_fd_sc_hd__o221a_1 _11002_ (.A1(\core.registers[2][3] ),
    .A2(net1340),
    .B1(_05913_),
    .B2(net1584),
    .C1(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__and3_1 _11003_ (.A(net1850),
    .B(\core.registers[21][3] ),
    .C(net1664),
    .X(_05916_));
 sky130_fd_sc_hd__a21o_1 _11004_ (.A1(\core.registers[20][3] ),
    .A2(net1498),
    .B1(net1584),
    .X(_05917_));
 sky130_fd_sc_hd__o31a_1 _11005_ (.A1(\core.registers[17][3] ),
    .A2(net1595),
    .A3(net1499),
    .B1(net1605),
    .X(_05918_));
 sky130_fd_sc_hd__o221a_1 _11006_ (.A1(\core.registers[16][3] ),
    .A2(net1340),
    .B1(_05916_),
    .B2(_05917_),
    .C1(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__o22a_1 _11007_ (.A1(net1728),
    .A2(\core.registers[23][3] ),
    .B1(net1541),
    .B2(\core.registers[22][3] ),
    .X(_05920_));
 sky130_fd_sc_hd__o31a_1 _11008_ (.A1(net1728),
    .A2(\core.registers[19][3] ),
    .A3(net1595),
    .B1(net1621),
    .X(_05921_));
 sky130_fd_sc_hd__o221a_1 _11009_ (.A1(\core.registers[18][3] ),
    .A2(net1340),
    .B1(_05920_),
    .B2(net1584),
    .C1(_05921_),
    .X(_05922_));
 sky130_fd_sc_hd__o31a_1 _11010_ (.A1(net1569),
    .A2(_05919_),
    .A3(_05922_),
    .B1(net1633),
    .X(_05923_));
 sky130_fd_sc_hd__o31a_1 _11011_ (.A1(net1573),
    .A2(_05912_),
    .A3(_05915_),
    .B1(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__or3_2 _11012_ (.A(net1159),
    .B(_05908_),
    .C(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__o211a_1 _11013_ (.A1(net1155),
    .A2(net1052),
    .B1(_05925_),
    .C1(net1265),
    .X(_05926_));
 sky130_fd_sc_hd__o21ba_1 _11014_ (.A1(\core.pipe0_currentInstruction[10] ),
    .A2(_04468_),
    .B1_N(_04481_),
    .X(_05927_));
 sky130_fd_sc_hd__o21ai_1 _11015_ (.A1(net1275),
    .A2(_05926_),
    .B1(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _11016_ (.A(\core.pipe0_currentInstruction[23] ),
    .B(_04481_),
    .Y(_05929_));
 sky130_fd_sc_hd__a21o_1 _11017_ (.A1(_05928_),
    .A2(_05929_),
    .B1(net1287),
    .X(_05930_));
 sky130_fd_sc_hd__inv_2 _11018_ (.A(net946),
    .Y(_05931_));
 sky130_fd_sc_hd__nor2_1 _11019_ (.A(net475),
    .B(net1283),
    .Y(_05932_));
 sky130_fd_sc_hd__o22a_1 _11020_ (.A1(net1693),
    .A2(\core.registers[23][3] ),
    .B1(net1410),
    .B2(\core.registers[22][3] ),
    .X(_05933_));
 sky130_fd_sc_hd__or3_1 _11021_ (.A(net1693),
    .B(\core.registers[19][3] ),
    .C(net1453),
    .X(_05934_));
 sky130_fd_sc_hd__o221a_1 _11022_ (.A1(\core.registers[18][3] ),
    .A2(net1338),
    .B1(_05933_),
    .B2(net1438),
    .C1(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__mux4_1 _11023_ (.A0(\core.registers[16][3] ),
    .A1(\core.registers[17][3] ),
    .A2(\core.registers[20][3] ),
    .A3(\core.registers[21][3] ),
    .S0(net1406),
    .S1(net1451),
    .X(_05936_));
 sky130_fd_sc_hd__mux2_1 _11024_ (.A0(_05935_),
    .A1(_05936_),
    .S(net1473),
    .X(_05937_));
 sky130_fd_sc_hd__o22a_1 _11025_ (.A1(net1691),
    .A2(\core.registers[7][3] ),
    .B1(net1407),
    .B2(\core.registers[6][3] ),
    .X(_05938_));
 sky130_fd_sc_hd__or3_1 _11026_ (.A(net1691),
    .B(\core.registers[3][3] ),
    .C(net1452),
    .X(_05939_));
 sky130_fd_sc_hd__o221a_1 _11027_ (.A1(\core.registers[2][3] ),
    .A2(net1334),
    .B1(_05938_),
    .B2(net1438),
    .C1(_05939_),
    .X(_05940_));
 sky130_fd_sc_hd__mux4_1 _11028_ (.A0(\core.registers[0][3] ),
    .A1(\core.registers[1][3] ),
    .A2(\core.registers[4][3] ),
    .A3(\core.registers[5][3] ),
    .S0(net1410),
    .S1(net1453),
    .X(_05941_));
 sky130_fd_sc_hd__mux2_1 _11029_ (.A0(_05940_),
    .A1(_05941_),
    .S(net1473),
    .X(_05942_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(_05937_),
    .A1(_05942_),
    .S(net1462),
    .X(_05943_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(\core.registers[10][3] ),
    .A1(\core.registers[11][3] ),
    .S(net1411),
    .X(_05944_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(\core.registers[8][3] ),
    .A1(\core.registers[9][3] ),
    .S(net1411),
    .X(_05945_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(_05944_),
    .A1(_05945_),
    .S(net1473),
    .X(_05946_));
 sky130_fd_sc_hd__nor2_1 _11034_ (.A(net1857),
    .B(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(\core.registers[24][3] ),
    .A1(\core.registers[25][3] ),
    .S(net1410),
    .X(_05948_));
 sky130_fd_sc_hd__a221o_1 _11036_ (.A1(net1696),
    .A2(\core.registers[26][3] ),
    .B1(\core.registers[27][3] ),
    .B2(net1417),
    .C1(net1711),
    .X(_05949_));
 sky130_fd_sc_hd__o21ai_1 _11037_ (.A1(net1874),
    .A2(_05948_),
    .B1(_05949_),
    .Y(_05950_));
 sky130_fd_sc_hd__a211o_1 _11038_ (.A1(net1857),
    .A2(_05950_),
    .B1(_05947_),
    .C1(net1865),
    .X(_05951_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(\core.registers[28][3] ),
    .A1(\core.registers[29][3] ),
    .S(net1411),
    .X(_05952_));
 sky130_fd_sc_hd__a221o_1 _11040_ (.A1(net1693),
    .A2(\core.registers[30][3] ),
    .B1(\core.registers[31][3] ),
    .B2(net1411),
    .C1(net1710),
    .X(_05953_));
 sky130_fd_sc_hd__o21a_1 _11041_ (.A1(net1874),
    .A2(_05952_),
    .B1(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__or2_1 _11042_ (.A(\core.registers[12][3] ),
    .B(net1408),
    .X(_05955_));
 sky130_fd_sc_hd__o21a_1 _11043_ (.A1(\core.registers[13][3] ),
    .A2(net1376),
    .B1(net1710),
    .X(_05956_));
 sky130_fd_sc_hd__a22o_1 _11044_ (.A1(net1693),
    .A2(\core.registers[14][3] ),
    .B1(\core.registers[15][3] ),
    .B2(net1411),
    .X(_05957_));
 sky130_fd_sc_hd__a221o_1 _11045_ (.A1(_05955_),
    .A2(_05956_),
    .B1(_05957_),
    .B2(net1874),
    .C1(net1857),
    .X(_05958_));
 sky130_fd_sc_hd__o211a_1 _11046_ (.A1(net1717),
    .A2(_05954_),
    .B1(_05958_),
    .C1(net1865),
    .X(_05959_));
 sky130_fd_sc_hd__nor2_1 _11047_ (.A(net1487),
    .B(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__a2bb2o_4 _11048_ (.A1_N(net1491),
    .A2_N(_05943_),
    .B1(_05951_),
    .B2(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__a2bb2o_4 _11049_ (.A1_N(_04663_),
    .A2_N(_05961_),
    .B1(net1052),
    .B2(net1070),
    .X(_05962_));
 sky130_fd_sc_hd__o21bai_4 _11050_ (.A1(net1287),
    .A2(_05962_),
    .B1_N(_05932_),
    .Y(_05963_));
 sky130_fd_sc_hd__inv_2 _11051_ (.A(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__nor2_1 _11052_ (.A(net887),
    .B(_05963_),
    .Y(_05965_));
 sky130_fd_sc_hd__nor2_2 _11053_ (.A(net946),
    .B(_05963_),
    .Y(_05966_));
 sky130_fd_sc_hd__nand2_2 _11054_ (.A(net946),
    .B(_05963_),
    .Y(_05967_));
 sky130_fd_sc_hd__nand2b_4 _11055_ (.A_N(_05966_),
    .B(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__a22o_1 _11056_ (.A1(\core.pipe1_resultRegister[2] ),
    .A2(net1239),
    .B1(net1270),
    .B2(\core.pipe1_csrData[2] ),
    .X(_05969_));
 sky130_fd_sc_hd__a21o_1 _11057_ (.A1(net1806),
    .A2(_05378_),
    .B1(net1810),
    .X(_05970_));
 sky130_fd_sc_hd__o211ai_1 _11058_ (.A1(_04558_),
    .A2(_05383_),
    .B1(_05970_),
    .C1(_05374_),
    .Y(_05971_));
 sky130_fd_sc_hd__mux2_8 _11059_ (.A0(net129),
    .A1(net134),
    .S(net1805),
    .X(_05972_));
 sky130_fd_sc_hd__o32ai_4 _11060_ (.A1(net1676),
    .A2(net1655),
    .A3(_05972_),
    .B1(net1659),
    .B2(\coreWBInterface.readDataBuffered[2] ),
    .Y(_05973_));
 sky130_fd_sc_hd__nor2_1 _11061_ (.A(net1812),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__a211o_1 _11062_ (.A1(\core.pipe1_loadResult[2] ),
    .A2(net1812),
    .B1(_04572_),
    .C1(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__a31o_2 _11063_ (.A1(net1189),
    .A2(_05971_),
    .A3(_05975_),
    .B1(_05969_),
    .X(_05976_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(\core.registers[8][2] ),
    .A1(\core.registers[9][2] ),
    .S(net1553),
    .X(_05977_));
 sky130_fd_sc_hd__mux2_1 _11065_ (.A0(\core.registers[10][2] ),
    .A1(\core.registers[11][2] ),
    .S(net1553),
    .X(_05978_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(\core.registers[24][2] ),
    .A1(\core.registers[25][2] ),
    .S(net1549),
    .X(_05979_));
 sky130_fd_sc_hd__a221o_1 _11067_ (.A1(net1731),
    .A2(\core.registers[26][2] ),
    .B1(\core.registers[27][2] ),
    .B2(net1555),
    .C1(net1740),
    .X(_05980_));
 sky130_fd_sc_hd__or2_1 _11068_ (.A(\core.registers[29][2] ),
    .B(net1502),
    .X(_05981_));
 sky130_fd_sc_hd__o211a_1 _11069_ (.A1(\core.registers[28][2] ),
    .A2(net1550),
    .B1(_05981_),
    .C1(net1740),
    .X(_05982_));
 sky130_fd_sc_hd__a31o_1 _11070_ (.A1(net1847),
    .A2(net1732),
    .A3(\core.registers[30][2] ),
    .B1(net1751),
    .X(_05983_));
 sky130_fd_sc_hd__a31o_1 _11071_ (.A1(net1847),
    .A2(\core.registers[31][2] ),
    .A3(net1550),
    .B1(_05983_),
    .X(_05984_));
 sky130_fd_sc_hd__or2_1 _11072_ (.A(\core.registers[17][2] ),
    .B(net1502),
    .X(_05985_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(\core.registers[12][2] ),
    .A1(\core.registers[13][2] ),
    .S(net1550),
    .X(_05986_));
 sky130_fd_sc_hd__mux2_1 _11074_ (.A0(\core.registers[14][2] ),
    .A1(\core.registers[15][2] ),
    .S(net1550),
    .X(_05987_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(_05986_),
    .A1(_05987_),
    .S(net1626),
    .X(_05988_));
 sky130_fd_sc_hd__o221a_1 _11076_ (.A1(_05982_),
    .A2(_05984_),
    .B1(_05988_),
    .B2(net1826),
    .C1(net1835),
    .X(_05989_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(_05977_),
    .A1(_05978_),
    .S(net1624),
    .X(_05990_));
 sky130_fd_sc_hd__o21a_1 _11078_ (.A1(net1847),
    .A2(_05979_),
    .B1(_05980_),
    .X(_05991_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(_05990_),
    .A1(_05991_),
    .S(net1826),
    .X(_05992_));
 sky130_fd_sc_hd__a211o_1 _11080_ (.A1(net1747),
    .A2(_05992_),
    .B1(_05989_),
    .C1(net1634),
    .X(_05993_));
 sky130_fd_sc_hd__or2_1 _11081_ (.A(\core.registers[7][2] ),
    .B(net1502),
    .X(_05994_));
 sky130_fd_sc_hd__o211a_1 _11082_ (.A1(\core.registers[6][2] ),
    .A2(net1562),
    .B1(_05994_),
    .C1(net1628),
    .X(_05995_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(\core.registers[4][2] ),
    .A1(\core.registers[5][2] ),
    .S(net1562),
    .X(_05996_));
 sky130_fd_sc_hd__a211o_1 _11084_ (.A1(net1607),
    .A2(_05996_),
    .B1(_05995_),
    .C1(net1582),
    .X(_05997_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(\core.registers[0][2] ),
    .A1(\core.registers[1][2] ),
    .S(net1564),
    .X(_05998_));
 sky130_fd_sc_hd__mux2_1 _11086_ (.A0(\core.registers[2][2] ),
    .A1(\core.registers[3][2] ),
    .S(net1564),
    .X(_05999_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(_05998_),
    .A1(_05999_),
    .S(net1628),
    .X(_06000_));
 sky130_fd_sc_hd__o211a_2 _11088_ (.A1(net1592),
    .A2(_06000_),
    .B1(_05997_),
    .C1(net1570),
    .X(_06001_));
 sky130_fd_sc_hd__o211a_1 _11089_ (.A1(\core.registers[16][2] ),
    .A2(net1555),
    .B1(_05985_),
    .C1(net1610),
    .X(_06002_));
 sky130_fd_sc_hd__mux2_1 _11090_ (.A0(\core.registers[18][2] ),
    .A1(\core.registers[19][2] ),
    .S(net1555),
    .X(_06003_));
 sky130_fd_sc_hd__a211o_1 _11091_ (.A1(net1625),
    .A2(_06003_),
    .B1(_06002_),
    .C1(net1592),
    .X(_06004_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(\core.registers[22][2] ),
    .A1(\core.registers[23][2] ),
    .S(net1554),
    .X(_06005_));
 sky130_fd_sc_hd__mux2_1 _11093_ (.A0(\core.registers[20][2] ),
    .A1(\core.registers[21][2] ),
    .S(net1554),
    .X(_06006_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(_06005_),
    .A1(_06006_),
    .S(net1610),
    .X(_06007_));
 sky130_fd_sc_hd__o211a_1 _11095_ (.A1(net1581),
    .A2(_06007_),
    .B1(_06004_),
    .C1(net1574),
    .X(_06008_));
 sky130_fd_sc_hd__o31a_4 _11096_ (.A1(net1638),
    .A2(_06001_),
    .A3(_06008_),
    .B1(_05993_),
    .X(_06009_));
 sky130_fd_sc_hd__o21a_1 _11097_ (.A1(net1159),
    .A2(_06009_),
    .B1(net1265),
    .X(_06010_));
 sky130_fd_sc_hd__o21ai_4 _11098_ (.A1(net1155),
    .A2(net1047),
    .B1(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__nor2_1 _11099_ (.A(\core.pipe0_currentInstruction[9] ),
    .B(_04468_),
    .Y(_06012_));
 sky130_fd_sc_hd__a211o_1 _11100_ (.A1(_04468_),
    .A2(_06011_),
    .B1(_06012_),
    .C1(_04481_),
    .X(_06013_));
 sky130_fd_sc_hd__nand2_1 _11101_ (.A(net1836),
    .B(_04481_),
    .Y(_06014_));
 sky130_fd_sc_hd__a21o_1 _11102_ (.A1(_06013_),
    .A2(_06014_),
    .B1(net1287),
    .X(_06015_));
 sky130_fd_sc_hd__nor2_1 _11103_ (.A(net472),
    .B(net1283),
    .Y(_06016_));
 sky130_fd_sc_hd__o22a_1 _11104_ (.A1(net1697),
    .A2(\core.registers[23][2] ),
    .B1(net1421),
    .B2(\core.registers[22][2] ),
    .X(_06017_));
 sky130_fd_sc_hd__or3_1 _11105_ (.A(net1697),
    .B(\core.registers[19][2] ),
    .C(net1456),
    .X(_06018_));
 sky130_fd_sc_hd__o221a_1 _11106_ (.A1(\core.registers[18][2] ),
    .A2(net1335),
    .B1(_06017_),
    .B2(net1441),
    .C1(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__mux4_1 _11107_ (.A0(\core.registers[16][2] ),
    .A1(\core.registers[17][2] ),
    .A2(\core.registers[20][2] ),
    .A3(\core.registers[21][2] ),
    .S0(net1421),
    .S1(net1455),
    .X(_06020_));
 sky130_fd_sc_hd__mux2_1 _11108_ (.A0(_06019_),
    .A1(_06020_),
    .S(net1474),
    .X(_06021_));
 sky130_fd_sc_hd__o22a_1 _11109_ (.A1(net1700),
    .A2(\core.registers[7][2] ),
    .B1(net1429),
    .B2(\core.registers[6][2] ),
    .X(_06022_));
 sky130_fd_sc_hd__or3_1 _11110_ (.A(net1699),
    .B(\core.registers[3][2] ),
    .C(net1458),
    .X(_06023_));
 sky130_fd_sc_hd__o221a_1 _11111_ (.A1(\core.registers[2][2] ),
    .A2(net1336),
    .B1(_06022_),
    .B2(net1441),
    .C1(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__mux4_1 _11112_ (.A0(\core.registers[0][2] ),
    .A1(\core.registers[1][2] ),
    .A2(\core.registers[4][2] ),
    .A3(\core.registers[5][2] ),
    .S0(net1428),
    .S1(net1458),
    .X(_06025_));
 sky130_fd_sc_hd__mux2_2 _11113_ (.A0(_06024_),
    .A1(_06025_),
    .S(net1475),
    .X(_06026_));
 sky130_fd_sc_hd__mux2_2 _11114_ (.A0(_06021_),
    .A1(_06026_),
    .S(net1463),
    .X(_06027_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(\core.registers[10][2] ),
    .A1(\core.registers[11][2] ),
    .S(net1420),
    .X(_06028_));
 sky130_fd_sc_hd__mux2_1 _11116_ (.A0(\core.registers[8][2] ),
    .A1(\core.registers[9][2] ),
    .S(net1420),
    .X(_06029_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(_06028_),
    .A1(_06029_),
    .S(net1474),
    .X(_06030_));
 sky130_fd_sc_hd__nor2_1 _11118_ (.A(net1859),
    .B(_06030_),
    .Y(_06031_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(\core.registers[24][2] ),
    .A1(\core.registers[25][2] ),
    .S(net1418),
    .X(_06032_));
 sky130_fd_sc_hd__a221o_1 _11120_ (.A1(net1695),
    .A2(\core.registers[26][2] ),
    .B1(\core.registers[27][2] ),
    .B2(net1418),
    .C1(net1712),
    .X(_06033_));
 sky130_fd_sc_hd__o21ai_1 _11121_ (.A1(net1876),
    .A2(_06032_),
    .B1(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__a211o_1 _11122_ (.A1(net1859),
    .A2(_06034_),
    .B1(_06031_),
    .C1(net1865),
    .X(_06035_));
 sky130_fd_sc_hd__a221o_1 _11123_ (.A1(net1696),
    .A2(\core.registers[30][2] ),
    .B1(\core.registers[31][2] ),
    .B2(net1418),
    .C1(net1712),
    .X(_06036_));
 sky130_fd_sc_hd__mux2_1 _11124_ (.A0(\core.registers[28][2] ),
    .A1(\core.registers[29][2] ),
    .S(net1418),
    .X(_06037_));
 sky130_fd_sc_hd__o21a_1 _11125_ (.A1(net1876),
    .A2(_06037_),
    .B1(_06036_),
    .X(_06038_));
 sky130_fd_sc_hd__or2_1 _11126_ (.A(\core.registers[12][2] ),
    .B(net1418),
    .X(_06039_));
 sky130_fd_sc_hd__o21a_1 _11127_ (.A1(\core.registers[13][2] ),
    .A2(net1376),
    .B1(net1712),
    .X(_06040_));
 sky130_fd_sc_hd__a22o_1 _11128_ (.A1(net1696),
    .A2(\core.registers[14][2] ),
    .B1(\core.registers[15][2] ),
    .B2(net1418),
    .X(_06041_));
 sky130_fd_sc_hd__a221o_1 _11129_ (.A1(_06039_),
    .A2(_06040_),
    .B1(_06041_),
    .B2(net1876),
    .C1(net1859),
    .X(_06042_));
 sky130_fd_sc_hd__o211a_1 _11130_ (.A1(net1718),
    .A2(_06038_),
    .B1(_06042_),
    .C1(net1864),
    .X(_06043_));
 sky130_fd_sc_hd__nor2_1 _11131_ (.A(net1488),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__a2bb2o_4 _11132_ (.A1_N(net1491),
    .A2_N(_06027_),
    .B1(_06035_),
    .B2(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__o2bb2a_2 _11133_ (.A1_N(net1070),
    .A2_N(net1047),
    .B1(_06045_),
    .B2(_04663_),
    .X(_06046_));
 sky130_fd_sc_hd__a21o_2 _11134_ (.A1(net1283),
    .A2(_06046_),
    .B1(_06016_),
    .X(_06047_));
 sky130_fd_sc_hd__inv_2 _11135_ (.A(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__and2_1 _11136_ (.A(net943),
    .B(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__nor2_1 _11137_ (.A(net943),
    .B(_06047_),
    .Y(_06050_));
 sky130_fd_sc_hd__and2_1 _11138_ (.A(net942),
    .B(_06047_),
    .X(_06051_));
 sky130_fd_sc_hd__inv_2 _11139_ (.A(_06051_),
    .Y(_06052_));
 sky130_fd_sc_hd__or2_4 _11140_ (.A(_06050_),
    .B(_06051_),
    .X(_06053_));
 sky130_fd_sc_hd__mux2_8 _11141_ (.A0(net118),
    .A1(net133),
    .S(net1805),
    .X(_06054_));
 sky130_fd_sc_hd__o32ai_4 _11142_ (.A1(net1676),
    .A2(net1655),
    .A3(_06054_),
    .B1(_04561_),
    .B2(\coreWBInterface.readDataBuffered[1] ),
    .Y(_06055_));
 sky130_fd_sc_hd__a21oi_1 _11143_ (.A1(\core.pipe1_loadResult[1] ),
    .A2(net1814),
    .B1(\core.pipe1_resultRegister[0] ),
    .Y(_06056_));
 sky130_fd_sc_hd__o21a_1 _11144_ (.A1(net1814),
    .A2(_06055_),
    .B1(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__a21o_1 _11145_ (.A1(net1810),
    .A2(_05461_),
    .B1(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__a21oi_1 _11146_ (.A1(net1190),
    .A2(_06058_),
    .B1(net1239),
    .Y(_06059_));
 sky130_fd_sc_hd__a31oi_1 _11147_ (.A1(_04557_),
    .A2(net1233),
    .A3(_05470_),
    .B1(_05462_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_1 _11148_ (.A(\core.pipe1_csrData[1] ),
    .B(net1268),
    .Y(_06061_));
 sky130_fd_sc_hd__o211a_1 _11149_ (.A1(_04524_),
    .A2(_04555_),
    .B1(_06061_),
    .C1(_04499_),
    .X(_06062_));
 sky130_fd_sc_hd__and2_1 _11150_ (.A(net1806),
    .B(_05466_),
    .X(_06063_));
 sky130_fd_sc_hd__a31o_1 _11151_ (.A1(net1187),
    .A2(_06060_),
    .A3(_06063_),
    .B1(_06062_),
    .X(_06064_));
 sky130_fd_sc_hd__o2bb2a_1 _11152_ (.A1_N(_04508_),
    .A2_N(_06064_),
    .B1(_06059_),
    .B2(net1809),
    .X(_06065_));
 sky130_fd_sc_hd__o221a_1 _11153_ (.A1(net1730),
    .A2(\core.registers[19][1] ),
    .B1(net1545),
    .B2(\core.registers[18][1] ),
    .C1(net1583),
    .X(_06066_));
 sky130_fd_sc_hd__o221a_1 _11154_ (.A1(net1733),
    .A2(\core.registers[23][1] ),
    .B1(net1559),
    .B2(\core.registers[22][1] ),
    .C1(net1594),
    .X(_06067_));
 sky130_fd_sc_hd__or3_1 _11155_ (.A(net1609),
    .B(_06066_),
    .C(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__mux2_1 _11156_ (.A0(\core.registers[16][1] ),
    .A1(\core.registers[17][1] ),
    .S(net1557),
    .X(_06069_));
 sky130_fd_sc_hd__o221a_1 _11157_ (.A1(net1851),
    .A2(\core.registers[20][1] ),
    .B1(\core.registers[21][1] ),
    .B2(net1501),
    .C1(net1594),
    .X(_06070_));
 sky130_fd_sc_hd__a211o_1 _11158_ (.A1(net1583),
    .A2(_06069_),
    .B1(_06070_),
    .C1(net1629),
    .X(_06071_));
 sky130_fd_sc_hd__o221a_1 _11159_ (.A1(net1733),
    .A2(\core.registers[3][1] ),
    .B1(net1565),
    .B2(\core.registers[2][1] ),
    .C1(net1581),
    .X(_06072_));
 sky130_fd_sc_hd__o221a_1 _11160_ (.A1(net1733),
    .A2(\core.registers[7][1] ),
    .B1(net1564),
    .B2(\core.registers[6][1] ),
    .C1(net1593),
    .X(_06073_));
 sky130_fd_sc_hd__mux2_1 _11161_ (.A0(\core.registers[0][1] ),
    .A1(\core.registers[1][1] ),
    .S(net1564),
    .X(_06074_));
 sky130_fd_sc_hd__o221a_1 _11162_ (.A1(net1850),
    .A2(\core.registers[4][1] ),
    .B1(\core.registers[5][1] ),
    .B2(net1501),
    .C1(net1593),
    .X(_06075_));
 sky130_fd_sc_hd__a211o_1 _11163_ (.A1(net1581),
    .A2(_06074_),
    .B1(_06075_),
    .C1(net1628),
    .X(_06076_));
 sky130_fd_sc_hd__o311a_2 _11164_ (.A1(net1608),
    .A2(_06072_),
    .A3(_06073_),
    .B1(_06076_),
    .C1(net1569),
    .X(_06077_));
 sky130_fd_sc_hd__a31o_1 _11165_ (.A1(net1573),
    .A2(_06068_),
    .A3(_06071_),
    .B1(_06077_),
    .X(_06078_));
 sky130_fd_sc_hd__mux2_1 _11166_ (.A0(\core.registers[8][1] ),
    .A1(\core.registers[9][1] ),
    .S(net1557),
    .X(_06079_));
 sky130_fd_sc_hd__a221o_1 _11167_ (.A1(net1732),
    .A2(\core.registers[10][1] ),
    .B1(\core.registers[11][1] ),
    .B2(net1557),
    .C1(net1609),
    .X(_06080_));
 sky130_fd_sc_hd__o21a_1 _11168_ (.A1(net1629),
    .A2(_06079_),
    .B1(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__or2_1 _11169_ (.A(\core.registers[13][1] ),
    .B(net1499),
    .X(_06082_));
 sky130_fd_sc_hd__o21a_1 _11170_ (.A1(\core.registers[12][1] ),
    .A2(net1544),
    .B1(net1606),
    .X(_06083_));
 sky130_fd_sc_hd__a22o_1 _11171_ (.A1(net1729),
    .A2(\core.registers[14][1] ),
    .B1(\core.registers[15][1] ),
    .B2(net1544),
    .X(_06084_));
 sky130_fd_sc_hd__a221o_1 _11172_ (.A1(_06082_),
    .A2(_06083_),
    .B1(_06084_),
    .B2(net1623),
    .C1(net1746),
    .X(_06085_));
 sky130_fd_sc_hd__o21a_1 _11173_ (.A1(net1835),
    .A2(_06081_),
    .B1(_06085_),
    .X(_06086_));
 sky130_fd_sc_hd__mux2_1 _11174_ (.A0(\core.registers[24][1] ),
    .A1(\core.registers[25][1] ),
    .S(net1545),
    .X(_06087_));
 sky130_fd_sc_hd__a221o_1 _11175_ (.A1(net1730),
    .A2(\core.registers[26][1] ),
    .B1(\core.registers[27][1] ),
    .B2(net1545),
    .C1(net1742),
    .X(_06088_));
 sky130_fd_sc_hd__o211a_1 _11176_ (.A1(net1846),
    .A2(_06087_),
    .B1(_06088_),
    .C1(net1746),
    .X(_06089_));
 sky130_fd_sc_hd__a21o_1 _11177_ (.A1(\core.registers[28][1] ),
    .A2(net1499),
    .B1(net1848),
    .X(_06090_));
 sky130_fd_sc_hd__a21o_1 _11178_ (.A1(\core.registers[29][1] ),
    .A2(net1544),
    .B1(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__a221o_1 _11179_ (.A1(net1730),
    .A2(\core.registers[30][1] ),
    .B1(\core.registers[31][1] ),
    .B2(net1544),
    .C1(net1743),
    .X(_06092_));
 sky130_fd_sc_hd__a311o_1 _11180_ (.A1(net1836),
    .A2(_06091_),
    .A3(_06092_),
    .B1(_06089_),
    .C1(net1751),
    .X(_06093_));
 sky130_fd_sc_hd__o211a_1 _11181_ (.A1(net1829),
    .A2(_06086_),
    .B1(_06093_),
    .C1(net1638),
    .X(_06094_));
 sky130_fd_sc_hd__a211o_2 _11182_ (.A1(net1633),
    .A2(_06078_),
    .B1(_06094_),
    .C1(net1160),
    .X(_06095_));
 sky130_fd_sc_hd__o211ai_4 _11183_ (.A1(net1156),
    .A2(net1041),
    .B1(_06095_),
    .C1(net1266),
    .Y(_06096_));
 sky130_fd_sc_hd__nor2_1 _11184_ (.A(\core.pipe0_currentInstruction[8] ),
    .B(_04468_),
    .Y(_06097_));
 sky130_fd_sc_hd__a211o_1 _11185_ (.A1(_04468_),
    .A2(_06096_),
    .B1(_06097_),
    .C1(_04481_),
    .X(_06098_));
 sky130_fd_sc_hd__nand2_1 _11186_ (.A(net1848),
    .B(_04481_),
    .Y(_06099_));
 sky130_fd_sc_hd__a21o_1 _11187_ (.A1(_06098_),
    .A2(_06099_),
    .B1(net1287),
    .X(_06100_));
 sky130_fd_sc_hd__inv_2 _11188_ (.A(net937),
    .Y(_06101_));
 sky130_fd_sc_hd__nor2_2 _11189_ (.A(net461),
    .B(net1283),
    .Y(_06102_));
 sky130_fd_sc_hd__o22a_1 _11190_ (.A1(net1701),
    .A2(\core.registers[23][1] ),
    .B1(net1425),
    .B2(\core.registers[22][1] ),
    .X(_06103_));
 sky130_fd_sc_hd__or3_1 _11191_ (.A(net1703),
    .B(\core.registers[19][1] ),
    .C(net1454),
    .X(_06104_));
 sky130_fd_sc_hd__o221a_1 _11192_ (.A1(\core.registers[18][1] ),
    .A2(net1338),
    .B1(_06103_),
    .B2(net1439),
    .C1(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__mux4_1 _11193_ (.A0(\core.registers[16][1] ),
    .A1(\core.registers[17][1] ),
    .A2(\core.registers[20][1] ),
    .A3(\core.registers[21][1] ),
    .S0(net1423),
    .S1(net1459),
    .X(_06106_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(_06105_),
    .A1(_06106_),
    .S(net1475),
    .X(_06107_));
 sky130_fd_sc_hd__o22a_1 _11195_ (.A1(net1699),
    .A2(\core.registers[7][1] ),
    .B1(net1428),
    .B2(\core.registers[6][1] ),
    .X(_06108_));
 sky130_fd_sc_hd__or3_1 _11196_ (.A(net1699),
    .B(\core.registers[3][1] ),
    .C(net1457),
    .X(_06109_));
 sky130_fd_sc_hd__o221a_1 _11197_ (.A1(\core.registers[2][1] ),
    .A2(net1335),
    .B1(_06108_),
    .B2(net1440),
    .C1(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__mux4_1 _11198_ (.A0(\core.registers[0][1] ),
    .A1(\core.registers[1][1] ),
    .A2(\core.registers[4][1] ),
    .A3(\core.registers[5][1] ),
    .S0(net1428),
    .S1(net1458),
    .X(_06111_));
 sky130_fd_sc_hd__mux2_2 _11199_ (.A0(_06110_),
    .A1(_06111_),
    .S(net1476),
    .X(_06112_));
 sky130_fd_sc_hd__mux2_1 _11200_ (.A0(_06107_),
    .A1(_06112_),
    .S(net1462),
    .X(_06113_));
 sky130_fd_sc_hd__or2_2 _11201_ (.A(net1491),
    .B(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__mux2_1 _11202_ (.A0(\core.registers[14][1] ),
    .A1(\core.registers[15][1] ),
    .S(net1414),
    .X(_06115_));
 sky130_fd_sc_hd__mux2_1 _11203_ (.A0(\core.registers[12][1] ),
    .A1(\core.registers[13][1] ),
    .S(net1414),
    .X(_06116_));
 sky130_fd_sc_hd__mux2_1 _11204_ (.A0(_06115_),
    .A1(_06116_),
    .S(net1477),
    .X(_06117_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(\core.registers[28][1] ),
    .A1(\core.registers[29][1] ),
    .S(net1413),
    .X(_06118_));
 sky130_fd_sc_hd__a221o_1 _11206_ (.A1(net1694),
    .A2(\core.registers[30][1] ),
    .B1(\core.registers[31][1] ),
    .B2(net1413),
    .C1(net1708),
    .X(_06119_));
 sky130_fd_sc_hd__o21ai_1 _11207_ (.A1(net1872),
    .A2(_06118_),
    .B1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__nand2_1 _11208_ (.A(net1857),
    .B(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__o211a_1 _11209_ (.A1(net1857),
    .A2(_06117_),
    .B1(_06121_),
    .C1(net1865),
    .X(_06122_));
 sky130_fd_sc_hd__a22o_1 _11210_ (.A1(net1703),
    .A2(\core.registers[26][1] ),
    .B1(\core.registers[27][1] ),
    .B2(net1413),
    .X(_06123_));
 sky130_fd_sc_hd__mux2_1 _11211_ (.A0(\core.registers[24][1] ),
    .A1(\core.registers[25][1] ),
    .S(net1413),
    .X(_06124_));
 sky130_fd_sc_hd__mux2_1 _11212_ (.A0(_06123_),
    .A1(_06124_),
    .S(net1711),
    .X(_06125_));
 sky130_fd_sc_hd__or2_1 _11213_ (.A(\core.registers[9][1] ),
    .B(net1378),
    .X(_06126_));
 sky130_fd_sc_hd__o21a_1 _11214_ (.A1(\core.registers[8][1] ),
    .A2(net1423),
    .B1(net1711),
    .X(_06127_));
 sky130_fd_sc_hd__a22o_1 _11215_ (.A1(net1701),
    .A2(\core.registers[10][1] ),
    .B1(\core.registers[11][1] ),
    .B2(net1423),
    .X(_06128_));
 sky130_fd_sc_hd__a221o_1 _11216_ (.A1(_06126_),
    .A2(_06127_),
    .B1(_06128_),
    .B2(net1877),
    .C1(net1857),
    .X(_06129_));
 sky130_fd_sc_hd__o211a_1 _11217_ (.A1(net1717),
    .A2(_06125_),
    .B1(_06129_),
    .C1(net1715),
    .X(_06130_));
 sky130_fd_sc_hd__o31ai_4 _11218_ (.A1(net1487),
    .A2(_06122_),
    .A3(_06130_),
    .B1(_06114_),
    .Y(_06131_));
 sky130_fd_sc_hd__o2bb2a_4 _11219_ (.A1_N(net1071),
    .A2_N(net1041),
    .B1(_06131_),
    .B2(_04663_),
    .X(_06132_));
 sky130_fd_sc_hd__a21oi_4 _11220_ (.A1(net1283),
    .A2(_06132_),
    .B1(_06102_),
    .Y(_06133_));
 sky130_fd_sc_hd__and2b_2 _11221_ (.A_N(net937),
    .B(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__nor2_1 _11222_ (.A(_06101_),
    .B(_06133_),
    .Y(_06135_));
 sky130_fd_sc_hd__xnor2_4 _11223_ (.A(net938),
    .B(_06133_),
    .Y(_06136_));
 sky130_fd_sc_hd__or2_4 _11224_ (.A(_06134_),
    .B(_06135_),
    .X(_06137_));
 sky130_fd_sc_hd__nand2_1 _11225_ (.A(\core.pipe1_csrData[0] ),
    .B(net1268),
    .Y(_06138_));
 sky130_fd_sc_hd__o211a_1 _11226_ (.A1(_04524_),
    .A2(_04555_),
    .B1(_06138_),
    .C1(_04499_),
    .X(_06139_));
 sky130_fd_sc_hd__mux2_8 _11227_ (.A0(net123),
    .A1(net158),
    .S(net1805),
    .X(_06140_));
 sky130_fd_sc_hd__o32a_1 _11228_ (.A1(net1674),
    .A2(net1660),
    .A3(_06140_),
    .B1(net1658),
    .B2(\coreWBInterface.readDataBuffered[24] ),
    .X(_06141_));
 sky130_fd_sc_hd__mux2_4 _11229_ (.A0(\core.pipe1_loadResult[24] ),
    .A1(_06141_),
    .S(net1757),
    .X(_06142_));
 sky130_fd_sc_hd__nand2_1 _11230_ (.A(_04949_),
    .B(_06142_),
    .Y(_06143_));
 sky130_fd_sc_hd__mux2_8 _11231_ (.A0(net169),
    .A1(net141),
    .S(net1805),
    .X(_06144_));
 sky130_fd_sc_hd__o32a_1 _11232_ (.A1(net1676),
    .A2(net1654),
    .A3(_06144_),
    .B1(net1659),
    .B2(\coreWBInterface.readDataBuffered[8] ),
    .X(_06145_));
 sky130_fd_sc_hd__mux2_1 _11233_ (.A0(\core.pipe1_loadResult[8] ),
    .A1(_06145_),
    .S(net1759),
    .X(_06146_));
 sky130_fd_sc_hd__or3b_1 _11234_ (.A(net1806),
    .B(_04935_),
    .C_N(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__and2_1 _11235_ (.A(net1810),
    .B(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__nand3_1 _11236_ (.A(_04557_),
    .B(net1233),
    .C(_06142_),
    .Y(_06149_));
 sky130_fd_sc_hd__a31o_1 _11237_ (.A1(net1187),
    .A2(_06148_),
    .A3(_06149_),
    .B1(_06139_),
    .X(_06150_));
 sky130_fd_sc_hd__mux2_8 _11238_ (.A0(net107),
    .A1(net132),
    .S(\localMemoryInterface.lastRBankSelect ),
    .X(_06151_));
 sky130_fd_sc_hd__o32a_1 _11239_ (.A1(net1676),
    .A2(net1655),
    .A3(_06151_),
    .B1(net1659),
    .B2(\coreWBInterface.readDataBuffered[0] ),
    .X(_06152_));
 sky130_fd_sc_hd__mux2_1 _11240_ (.A0(\core.pipe1_loadResult[0] ),
    .A1(_06152_),
    .S(net1759),
    .X(_06153_));
 sky130_fd_sc_hd__mux2_8 _11241_ (.A0(net114),
    .A1(net149),
    .S(net1805),
    .X(_06154_));
 sky130_fd_sc_hd__o32a_1 _11242_ (.A1(net1673),
    .A2(net1651),
    .A3(_06154_),
    .B1(net1657),
    .B2(\coreWBInterface.readDataBuffered[16] ),
    .X(_06155_));
 sky130_fd_sc_hd__mux2_4 _11243_ (.A0(\core.pipe1_loadResult[16] ),
    .A1(_06155_),
    .S(net1758),
    .X(_06156_));
 sky130_fd_sc_hd__a31o_1 _11244_ (.A1(_04549_),
    .A2(_04558_),
    .A3(_06156_),
    .B1(_04401_),
    .X(_06157_));
 sky130_fd_sc_hd__o21ai_1 _11245_ (.A1(net1809),
    .A2(_06153_),
    .B1(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__a21oi_1 _11246_ (.A1(net1187),
    .A2(_06158_),
    .B1(net1239),
    .Y(_06159_));
 sky130_fd_sc_hd__o2bb2a_2 _11247_ (.A1_N(_04508_),
    .A2_N(_06150_),
    .B1(_06159_),
    .B2(net1810),
    .X(_06160_));
 sky130_fd_sc_hd__mux2_1 _11248_ (.A0(\core.registers[14][0] ),
    .A1(\core.registers[15][0] ),
    .S(net1535),
    .X(_06161_));
 sky130_fd_sc_hd__mux2_1 _11249_ (.A0(\core.registers[12][0] ),
    .A1(\core.registers[13][0] ),
    .S(net1540),
    .X(_06162_));
 sky130_fd_sc_hd__mux2_1 _11250_ (.A0(_06161_),
    .A1(_06162_),
    .S(net1605),
    .X(_06163_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(\core.registers[28][0] ),
    .A1(\core.registers[29][0] ),
    .S(net1540),
    .X(_06164_));
 sky130_fd_sc_hd__a221o_1 _11252_ (.A1(net1729),
    .A2(\core.registers[30][0] ),
    .B1(\core.registers[31][0] ),
    .B2(net1540),
    .C1(net1743),
    .X(_06165_));
 sky130_fd_sc_hd__o21a_1 _11253_ (.A1(net1848),
    .A2(_06164_),
    .B1(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__mux2_1 _11254_ (.A0(\core.registers[8][0] ),
    .A1(\core.registers[9][0] ),
    .S(net1535),
    .X(_06167_));
 sky130_fd_sc_hd__mux2_1 _11255_ (.A0(\core.registers[10][0] ),
    .A1(\core.registers[11][0] ),
    .S(net1535),
    .X(_06168_));
 sky130_fd_sc_hd__mux2_1 _11256_ (.A0(_06167_),
    .A1(_06168_),
    .S(net1620),
    .X(_06169_));
 sky130_fd_sc_hd__mux2_1 _11257_ (.A0(\core.registers[24][0] ),
    .A1(\core.registers[25][0] ),
    .S(net1540),
    .X(_06170_));
 sky130_fd_sc_hd__a22o_1 _11258_ (.A1(net1729),
    .A2(\core.registers[26][0] ),
    .B1(\core.registers[27][0] ),
    .B2(net1540),
    .X(_06171_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(_06170_),
    .A1(_06171_),
    .S(net1848),
    .X(_06172_));
 sky130_fd_sc_hd__mux4_2 _11260_ (.A0(_06163_),
    .A1(_06166_),
    .A2(_06169_),
    .A3(_06172_),
    .S0(net1829),
    .S1(net1746),
    .X(_06173_));
 sky130_fd_sc_hd__and3_1 _11261_ (.A(net1850),
    .B(\core.registers[5][0] ),
    .C(net1664),
    .X(_06174_));
 sky130_fd_sc_hd__a211o_1 _11262_ (.A1(\core.registers[4][0] ),
    .A2(net1498),
    .B1(_06174_),
    .C1(net1579),
    .X(_06175_));
 sky130_fd_sc_hd__o31a_1 _11263_ (.A1(\core.registers[1][0] ),
    .A2(net1590),
    .A3(net1498),
    .B1(net1605),
    .X(_06176_));
 sky130_fd_sc_hd__o211a_1 _11264_ (.A1(\core.registers[0][0] ),
    .A2(net1339),
    .B1(_06175_),
    .C1(_06176_),
    .X(_06177_));
 sky130_fd_sc_hd__o22a_1 _11265_ (.A1(net1726),
    .A2(\core.registers[7][0] ),
    .B1(net1537),
    .B2(\core.registers[6][0] ),
    .X(_06178_));
 sky130_fd_sc_hd__o31a_1 _11266_ (.A1(net1726),
    .A2(\core.registers[3][0] ),
    .A3(net1590),
    .B1(net1620),
    .X(_06179_));
 sky130_fd_sc_hd__o221a_1 _11267_ (.A1(\core.registers[2][0] ),
    .A2(net1339),
    .B1(_06178_),
    .B2(net1579),
    .C1(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__and3_1 _11268_ (.A(net1850),
    .B(\core.registers[21][0] ),
    .C(net1662),
    .X(_06181_));
 sky130_fd_sc_hd__a21o_1 _11269_ (.A1(\core.registers[20][0] ),
    .A2(net1498),
    .B1(net1580),
    .X(_06182_));
 sky130_fd_sc_hd__o31a_1 _11270_ (.A1(\core.registers[17][0] ),
    .A2(net1590),
    .A3(net1498),
    .B1(net1605),
    .X(_06183_));
 sky130_fd_sc_hd__o221a_1 _11271_ (.A1(\core.registers[16][0] ),
    .A2(net1339),
    .B1(_06181_),
    .B2(_06182_),
    .C1(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__o22a_1 _11272_ (.A1(net1727),
    .A2(\core.registers[23][0] ),
    .B1(net1537),
    .B2(\core.registers[22][0] ),
    .X(_06185_));
 sky130_fd_sc_hd__o31a_1 _11273_ (.A1(net1727),
    .A2(\core.registers[19][0] ),
    .A3(net1591),
    .B1(net1622),
    .X(_06186_));
 sky130_fd_sc_hd__o221a_1 _11274_ (.A1(\core.registers[18][0] ),
    .A2(net1339),
    .B1(_06185_),
    .B2(net1579),
    .C1(_06186_),
    .X(_06187_));
 sky130_fd_sc_hd__or3_1 _11275_ (.A(net1569),
    .B(_06184_),
    .C(_06187_),
    .X(_06188_));
 sky130_fd_sc_hd__o311a_1 _11276_ (.A1(net1573),
    .A2(_06177_),
    .A3(_06180_),
    .B1(_06188_),
    .C1(net1633),
    .X(_06189_));
 sky130_fd_sc_hd__a211o_1 _11277_ (.A1(net1637),
    .A2(_06173_),
    .B1(_06189_),
    .C1(net1159),
    .X(_06190_));
 sky130_fd_sc_hd__o211a_1 _11278_ (.A1(net1156),
    .A2(net1038),
    .B1(_06190_),
    .C1(net1266),
    .X(_06191_));
 sky130_fd_sc_hd__o21ba_1 _11279_ (.A1(\core.pipe0_currentInstruction[7] ),
    .A2(_04468_),
    .B1_N(_04481_),
    .X(_06192_));
 sky130_fd_sc_hd__o21ai_2 _11280_ (.A1(net1275),
    .A2(_06191_),
    .B1(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__nand2_1 _11281_ (.A(net1852),
    .B(_04481_),
    .Y(_06194_));
 sky130_fd_sc_hd__a21oi_1 _11282_ (.A1(_06193_),
    .A2(_06194_),
    .B1(net1287),
    .Y(_06195_));
 sky130_fd_sc_hd__a21o_4 _11283_ (.A1(_06193_),
    .A2(_06194_),
    .B1(net1287),
    .X(_06196_));
 sky130_fd_sc_hd__o22a_1 _11284_ (.A1(net1691),
    .A2(\core.registers[23][0] ),
    .B1(net1406),
    .B2(\core.registers[22][0] ),
    .X(_06197_));
 sky130_fd_sc_hd__or3_1 _11285_ (.A(net1689),
    .B(\core.registers[19][0] ),
    .C(net1451),
    .X(_06198_));
 sky130_fd_sc_hd__o221a_1 _11286_ (.A1(\core.registers[18][0] ),
    .A2(net1334),
    .B1(_06197_),
    .B2(net1438),
    .C1(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__mux4_1 _11287_ (.A0(\core.registers[16][0] ),
    .A1(\core.registers[17][0] ),
    .A2(\core.registers[20][0] ),
    .A3(\core.registers[21][0] ),
    .S0(net1406),
    .S1(net1451),
    .X(_06200_));
 sky130_fd_sc_hd__mux2_1 _11288_ (.A0(_06199_),
    .A1(_06200_),
    .S(net1472),
    .X(_06201_));
 sky130_fd_sc_hd__o22a_1 _11289_ (.A1(net1691),
    .A2(\core.registers[7][0] ),
    .B1(net1406),
    .B2(\core.registers[6][0] ),
    .X(_06202_));
 sky130_fd_sc_hd__or3_1 _11290_ (.A(net1689),
    .B(\core.registers[3][0] ),
    .C(net1451),
    .X(_06203_));
 sky130_fd_sc_hd__o221a_1 _11291_ (.A1(\core.registers[2][0] ),
    .A2(net1334),
    .B1(_06202_),
    .B2(net1438),
    .C1(_06203_),
    .X(_06204_));
 sky130_fd_sc_hd__mux4_1 _11292_ (.A0(\core.registers[0][0] ),
    .A1(\core.registers[1][0] ),
    .A2(\core.registers[4][0] ),
    .A3(\core.registers[5][0] ),
    .S0(net1406),
    .S1(net1452),
    .X(_06205_));
 sky130_fd_sc_hd__mux2_1 _11293_ (.A0(_06204_),
    .A1(_06205_),
    .S(net1472),
    .X(_06206_));
 sky130_fd_sc_hd__mux2_1 _11294_ (.A0(_06201_),
    .A1(_06206_),
    .S(net1462),
    .X(_06207_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(\core.registers[14][0] ),
    .A1(\core.registers[15][0] ),
    .S(net1404),
    .X(_06208_));
 sky130_fd_sc_hd__mux2_1 _11296_ (.A0(\core.registers[12][0] ),
    .A1(\core.registers[13][0] ),
    .S(net1409),
    .X(_06209_));
 sky130_fd_sc_hd__mux2_1 _11297_ (.A0(_06208_),
    .A1(_06209_),
    .S(net1472),
    .X(_06210_));
 sky130_fd_sc_hd__mux2_1 _11298_ (.A0(\core.registers[28][0] ),
    .A1(\core.registers[29][0] ),
    .S(net1409),
    .X(_06211_));
 sky130_fd_sc_hd__a221o_1 _11299_ (.A1(net1692),
    .A2(\core.registers[30][0] ),
    .B1(\core.registers[31][0] ),
    .B2(net1409),
    .C1(net1707),
    .X(_06212_));
 sky130_fd_sc_hd__o21a_1 _11300_ (.A1(net1872),
    .A2(_06211_),
    .B1(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__mux2_1 _11301_ (.A0(_06210_),
    .A1(_06213_),
    .S(net1856),
    .X(_06214_));
 sky130_fd_sc_hd__a22o_1 _11302_ (.A1(net1692),
    .A2(\core.registers[26][0] ),
    .B1(\core.registers[27][0] ),
    .B2(net1409),
    .X(_06215_));
 sky130_fd_sc_hd__mux2_1 _11303_ (.A0(\core.registers[24][0] ),
    .A1(\core.registers[25][0] ),
    .S(net1409),
    .X(_06216_));
 sky130_fd_sc_hd__mux2_1 _11304_ (.A0(_06215_),
    .A1(_06216_),
    .S(net1707),
    .X(_06217_));
 sky130_fd_sc_hd__or2_1 _11305_ (.A(\core.registers[9][0] ),
    .B(net1377),
    .X(_06218_));
 sky130_fd_sc_hd__o21a_1 _11306_ (.A1(\core.registers[8][0] ),
    .A2(net1404),
    .B1(net1707),
    .X(_06219_));
 sky130_fd_sc_hd__a22o_1 _11307_ (.A1(net1690),
    .A2(\core.registers[10][0] ),
    .B1(\core.registers[11][0] ),
    .B2(net1404),
    .X(_06220_));
 sky130_fd_sc_hd__a221o_1 _11308_ (.A1(_06218_),
    .A2(_06219_),
    .B1(_06220_),
    .B2(net1872),
    .C1(net1856),
    .X(_06221_));
 sky130_fd_sc_hd__o211a_1 _11309_ (.A1(net1718),
    .A2(_06217_),
    .B1(_06221_),
    .C1(net1715),
    .X(_06222_));
 sky130_fd_sc_hd__a211o_2 _11310_ (.A1(net1866),
    .A2(_06214_),
    .B1(_06222_),
    .C1(net1488),
    .X(_06223_));
 sky130_fd_sc_hd__o21ai_2 _11311_ (.A1(net1492),
    .A2(_06207_),
    .B1(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__o2bb2a_2 _11312_ (.A1_N(net1071),
    .A2_N(net1038),
    .B1(_06224_),
    .B2(_04663_),
    .X(_06225_));
 sky130_fd_sc_hd__nand2_1 _11313_ (.A(net450),
    .B(net1287),
    .Y(_06226_));
 sky130_fd_sc_hd__o21ai_4 _11314_ (.A1(net1287),
    .A2(_06225_),
    .B1(_06226_),
    .Y(_06227_));
 sky130_fd_sc_hd__nor2_1 _11315_ (.A(net931),
    .B(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__a2bb2o_4 _11316_ (.A1_N(_06136_),
    .A2_N(_06228_),
    .B1(net938),
    .B2(_06133_),
    .X(_06229_));
 sky130_fd_sc_hd__a21o_1 _11317_ (.A1(_06053_),
    .A2(_06229_),
    .B1(_06049_),
    .X(_06230_));
 sky130_fd_sc_hd__a21o_2 _11318_ (.A1(_05968_),
    .A2(_06230_),
    .B1(_05965_),
    .X(_06231_));
 sky130_fd_sc_hd__and3_1 _11319_ (.A(_05799_),
    .B(_05883_),
    .C(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__nand2_1 _11320_ (.A(net947),
    .B(_05880_),
    .Y(_06233_));
 sky130_fd_sc_hd__or2_1 _11321_ (.A(_05798_),
    .B(_06233_),
    .X(_06234_));
 sky130_fd_sc_hd__nand2b_1 _11322_ (.A_N(_05763_),
    .B(_05795_),
    .Y(_06235_));
 sky130_fd_sc_hd__nand2_2 _11323_ (.A(_06234_),
    .B(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__o31a_1 _11324_ (.A1(_05717_),
    .A2(_06232_),
    .A3(_06236_),
    .B1(_05718_),
    .X(_06237_));
 sky130_fd_sc_hd__a221o_1 _11325_ (.A1(\core.pipe1_resultRegister[8] ),
    .A2(_04498_),
    .B1(net1268),
    .B2(\core.pipe1_csrData[8] ),
    .C1(_04599_),
    .X(_06238_));
 sky130_fd_sc_hd__and3_1 _11326_ (.A(_04571_),
    .B(_04936_),
    .C(_06147_),
    .X(_06239_));
 sky130_fd_sc_hd__a21boi_1 _11327_ (.A1(_04944_),
    .A2(_06156_),
    .B1_N(_04945_),
    .Y(_06240_));
 sky130_fd_sc_hd__a21o_1 _11328_ (.A1(_04950_),
    .A2(_06143_),
    .B1(_04582_),
    .X(_06241_));
 sky130_fd_sc_hd__o211a_1 _11329_ (.A1(_04551_),
    .A2(_06240_),
    .B1(_06241_),
    .C1(_04948_),
    .X(_06242_));
 sky130_fd_sc_hd__o21ai_1 _11330_ (.A1(_06239_),
    .A2(_06242_),
    .B1(net1189),
    .Y(_06243_));
 sky130_fd_sc_hd__a22o_1 _11331_ (.A1(\core.pipe1_resultRegister[8] ),
    .A2(_04507_),
    .B1(_06238_),
    .B2(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(\core.registers[8][8] ),
    .A1(\core.registers[9][8] ),
    .S(net1549),
    .X(_06245_));
 sky130_fd_sc_hd__mux2_1 _11333_ (.A0(\core.registers[10][8] ),
    .A1(\core.registers[11][8] ),
    .S(net1547),
    .X(_06246_));
 sky130_fd_sc_hd__mux2_1 _11334_ (.A0(_06245_),
    .A1(_06246_),
    .S(net1626),
    .X(_06247_));
 sky130_fd_sc_hd__mux2_1 _11335_ (.A0(\core.registers[24][8] ),
    .A1(\core.registers[25][8] ),
    .S(net1549),
    .X(_06248_));
 sky130_fd_sc_hd__and3_1 _11336_ (.A(net1844),
    .B(\core.registers[27][8] ),
    .C(net1549),
    .X(_06249_));
 sky130_fd_sc_hd__a211o_1 _11337_ (.A1(\core.registers[26][8] ),
    .A2(_04608_),
    .B1(_06249_),
    .C1(net1750),
    .X(_06250_));
 sky130_fd_sc_hd__a21o_1 _11338_ (.A1(net1739),
    .A2(_06248_),
    .B1(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__mux2_1 _11339_ (.A0(\core.registers[28][8] ),
    .A1(\core.registers[29][8] ),
    .S(net1549),
    .X(_06252_));
 sky130_fd_sc_hd__a221o_1 _11340_ (.A1(net1732),
    .A2(\core.registers[30][8] ),
    .B1(\core.registers[31][8] ),
    .B2(net1549),
    .C1(net1741),
    .X(_06253_));
 sky130_fd_sc_hd__mux2_1 _11341_ (.A0(\core.registers[12][8] ),
    .A1(\core.registers[13][8] ),
    .S(net1549),
    .X(_06254_));
 sky130_fd_sc_hd__mux2_1 _11342_ (.A0(\core.registers[14][8] ),
    .A1(\core.registers[15][8] ),
    .S(net1549),
    .X(_06255_));
 sky130_fd_sc_hd__mux2_1 _11343_ (.A0(_06254_),
    .A1(_06255_),
    .S(net1626),
    .X(_06256_));
 sky130_fd_sc_hd__o21a_1 _11344_ (.A1(net1845),
    .A2(_06252_),
    .B1(_06253_),
    .X(_06257_));
 sky130_fd_sc_hd__mux2_1 _11345_ (.A0(_06256_),
    .A1(_06257_),
    .S(net1827),
    .X(_06258_));
 sky130_fd_sc_hd__o211a_1 _11346_ (.A1(net1827),
    .A2(_06247_),
    .B1(_06251_),
    .C1(net1747),
    .X(_06259_));
 sky130_fd_sc_hd__a211o_1 _11347_ (.A1(net1834),
    .A2(_06258_),
    .B1(_06259_),
    .C1(net1633),
    .X(_06260_));
 sky130_fd_sc_hd__or2_1 _11348_ (.A(\core.registers[22][8] ),
    .B(net1558),
    .X(_06261_));
 sky130_fd_sc_hd__or2_1 _11349_ (.A(\core.registers[1][8] ),
    .B(net1501),
    .X(_06262_));
 sky130_fd_sc_hd__or2_1 _11350_ (.A(\core.registers[6][8] ),
    .B(net1558),
    .X(_06263_));
 sky130_fd_sc_hd__o211a_1 _11351_ (.A1(net1733),
    .A2(\core.registers[7][8] ),
    .B1(net1629),
    .C1(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__mux2_1 _11352_ (.A0(\core.registers[4][8] ),
    .A1(\core.registers[5][8] ),
    .S(net1559),
    .X(_06265_));
 sky130_fd_sc_hd__a211o_1 _11353_ (.A1(net1609),
    .A2(_06265_),
    .B1(_06264_),
    .C1(net1583),
    .X(_06266_));
 sky130_fd_sc_hd__o211a_1 _11354_ (.A1(\core.registers[0][8] ),
    .A2(net1559),
    .B1(_06262_),
    .C1(net1609),
    .X(_06267_));
 sky130_fd_sc_hd__mux2_1 _11355_ (.A0(\core.registers[2][8] ),
    .A1(\core.registers[3][8] ),
    .S(net1559),
    .X(_06268_));
 sky130_fd_sc_hd__a211o_1 _11356_ (.A1(net1629),
    .A2(_06268_),
    .B1(_06267_),
    .C1(net1594),
    .X(_06269_));
 sky130_fd_sc_hd__mux2_1 _11357_ (.A0(\core.registers[16][8] ),
    .A1(\core.registers[17][8] ),
    .S(net1558),
    .X(_06270_));
 sky130_fd_sc_hd__mux2_1 _11358_ (.A0(\core.registers[18][8] ),
    .A1(\core.registers[19][8] ),
    .S(net1559),
    .X(_06271_));
 sky130_fd_sc_hd__mux2_1 _11359_ (.A0(_06270_),
    .A1(_06271_),
    .S(net1629),
    .X(_06272_));
 sky130_fd_sc_hd__o211a_1 _11360_ (.A1(net1733),
    .A2(\core.registers[23][8] ),
    .B1(net1629),
    .C1(_06261_),
    .X(_06273_));
 sky130_fd_sc_hd__mux2_1 _11361_ (.A0(\core.registers[20][8] ),
    .A1(\core.registers[21][8] ),
    .S(net1558),
    .X(_06274_));
 sky130_fd_sc_hd__a211o_1 _11362_ (.A1(net1609),
    .A2(_06274_),
    .B1(_06273_),
    .C1(net1582),
    .X(_06275_));
 sky130_fd_sc_hd__o211a_1 _11363_ (.A1(net1594),
    .A2(_06272_),
    .B1(_06275_),
    .C1(net1574),
    .X(_06276_));
 sky130_fd_sc_hd__a311o_1 _11364_ (.A1(net1570),
    .A2(_06266_),
    .A3(_06269_),
    .B1(_06276_),
    .C1(net1638),
    .X(_06277_));
 sky130_fd_sc_hd__a21o_2 _11365_ (.A1(_06260_),
    .A2(_06277_),
    .B1(net1160),
    .X(_06278_));
 sky130_fd_sc_hd__o211a_4 _11366_ (.A1(net1155),
    .A2(net961),
    .B1(_06278_),
    .C1(net1265),
    .X(_06279_));
 sky130_fd_sc_hd__or2_1 _11367_ (.A(net1819),
    .B(_04484_),
    .X(_06280_));
 sky130_fd_sc_hd__o211a_1 _11368_ (.A1(net1194),
    .A2(_06279_),
    .B1(_06280_),
    .C1(net1282),
    .X(_06281_));
 sky130_fd_sc_hd__mux2_1 _11369_ (.A0(\core.registers[28][8] ),
    .A1(\core.registers[29][8] ),
    .S(net1417),
    .X(_06282_));
 sky130_fd_sc_hd__a221o_1 _11370_ (.A1(net1696),
    .A2(\core.registers[30][8] ),
    .B1(\core.registers[31][8] ),
    .B2(net1417),
    .C1(net1712),
    .X(_06283_));
 sky130_fd_sc_hd__o21a_1 _11371_ (.A1(net1876),
    .A2(_06282_),
    .B1(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__mux2_1 _11372_ (.A0(\core.registers[14][8] ),
    .A1(\core.registers[15][8] ),
    .S(net1417),
    .X(_06285_));
 sky130_fd_sc_hd__mux2_1 _11373_ (.A0(\core.registers[12][8] ),
    .A1(\core.registers[13][8] ),
    .S(net1417),
    .X(_06286_));
 sky130_fd_sc_hd__mux2_1 _11374_ (.A0(_06285_),
    .A1(_06286_),
    .S(net1474),
    .X(_06287_));
 sky130_fd_sc_hd__mux2_1 _11375_ (.A0(_06284_),
    .A1(_06287_),
    .S(net1717),
    .X(_06288_));
 sky130_fd_sc_hd__a22o_1 _11376_ (.A1(net1695),
    .A2(\core.registers[26][8] ),
    .B1(\core.registers[27][8] ),
    .B2(net1417),
    .X(_06289_));
 sky130_fd_sc_hd__mux2_1 _11377_ (.A0(\core.registers[24][8] ),
    .A1(\core.registers[25][8] ),
    .S(net1417),
    .X(_06290_));
 sky130_fd_sc_hd__mux2_1 _11378_ (.A0(_06289_),
    .A1(_06290_),
    .S(net1710),
    .X(_06291_));
 sky130_fd_sc_hd__or2_1 _11379_ (.A(\core.registers[9][8] ),
    .B(net1376),
    .X(_06292_));
 sky130_fd_sc_hd__o21a_1 _11380_ (.A1(\core.registers[8][8] ),
    .A2(net1417),
    .B1(net1709),
    .X(_06293_));
 sky130_fd_sc_hd__a22o_1 _11381_ (.A1(net1695),
    .A2(\core.registers[10][8] ),
    .B1(\core.registers[11][8] ),
    .B2(net1415),
    .X(_06294_));
 sky130_fd_sc_hd__a221o_1 _11382_ (.A1(_06292_),
    .A2(_06293_),
    .B1(_06294_),
    .B2(net1875),
    .C1(net1858),
    .X(_06295_));
 sky130_fd_sc_hd__o21a_1 _11383_ (.A1(net1717),
    .A2(_06291_),
    .B1(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__mux2_2 _11384_ (.A0(_06296_),
    .A1(_06288_),
    .S(net1865),
    .X(_06297_));
 sky130_fd_sc_hd__o22a_1 _11385_ (.A1(net1701),
    .A2(\core.registers[23][8] ),
    .B1(net1425),
    .B2(\core.registers[22][8] ),
    .X(_06298_));
 sky130_fd_sc_hd__or3_1 _11386_ (.A(net1701),
    .B(\core.registers[19][8] ),
    .C(net1459),
    .X(_06299_));
 sky130_fd_sc_hd__o221a_1 _11387_ (.A1(\core.registers[18][8] ),
    .A2(net1337),
    .B1(_06298_),
    .B2(net1440),
    .C1(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__mux4_1 _11388_ (.A0(\core.registers[16][8] ),
    .A1(\core.registers[17][8] ),
    .A2(\core.registers[20][8] ),
    .A3(\core.registers[21][8] ),
    .S0(net1424),
    .S1(net1459),
    .X(_06301_));
 sky130_fd_sc_hd__mux2_1 _11389_ (.A0(_06300_),
    .A1(_06301_),
    .S(net1475),
    .X(_06302_));
 sky130_fd_sc_hd__o22a_1 _11390_ (.A1(net1701),
    .A2(\core.registers[7][8] ),
    .B1(net1423),
    .B2(\core.registers[6][8] ),
    .X(_06303_));
 sky130_fd_sc_hd__or3_1 _11391_ (.A(net1701),
    .B(\core.registers[3][8] ),
    .C(net1459),
    .X(_06304_));
 sky130_fd_sc_hd__o221a_1 _11392_ (.A1(\core.registers[2][8] ),
    .A2(net1337),
    .B1(_06303_),
    .B2(net1440),
    .C1(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__mux4_1 _11393_ (.A0(\core.registers[0][8] ),
    .A1(\core.registers[1][8] ),
    .A2(\core.registers[4][8] ),
    .A3(\core.registers[5][8] ),
    .S0(net1425),
    .S1(net1459),
    .X(_06306_));
 sky130_fd_sc_hd__mux2_1 _11394_ (.A0(_06305_),
    .A1(_06306_),
    .S(net1475),
    .X(_06307_));
 sky130_fd_sc_hd__mux2_1 _11395_ (.A0(_06302_),
    .A1(_06307_),
    .S(net1463),
    .X(_06308_));
 sky130_fd_sc_hd__mux2_4 _11396_ (.A0(_06297_),
    .A1(_06308_),
    .S(net1488),
    .X(_06309_));
 sky130_fd_sc_hd__a22o_4 _11397_ (.A1(net1070),
    .A2(net961),
    .B1(_06309_),
    .B2(net1067),
    .X(_06310_));
 sky130_fd_sc_hd__mux2_2 _11398_ (.A0(net480),
    .A1(_06310_),
    .S(net1282),
    .X(_06311_));
 sky130_fd_sc_hd__and2_2 _11399_ (.A(_06281_),
    .B(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__nor2_1 _11400_ (.A(_06281_),
    .B(_06311_),
    .Y(_06313_));
 sky130_fd_sc_hd__nor2_2 _11401_ (.A(_06312_),
    .B(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__inv_2 _11402_ (.A(_06314_),
    .Y(_06315_));
 sky130_fd_sc_hd__o311a_4 _11403_ (.A1(_05717_),
    .A2(_06232_),
    .A3(_06236_),
    .B1(_06315_),
    .C1(_05718_),
    .X(_06316_));
 sky130_fd_sc_hd__and2b_2 _11404_ (.A_N(_06281_),
    .B(_06311_),
    .X(_06317_));
 sky130_fd_sc_hd__or2_1 _11405_ (.A(_05557_),
    .B(_06317_),
    .X(_06318_));
 sky130_fd_sc_hd__or3_1 _11406_ (.A(_05368_),
    .B(_05455_),
    .C(_05555_),
    .X(_06319_));
 sky130_fd_sc_hd__a21bo_1 _11407_ (.A1(_05552_),
    .A2(_06317_),
    .B1_N(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__a311o_1 _11408_ (.A1(_05369_),
    .A2(_05421_),
    .A3(_05452_),
    .B1(_05553_),
    .C1(_06320_),
    .X(_06321_));
 sky130_fd_sc_hd__and2_1 _11409_ (.A(_05281_),
    .B(net2012),
    .X(_06322_));
 sky130_fd_sc_hd__a31oi_4 _11410_ (.A1(_05281_),
    .A2(_05552_),
    .A3(_06316_),
    .B1(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__and2b_1 _11411_ (.A_N(_05078_),
    .B(_05108_),
    .X(_06324_));
 sky130_fd_sc_hd__and2b_1 _11412_ (.A_N(_04991_),
    .B(_05023_),
    .X(_06325_));
 sky130_fd_sc_hd__a21oi_2 _11413_ (.A1(_05111_),
    .A2(_06325_),
    .B1(_06324_),
    .Y(_06326_));
 sky130_fd_sc_hd__nand2b_1 _11414_ (.A_N(_05244_),
    .B(_05276_),
    .Y(_06327_));
 sky130_fd_sc_hd__or2_1 _11415_ (.A(_05192_),
    .B(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__nand2b_1 _11416_ (.A_N(_05157_),
    .B(_05187_),
    .Y(_06329_));
 sky130_fd_sc_hd__o311a_2 _11417_ (.A1(_05192_),
    .A2(_05280_),
    .A3(_06326_),
    .B1(_06328_),
    .C1(_06329_),
    .X(_06330_));
 sky130_fd_sc_hd__mux2_1 _11418_ (.A0(\core.registers[8][17] ),
    .A1(\core.registers[9][17] ),
    .S(net1515),
    .X(_06331_));
 sky130_fd_sc_hd__mux2_1 _11419_ (.A0(\core.registers[10][17] ),
    .A1(\core.registers[11][17] ),
    .S(net1516),
    .X(_06332_));
 sky130_fd_sc_hd__mux2_1 _11420_ (.A0(\core.registers[24][17] ),
    .A1(\core.registers[25][17] ),
    .S(net1520),
    .X(_06333_));
 sky130_fd_sc_hd__a221o_1 _11421_ (.A1(net1721),
    .A2(\core.registers[26][17] ),
    .B1(\core.registers[27][17] ),
    .B2(net1520),
    .C1(net1738),
    .X(_06334_));
 sky130_fd_sc_hd__or2_1 _11422_ (.A(\core.registers[29][17] ),
    .B(net1495),
    .X(_06335_));
 sky130_fd_sc_hd__o211a_1 _11423_ (.A1(\core.registers[28][17] ),
    .A2(net1520),
    .B1(_06335_),
    .C1(net1738),
    .X(_06336_));
 sky130_fd_sc_hd__a31o_1 _11424_ (.A1(net1840),
    .A2(net1721),
    .A3(\core.registers[30][17] ),
    .B1(net1748),
    .X(_06337_));
 sky130_fd_sc_hd__a31o_1 _11425_ (.A1(net1840),
    .A2(\core.registers[31][17] ),
    .A3(net1520),
    .B1(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__or2_1 _11426_ (.A(\core.registers[1][17] ),
    .B(net1494),
    .X(_06339_));
 sky130_fd_sc_hd__or2_1 _11427_ (.A(\core.registers[6][17] ),
    .B(net1518),
    .X(_06340_));
 sky130_fd_sc_hd__or2_1 _11428_ (.A(\core.registers[17][17] ),
    .B(net1494),
    .X(_06341_));
 sky130_fd_sc_hd__mux2_1 _11429_ (.A0(\core.registers[12][17] ),
    .A1(\core.registers[13][17] ),
    .S(net1514),
    .X(_06342_));
 sky130_fd_sc_hd__mux2_1 _11430_ (.A0(\core.registers[14][17] ),
    .A1(\core.registers[15][17] ),
    .S(net1514),
    .X(_06343_));
 sky130_fd_sc_hd__mux2_2 _11431_ (.A0(_06342_),
    .A1(_06343_),
    .S(net1614),
    .X(_06344_));
 sky130_fd_sc_hd__o221a_1 _11432_ (.A1(_06336_),
    .A2(_06338_),
    .B1(_06344_),
    .B2(net1825),
    .C1(net1832),
    .X(_06345_));
 sky130_fd_sc_hd__mux2_1 _11433_ (.A0(_06331_),
    .A1(_06332_),
    .S(net1614),
    .X(_06346_));
 sky130_fd_sc_hd__o21a_1 _11434_ (.A1(net1843),
    .A2(_06333_),
    .B1(_06334_),
    .X(_06347_));
 sky130_fd_sc_hd__mux2_1 _11435_ (.A0(_06346_),
    .A1(_06347_),
    .S(net1825),
    .X(_06348_));
 sky130_fd_sc_hd__a211o_1 _11436_ (.A1(net1744),
    .A2(_06348_),
    .B1(_06345_),
    .C1(net1631),
    .X(_06349_));
 sky130_fd_sc_hd__o211a_1 _11437_ (.A1(net1721),
    .A2(\core.registers[7][17] ),
    .B1(net1614),
    .C1(_06340_),
    .X(_06350_));
 sky130_fd_sc_hd__mux2_1 _11438_ (.A0(\core.registers[4][17] ),
    .A1(\core.registers[5][17] ),
    .S(net1517),
    .X(_06351_));
 sky130_fd_sc_hd__a211o_1 _11439_ (.A1(net1599),
    .A2(_06351_),
    .B1(_06350_),
    .C1(net1575),
    .X(_06352_));
 sky130_fd_sc_hd__o211a_1 _11440_ (.A1(\core.registers[0][17] ),
    .A2(net1519),
    .B1(_06339_),
    .C1(net1600),
    .X(_06353_));
 sky130_fd_sc_hd__mux2_1 _11441_ (.A0(\core.registers[2][17] ),
    .A1(\core.registers[3][17] ),
    .S(net1518),
    .X(_06354_));
 sky130_fd_sc_hd__a211o_1 _11442_ (.A1(net1615),
    .A2(_06354_),
    .B1(_06353_),
    .C1(net1586),
    .X(_06355_));
 sky130_fd_sc_hd__o211a_1 _11443_ (.A1(\core.registers[16][17] ),
    .A2(net1517),
    .B1(_06341_),
    .C1(net1599),
    .X(_06356_));
 sky130_fd_sc_hd__mux2_1 _11444_ (.A0(\core.registers[18][17] ),
    .A1(\core.registers[19][17] ),
    .S(net1517),
    .X(_06357_));
 sky130_fd_sc_hd__a211o_1 _11445_ (.A1(net1615),
    .A2(_06357_),
    .B1(_06356_),
    .C1(net1587),
    .X(_06358_));
 sky130_fd_sc_hd__mux2_1 _11446_ (.A0(\core.registers[22][17] ),
    .A1(\core.registers[23][17] ),
    .S(net1518),
    .X(_06359_));
 sky130_fd_sc_hd__mux2_1 _11447_ (.A0(\core.registers[20][17] ),
    .A1(\core.registers[21][17] ),
    .S(net1517),
    .X(_06360_));
 sky130_fd_sc_hd__mux2_1 _11448_ (.A0(_06359_),
    .A1(_06360_),
    .S(net1599),
    .X(_06361_));
 sky130_fd_sc_hd__o211a_1 _11449_ (.A1(net1575),
    .A2(_06361_),
    .B1(_06358_),
    .C1(net1571),
    .X(_06362_));
 sky130_fd_sc_hd__a311o_2 _11450_ (.A1(net1567),
    .A2(_06352_),
    .A3(_06355_),
    .B1(_06362_),
    .C1(net1635),
    .X(_06363_));
 sky130_fd_sc_hd__a21o_1 _11451_ (.A1(_06349_),
    .A2(_06363_),
    .B1(net1157),
    .X(_06364_));
 sky130_fd_sc_hd__a21o_4 _11452_ (.A1(net1234),
    .A2(_05465_),
    .B1(net1236),
    .X(_06365_));
 sky130_fd_sc_hd__a22o_1 _11453_ (.A1(\core.pipe1_resultRegister[17] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[17] ),
    .X(_06366_));
 sky130_fd_sc_hd__a21o_2 _11454_ (.A1(net1188),
    .A2(_06365_),
    .B1(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__o211ai_2 _11455_ (.A1(net1153),
    .A2(_06367_),
    .B1(_06364_),
    .C1(net1263),
    .Y(_06368_));
 sky130_fd_sc_hd__o21ai_1 _11456_ (.A1(net1192),
    .A2(_06368_),
    .B1(net1161),
    .Y(_06369_));
 sky130_fd_sc_hd__o21a_1 _11457_ (.A1(net1863),
    .A2(net1278),
    .B1(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__and3_1 _11458_ (.A(\core.pipe0_currentInstruction[15] ),
    .B(\core.registers[23][17] ),
    .C(net1666),
    .X(_06371_));
 sky130_fd_sc_hd__mux2_1 _11459_ (.A0(\core.registers[28][17] ),
    .A1(\core.registers[29][17] ),
    .S(net1392),
    .X(_06372_));
 sky130_fd_sc_hd__mux2_1 _11460_ (.A0(\core.registers[30][17] ),
    .A1(\core.registers[31][17] ),
    .S(net1392),
    .X(_06373_));
 sky130_fd_sc_hd__mux2_1 _11461_ (.A0(_06372_),
    .A1(_06373_),
    .S(net1479),
    .X(_06374_));
 sky130_fd_sc_hd__mux2_1 _11462_ (.A0(\core.registers[26][17] ),
    .A1(\core.registers[27][17] ),
    .S(net1392),
    .X(_06375_));
 sky130_fd_sc_hd__mux2_1 _11463_ (.A0(\core.registers[24][17] ),
    .A1(\core.registers[25][17] ),
    .S(net1392),
    .X(_06376_));
 sky130_fd_sc_hd__or2_1 _11464_ (.A(net1479),
    .B(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__o211a_1 _11465_ (.A1(net1468),
    .A2(_06375_),
    .B1(_06377_),
    .C1(net1437),
    .X(_06378_));
 sky130_fd_sc_hd__a211o_2 _11466_ (.A1(net1446),
    .A2(_06374_),
    .B1(_06378_),
    .C1(net1484),
    .X(_06379_));
 sky130_fd_sc_hd__a211o_1 _11467_ (.A1(net1682),
    .A2(\core.registers[22][17] ),
    .B1(net1468),
    .C1(_06371_),
    .X(_06380_));
 sky130_fd_sc_hd__mux2_1 _11468_ (.A0(\core.registers[20][17] ),
    .A1(\core.registers[21][17] ),
    .S(net1390),
    .X(_06381_));
 sky130_fd_sc_hd__o211a_1 _11469_ (.A1(net1478),
    .A2(_06381_),
    .B1(_06380_),
    .C1(net1445),
    .X(_06382_));
 sky130_fd_sc_hd__mux2_1 _11470_ (.A0(\core.registers[16][17] ),
    .A1(\core.registers[17][17] ),
    .S(net1390),
    .X(_06383_));
 sky130_fd_sc_hd__or2_1 _11471_ (.A(net1478),
    .B(_06383_),
    .X(_06384_));
 sky130_fd_sc_hd__mux2_1 _11472_ (.A0(\core.registers[18][17] ),
    .A1(\core.registers[19][17] ),
    .S(net1390),
    .X(_06385_));
 sky130_fd_sc_hd__o211a_1 _11473_ (.A1(net1467),
    .A2(_06385_),
    .B1(_06384_),
    .C1(net1434),
    .X(_06386_));
 sky130_fd_sc_hd__o311a_1 _11474_ (.A1(net1489),
    .A2(_06382_),
    .A3(_06386_),
    .B1(net1464),
    .C1(_06379_),
    .X(_06387_));
 sky130_fd_sc_hd__mux2_1 _11475_ (.A0(\core.registers[2][17] ),
    .A1(\core.registers[3][17] ),
    .S(net1391),
    .X(_06388_));
 sky130_fd_sc_hd__mux2_1 _11476_ (.A0(\core.registers[0][17] ),
    .A1(\core.registers[1][17] ),
    .S(net1391),
    .X(_06389_));
 sky130_fd_sc_hd__or2_1 _11477_ (.A(net1479),
    .B(_06389_),
    .X(_06390_));
 sky130_fd_sc_hd__o211a_1 _11478_ (.A1(net1468),
    .A2(_06388_),
    .B1(_06390_),
    .C1(net1434),
    .X(_06391_));
 sky130_fd_sc_hd__mux2_1 _11479_ (.A0(\core.registers[4][17] ),
    .A1(\core.registers[5][17] ),
    .S(net1390),
    .X(_06392_));
 sky130_fd_sc_hd__mux2_1 _11480_ (.A0(\core.registers[6][17] ),
    .A1(\core.registers[7][17] ),
    .S(net1391),
    .X(_06393_));
 sky130_fd_sc_hd__mux2_1 _11481_ (.A0(_06392_),
    .A1(_06393_),
    .S(net1478),
    .X(_06394_));
 sky130_fd_sc_hd__a211o_1 _11482_ (.A1(net1446),
    .A2(_06394_),
    .B1(_06391_),
    .C1(net1490),
    .X(_06395_));
 sky130_fd_sc_hd__mux2_1 _11483_ (.A0(\core.registers[10][17] ),
    .A1(\core.registers[11][17] ),
    .S(net1389),
    .X(_06396_));
 sky130_fd_sc_hd__mux2_1 _11484_ (.A0(\core.registers[8][17] ),
    .A1(\core.registers[9][17] ),
    .S(net1389),
    .X(_06397_));
 sky130_fd_sc_hd__or2_1 _11485_ (.A(net1478),
    .B(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__o211a_1 _11486_ (.A1(net1467),
    .A2(_06396_),
    .B1(_06398_),
    .C1(net1434),
    .X(_06399_));
 sky130_fd_sc_hd__mux2_1 _11487_ (.A0(\core.registers[12][17] ),
    .A1(\core.registers[13][17] ),
    .S(net1388),
    .X(_06400_));
 sky130_fd_sc_hd__mux2_1 _11488_ (.A0(\core.registers[14][17] ),
    .A1(\core.registers[15][17] ),
    .S(net1388),
    .X(_06401_));
 sky130_fd_sc_hd__mux2_1 _11489_ (.A0(_06400_),
    .A1(_06401_),
    .S(net1478),
    .X(_06402_));
 sky130_fd_sc_hd__a211o_1 _11490_ (.A1(net1445),
    .A2(_06402_),
    .B1(_06399_),
    .C1(net1485),
    .X(_06403_));
 sky130_fd_sc_hd__a31o_1 _11491_ (.A1(net1460),
    .A2(_06395_),
    .A3(_06403_),
    .B1(_06387_),
    .X(_06404_));
 sky130_fd_sc_hd__a22o_2 _11492_ (.A1(net1068),
    .A2(net1131),
    .B1(_06404_),
    .B2(net1065),
    .X(_06405_));
 sky130_fd_sc_hd__mux2_4 _11493_ (.A0(net458),
    .A1(_06405_),
    .S(net1279),
    .X(_06406_));
 sky130_fd_sc_hd__or2_2 _11494_ (.A(_06370_),
    .B(_06406_),
    .X(_06407_));
 sky130_fd_sc_hd__nand2_1 _11495_ (.A(_06370_),
    .B(_06406_),
    .Y(_06408_));
 sky130_fd_sc_hd__inv_2 _11496_ (.A(_06408_),
    .Y(_06409_));
 sky130_fd_sc_hd__and2_4 _11497_ (.A(_06407_),
    .B(_06408_),
    .X(_06410_));
 sky130_fd_sc_hd__or2_1 _11498_ (.A(\core.registers[1][16] ),
    .B(net1494),
    .X(_06411_));
 sky130_fd_sc_hd__or2_1 _11499_ (.A(\core.registers[6][16] ),
    .B(net1514),
    .X(_06412_));
 sky130_fd_sc_hd__or2_1 _11500_ (.A(\core.registers[17][16] ),
    .B(net1493),
    .X(_06413_));
 sky130_fd_sc_hd__or2_1 _11501_ (.A(\core.registers[28][16] ),
    .B(net1507),
    .X(_06414_));
 sky130_fd_sc_hd__o211a_1 _11502_ (.A1(\core.registers[29][16] ),
    .A2(net1493),
    .B1(_06414_),
    .C1(net1736),
    .X(_06415_));
 sky130_fd_sc_hd__a31o_1 _11503_ (.A1(net1840),
    .A2(net1719),
    .A3(\core.registers[30][16] ),
    .B1(net1749),
    .X(_06416_));
 sky130_fd_sc_hd__a31o_1 _11504_ (.A1(net1840),
    .A2(\core.registers[31][16] ),
    .A3(net1508),
    .B1(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__mux2_1 _11505_ (.A0(\core.registers[8][16] ),
    .A1(\core.registers[9][16] ),
    .S(net1506),
    .X(_06418_));
 sky130_fd_sc_hd__mux2_1 _11506_ (.A0(\core.registers[10][16] ),
    .A1(\core.registers[11][16] ),
    .S(net1506),
    .X(_06419_));
 sky130_fd_sc_hd__mux2_1 _11507_ (.A0(\core.registers[24][16] ),
    .A1(\core.registers[25][16] ),
    .S(net1507),
    .X(_06420_));
 sky130_fd_sc_hd__a221o_1 _11508_ (.A1(net1720),
    .A2(\core.registers[26][16] ),
    .B1(\core.registers[27][16] ),
    .B2(net1507),
    .C1(net1735),
    .X(_06421_));
 sky130_fd_sc_hd__mux2_1 _11509_ (.A0(\core.registers[12][16] ),
    .A1(\core.registers[13][16] ),
    .S(net1506),
    .X(_06422_));
 sky130_fd_sc_hd__mux2_1 _11510_ (.A0(\core.registers[14][16] ),
    .A1(\core.registers[15][16] ),
    .S(net1507),
    .X(_06423_));
 sky130_fd_sc_hd__mux2_1 _11511_ (.A0(_06422_),
    .A1(_06423_),
    .S(net1611),
    .X(_06424_));
 sky130_fd_sc_hd__o221a_1 _11512_ (.A1(_06415_),
    .A2(_06417_),
    .B1(_06424_),
    .B2(net1824),
    .C1(net1832),
    .X(_06425_));
 sky130_fd_sc_hd__mux2_1 _11513_ (.A0(_06418_),
    .A1(_06419_),
    .S(net1613),
    .X(_06426_));
 sky130_fd_sc_hd__o21a_1 _11514_ (.A1(net1840),
    .A2(_06420_),
    .B1(_06421_),
    .X(_06427_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(_06426_),
    .A1(_06427_),
    .S(net1824),
    .X(_06428_));
 sky130_fd_sc_hd__a211o_1 _11516_ (.A1(net1744),
    .A2(_06428_),
    .B1(_06425_),
    .C1(net1631),
    .X(_06429_));
 sky130_fd_sc_hd__o211a_1 _11517_ (.A1(net1719),
    .A2(\core.registers[7][16] ),
    .B1(net1614),
    .C1(_06412_),
    .X(_06430_));
 sky130_fd_sc_hd__mux2_1 _11518_ (.A0(\core.registers[4][16] ),
    .A1(\core.registers[5][16] ),
    .S(net1514),
    .X(_06431_));
 sky130_fd_sc_hd__a211o_1 _11519_ (.A1(net1598),
    .A2(_06431_),
    .B1(_06430_),
    .C1(net1575),
    .X(_06432_));
 sky130_fd_sc_hd__o211a_1 _11520_ (.A1(\core.registers[0][16] ),
    .A2(net1514),
    .B1(_06411_),
    .C1(net1600),
    .X(_06433_));
 sky130_fd_sc_hd__mux2_1 _11521_ (.A0(\core.registers[2][16] ),
    .A1(\core.registers[3][16] ),
    .S(net1514),
    .X(_06434_));
 sky130_fd_sc_hd__a211o_1 _11522_ (.A1(net1611),
    .A2(_06434_),
    .B1(_06433_),
    .C1(net1586),
    .X(_06435_));
 sky130_fd_sc_hd__o211a_1 _11523_ (.A1(\core.registers[16][16] ),
    .A2(net1506),
    .B1(_06413_),
    .C1(net1598),
    .X(_06436_));
 sky130_fd_sc_hd__mux2_1 _11524_ (.A0(\core.registers[18][16] ),
    .A1(\core.registers[19][16] ),
    .S(net1506),
    .X(_06437_));
 sky130_fd_sc_hd__a211o_1 _11525_ (.A1(net1611),
    .A2(_06437_),
    .B1(_06436_),
    .C1(net1586),
    .X(_06438_));
 sky130_fd_sc_hd__mux2_1 _11526_ (.A0(\core.registers[22][16] ),
    .A1(\core.registers[23][16] ),
    .S(net1507),
    .X(_06439_));
 sky130_fd_sc_hd__mux2_1 _11527_ (.A0(\core.registers[20][16] ),
    .A1(\core.registers[21][16] ),
    .S(net1506),
    .X(_06440_));
 sky130_fd_sc_hd__mux2_1 _11528_ (.A0(_06439_),
    .A1(_06440_),
    .S(net1598),
    .X(_06441_));
 sky130_fd_sc_hd__o211a_1 _11529_ (.A1(net1575),
    .A2(_06441_),
    .B1(_06438_),
    .C1(net1571),
    .X(_06442_));
 sky130_fd_sc_hd__a311o_1 _11530_ (.A1(net1567),
    .A2(_06432_),
    .A3(_06435_),
    .B1(_06442_),
    .C1(net1635),
    .X(_06443_));
 sky130_fd_sc_hd__a21o_2 _11531_ (.A1(_06429_),
    .A2(_06443_),
    .B1(net1157),
    .X(_06444_));
 sky130_fd_sc_hd__a21o_4 _11532_ (.A1(net1234),
    .A2(_06156_),
    .B1(net2014),
    .X(_06445_));
 sky130_fd_sc_hd__a22o_1 _11533_ (.A1(\core.pipe1_resultRegister[16] ),
    .A2(net1240),
    .B1(_04520_),
    .B2(\core.pipe1_csrData[16] ),
    .X(_06446_));
 sky130_fd_sc_hd__a21o_4 _11534_ (.A1(net1191),
    .A2(_06445_),
    .B1(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__o211ai_4 _11535_ (.A1(net1153),
    .A2(_06447_),
    .B1(_06444_),
    .C1(net1263),
    .Y(_06448_));
 sky130_fd_sc_hd__o21a_1 _11536_ (.A1(net1193),
    .A2(_06448_),
    .B1(net1162),
    .X(_06449_));
 sky130_fd_sc_hd__a21oi_2 _11537_ (.A1(net1714),
    .A2(net1286),
    .B1(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__or2_1 _11538_ (.A(\core.registers[13][16] ),
    .B(net1373),
    .X(_06451_));
 sky130_fd_sc_hd__o211a_1 _11539_ (.A1(\core.registers[12][16] ),
    .A2(net1381),
    .B1(_06451_),
    .C1(net1444),
    .X(_06452_));
 sky130_fd_sc_hd__a31o_1 _11540_ (.A1(\core.registers[9][16] ),
    .A2(net1431),
    .A3(net1381),
    .B1(net1480),
    .X(_06453_));
 sky130_fd_sc_hd__a311o_1 _11541_ (.A1(\core.registers[8][16] ),
    .A2(net1431),
    .A3(net1373),
    .B1(_06452_),
    .C1(_06453_),
    .X(_06454_));
 sky130_fd_sc_hd__a22o_1 _11542_ (.A1(net1677),
    .A2(\core.registers[10][16] ),
    .B1(\core.registers[11][16] ),
    .B2(net1381),
    .X(_06455_));
 sky130_fd_sc_hd__a22o_1 _11543_ (.A1(net1677),
    .A2(\core.registers[14][16] ),
    .B1(\core.registers[15][16] ),
    .B2(net1381),
    .X(_06456_));
 sky130_fd_sc_hd__a21o_1 _11544_ (.A1(net1444),
    .A2(_06456_),
    .B1(net1465),
    .X(_06457_));
 sky130_fd_sc_hd__a21o_1 _11545_ (.A1(net1431),
    .A2(_06455_),
    .B1(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__a22o_1 _11546_ (.A1(net1677),
    .A2(\core.registers[6][16] ),
    .B1(\core.registers[7][16] ),
    .B2(net1388),
    .X(_06459_));
 sky130_fd_sc_hd__a22o_1 _11547_ (.A1(net1677),
    .A2(\core.registers[2][16] ),
    .B1(\core.registers[3][16] ),
    .B2(net1388),
    .X(_06460_));
 sky130_fd_sc_hd__mux2_1 _11548_ (.A0(_06459_),
    .A1(_06460_),
    .S(net1431),
    .X(_06461_));
 sky130_fd_sc_hd__mux4_1 _11549_ (.A0(\core.registers[0][16] ),
    .A1(\core.registers[1][16] ),
    .A2(\core.registers[4][16] ),
    .A3(\core.registers[5][16] ),
    .S0(net1388),
    .S1(net1444),
    .X(_06462_));
 sky130_fd_sc_hd__a31o_1 _11550_ (.A1(net1485),
    .A2(net1465),
    .A3(_06462_),
    .B1(net1464),
    .X(_06463_));
 sky130_fd_sc_hd__a31o_1 _11551_ (.A1(net1485),
    .A2(net1480),
    .A3(_06461_),
    .B1(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__a31o_2 _11552_ (.A1(net1489),
    .A2(_06454_),
    .A3(_06458_),
    .B1(_06464_),
    .X(_06465_));
 sky130_fd_sc_hd__or2_1 _11553_ (.A(\core.registers[29][16] ),
    .B(net1373),
    .X(_06466_));
 sky130_fd_sc_hd__o211a_1 _11554_ (.A1(\core.registers[28][16] ),
    .A2(net1382),
    .B1(_06466_),
    .C1(net1444),
    .X(_06467_));
 sky130_fd_sc_hd__a31o_1 _11555_ (.A1(\core.registers[25][16] ),
    .A2(net1431),
    .A3(net1382),
    .B1(net1480),
    .X(_06468_));
 sky130_fd_sc_hd__a311o_1 _11556_ (.A1(\core.registers[24][16] ),
    .A2(net1431),
    .A3(net1373),
    .B1(_06467_),
    .C1(_06468_),
    .X(_06469_));
 sky130_fd_sc_hd__a22o_1 _11557_ (.A1(net1683),
    .A2(\core.registers[26][16] ),
    .B1(\core.registers[27][16] ),
    .B2(net1382),
    .X(_06470_));
 sky130_fd_sc_hd__a22o_1 _11558_ (.A1(net1678),
    .A2(\core.registers[30][16] ),
    .B1(\core.registers[31][16] ),
    .B2(net1387),
    .X(_06471_));
 sky130_fd_sc_hd__a21o_1 _11559_ (.A1(net1444),
    .A2(_06471_),
    .B1(net1465),
    .X(_06472_));
 sky130_fd_sc_hd__a21o_1 _11560_ (.A1(net1433),
    .A2(_06470_),
    .B1(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__a22o_1 _11561_ (.A1(net1677),
    .A2(\core.registers[22][16] ),
    .B1(\core.registers[23][16] ),
    .B2(net1381),
    .X(_06474_));
 sky130_fd_sc_hd__a22o_1 _11562_ (.A1(net1677),
    .A2(\core.registers[18][16] ),
    .B1(\core.registers[19][16] ),
    .B2(net1381),
    .X(_06475_));
 sky130_fd_sc_hd__mux2_1 _11563_ (.A0(_06474_),
    .A1(_06475_),
    .S(net1431),
    .X(_06476_));
 sky130_fd_sc_hd__mux4_2 _11564_ (.A0(\core.registers[16][16] ),
    .A1(\core.registers[17][16] ),
    .A2(\core.registers[20][16] ),
    .A3(\core.registers[21][16] ),
    .S0(net1382),
    .S1(net1444),
    .X(_06477_));
 sky130_fd_sc_hd__a31o_1 _11565_ (.A1(net1484),
    .A2(net1465),
    .A3(_06477_),
    .B1(net1460),
    .X(_06478_));
 sky130_fd_sc_hd__a31o_1 _11566_ (.A1(net1485),
    .A2(net1480),
    .A3(_06476_),
    .B1(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__a31o_1 _11567_ (.A1(net1489),
    .A2(_06469_),
    .A3(_06473_),
    .B1(_06479_),
    .X(_06480_));
 sky130_fd_sc_hd__nand2_4 _11568_ (.A(_06465_),
    .B(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__o2bb2a_1 _11569_ (.A1_N(net1068),
    .A2_N(_06447_),
    .B1(_06481_),
    .B2(_04663_),
    .X(_06482_));
 sky130_fd_sc_hd__inv_2 _11570_ (.A(_06482_),
    .Y(_06483_));
 sky130_fd_sc_hd__mux2_4 _11571_ (.A0(net457),
    .A1(_06483_),
    .S(net1279),
    .X(_06484_));
 sky130_fd_sc_hd__nor2_2 _11572_ (.A(_06450_),
    .B(_06484_),
    .Y(_06485_));
 sky130_fd_sc_hd__inv_2 _11573_ (.A(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__and2_2 _11574_ (.A(_06450_),
    .B(_06484_),
    .X(_06487_));
 sky130_fd_sc_hd__nor2_4 _11575_ (.A(_06485_),
    .B(_06487_),
    .Y(_06488_));
 sky130_fd_sc_hd__mux2_1 _11576_ (.A0(\core.registers[8][19] ),
    .A1(\core.registers[9][19] ),
    .S(net1513),
    .X(_06489_));
 sky130_fd_sc_hd__mux2_1 _11577_ (.A0(\core.registers[10][19] ),
    .A1(\core.registers[11][19] ),
    .S(net1510),
    .X(_06490_));
 sky130_fd_sc_hd__mux2_1 _11578_ (.A0(\core.registers[24][19] ),
    .A1(\core.registers[25][19] ),
    .S(net1524),
    .X(_06491_));
 sky130_fd_sc_hd__a221o_1 _11579_ (.A1(net1722),
    .A2(\core.registers[26][19] ),
    .B1(\core.registers[27][19] ),
    .B2(net1524),
    .C1(net1736),
    .X(_06492_));
 sky130_fd_sc_hd__or2_1 _11580_ (.A(\core.registers[28][19] ),
    .B(net1524),
    .X(_06493_));
 sky130_fd_sc_hd__o211a_1 _11581_ (.A1(\core.registers[29][19] ),
    .A2(net1496),
    .B1(_06493_),
    .C1(net1736),
    .X(_06494_));
 sky130_fd_sc_hd__a31o_1 _11582_ (.A1(net1839),
    .A2(net1720),
    .A3(\core.registers[30][19] ),
    .B1(net1748),
    .X(_06495_));
 sky130_fd_sc_hd__a31o_1 _11583_ (.A1(net1839),
    .A2(\core.registers[31][19] ),
    .A3(net1510),
    .B1(_06495_),
    .X(_06496_));
 sky130_fd_sc_hd__or2_1 _11584_ (.A(\core.registers[1][19] ),
    .B(net1493),
    .X(_06497_));
 sky130_fd_sc_hd__or2_1 _11585_ (.A(\core.registers[6][19] ),
    .B(net1512),
    .X(_06498_));
 sky130_fd_sc_hd__or2_1 _11586_ (.A(\core.registers[17][19] ),
    .B(net1495),
    .X(_06499_));
 sky130_fd_sc_hd__mux2_1 _11587_ (.A0(\core.registers[12][19] ),
    .A1(\core.registers[13][19] ),
    .S(net1510),
    .X(_06500_));
 sky130_fd_sc_hd__mux2_1 _11588_ (.A0(\core.registers[14][19] ),
    .A1(\core.registers[15][19] ),
    .S(net1510),
    .X(_06501_));
 sky130_fd_sc_hd__mux2_1 _11589_ (.A0(_06500_),
    .A1(_06501_),
    .S(net1612),
    .X(_06502_));
 sky130_fd_sc_hd__o221a_1 _11590_ (.A1(_06494_),
    .A2(_06496_),
    .B1(_06502_),
    .B2(net1824),
    .C1(net1832),
    .X(_06503_));
 sky130_fd_sc_hd__mux2_1 _11591_ (.A0(_06489_),
    .A1(_06490_),
    .S(net1612),
    .X(_06504_));
 sky130_fd_sc_hd__o21a_1 _11592_ (.A1(net1839),
    .A2(_06491_),
    .B1(_06492_),
    .X(_06505_));
 sky130_fd_sc_hd__mux2_1 _11593_ (.A0(_06504_),
    .A1(_06505_),
    .S(net1824),
    .X(_06506_));
 sky130_fd_sc_hd__a211o_1 _11594_ (.A1(net1744),
    .A2(_06506_),
    .B1(_06503_),
    .C1(net1631),
    .X(_06507_));
 sky130_fd_sc_hd__o211a_1 _11595_ (.A1(net1721),
    .A2(\core.registers[7][19] ),
    .B1(net1612),
    .C1(_06498_),
    .X(_06508_));
 sky130_fd_sc_hd__mux2_1 _11596_ (.A0(\core.registers[4][19] ),
    .A1(\core.registers[5][19] ),
    .S(net1513),
    .X(_06509_));
 sky130_fd_sc_hd__a211o_1 _11597_ (.A1(net1597),
    .A2(_06509_),
    .B1(_06508_),
    .C1(net1585),
    .X(_06510_));
 sky130_fd_sc_hd__o211a_1 _11598_ (.A1(\core.registers[0][19] ),
    .A2(net1512),
    .B1(_06497_),
    .C1(net1597),
    .X(_06511_));
 sky130_fd_sc_hd__mux2_1 _11599_ (.A0(\core.registers[2][19] ),
    .A1(\core.registers[3][19] ),
    .S(net1513),
    .X(_06512_));
 sky130_fd_sc_hd__a211o_1 _11600_ (.A1(net1612),
    .A2(_06512_),
    .B1(_06511_),
    .C1(net1596),
    .X(_06513_));
 sky130_fd_sc_hd__o211a_1 _11601_ (.A1(\core.registers[16][19] ),
    .A2(net1512),
    .B1(_06499_),
    .C1(net1598),
    .X(_06514_));
 sky130_fd_sc_hd__mux2_1 _11602_ (.A0(\core.registers[18][19] ),
    .A1(\core.registers[19][19] ),
    .S(net1512),
    .X(_06515_));
 sky130_fd_sc_hd__a211o_1 _11603_ (.A1(net1612),
    .A2(_06515_),
    .B1(_06514_),
    .C1(net1587),
    .X(_06516_));
 sky130_fd_sc_hd__mux2_1 _11604_ (.A0(\core.registers[22][19] ),
    .A1(\core.registers[23][19] ),
    .S(net1512),
    .X(_06517_));
 sky130_fd_sc_hd__mux2_1 _11605_ (.A0(\core.registers[20][19] ),
    .A1(\core.registers[21][19] ),
    .S(net1512),
    .X(_06518_));
 sky130_fd_sc_hd__mux2_1 _11606_ (.A0(_06517_),
    .A1(_06518_),
    .S(net1597),
    .X(_06519_));
 sky130_fd_sc_hd__o211a_1 _11607_ (.A1(net1576),
    .A2(_06519_),
    .B1(_06516_),
    .C1(net1571),
    .X(_06520_));
 sky130_fd_sc_hd__a311o_1 _11608_ (.A1(net1567),
    .A2(_06510_),
    .A3(_06513_),
    .B1(_06520_),
    .C1(net1635),
    .X(_06521_));
 sky130_fd_sc_hd__a21o_1 _11609_ (.A1(_06507_),
    .A2(_06521_),
    .B1(net1157),
    .X(_06522_));
 sky130_fd_sc_hd__a21o_4 _11610_ (.A1(net1234),
    .A2(_05289_),
    .B1(net1237),
    .X(_06523_));
 sky130_fd_sc_hd__a22o_1 _11611_ (.A1(\core.pipe1_resultRegister[19] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[19] ),
    .X(_06524_));
 sky130_fd_sc_hd__a21o_1 _11612_ (.A1(net1188),
    .A2(_06523_),
    .B1(_06524_),
    .X(_06525_));
 sky130_fd_sc_hd__o211ai_2 _11613_ (.A1(net1153),
    .A2(net1123),
    .B1(_06522_),
    .C1(net1263),
    .Y(_06526_));
 sky130_fd_sc_hd__o21ai_1 _11614_ (.A1(net1192),
    .A2(_06526_),
    .B1(net1161),
    .Y(_06527_));
 sky130_fd_sc_hd__o21a_1 _11615_ (.A1(net1855),
    .A2(net1278),
    .B1(_06527_),
    .X(_06528_));
 sky130_fd_sc_hd__or2_1 _11616_ (.A(\core.registers[13][19] ),
    .B(net1373),
    .X(_06529_));
 sky130_fd_sc_hd__o211a_1 _11617_ (.A1(\core.registers[12][19] ),
    .A2(net1384),
    .B1(_06529_),
    .C1(net1442),
    .X(_06530_));
 sky130_fd_sc_hd__a31o_1 _11618_ (.A1(\core.registers[9][19] ),
    .A2(net1432),
    .A3(net1384),
    .B1(net1480),
    .X(_06531_));
 sky130_fd_sc_hd__a311o_1 _11619_ (.A1(\core.registers[8][19] ),
    .A2(net1432),
    .A3(net1378),
    .B1(_06530_),
    .C1(_06531_),
    .X(_06532_));
 sky130_fd_sc_hd__a22o_1 _11620_ (.A1(net1681),
    .A2(\core.registers[10][19] ),
    .B1(\core.registers[11][19] ),
    .B2(net1384),
    .X(_06533_));
 sky130_fd_sc_hd__a22o_1 _11621_ (.A1(net1679),
    .A2(\core.registers[14][19] ),
    .B1(\core.registers[15][19] ),
    .B2(net1384),
    .X(_06534_));
 sky130_fd_sc_hd__a21o_1 _11622_ (.A1(net1442),
    .A2(_06534_),
    .B1(net1466),
    .X(_06535_));
 sky130_fd_sc_hd__a21o_1 _11623_ (.A1(net1432),
    .A2(_06533_),
    .B1(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__a22o_1 _11624_ (.A1(net1680),
    .A2(\core.registers[6][19] ),
    .B1(\core.registers[7][19] ),
    .B2(net1385),
    .X(_06537_));
 sky130_fd_sc_hd__a22o_1 _11625_ (.A1(net1680),
    .A2(\core.registers[2][19] ),
    .B1(\core.registers[3][19] ),
    .B2(net1386),
    .X(_06538_));
 sky130_fd_sc_hd__mux2_1 _11626_ (.A0(_06537_),
    .A1(_06538_),
    .S(net1432),
    .X(_06539_));
 sky130_fd_sc_hd__mux4_1 _11627_ (.A0(\core.registers[0][19] ),
    .A1(\core.registers[1][19] ),
    .A2(\core.registers[4][19] ),
    .A3(\core.registers[5][19] ),
    .S0(net1385),
    .S1(net1443),
    .X(_06540_));
 sky130_fd_sc_hd__a31o_1 _11628_ (.A1(net1485),
    .A2(net1466),
    .A3(_06540_),
    .B1(net1464),
    .X(_06541_));
 sky130_fd_sc_hd__a31o_1 _11629_ (.A1(net1484),
    .A2(net1481),
    .A3(_06539_),
    .B1(_06541_),
    .X(_06542_));
 sky130_fd_sc_hd__a31o_1 _11630_ (.A1(net1489),
    .A2(_06532_),
    .A3(_06536_),
    .B1(_06542_),
    .X(_06543_));
 sky130_fd_sc_hd__or2_1 _11631_ (.A(\core.registers[29][19] ),
    .B(net1374),
    .X(_06544_));
 sky130_fd_sc_hd__o211a_1 _11632_ (.A1(\core.registers[28][19] ),
    .A2(net1395),
    .B1(_06544_),
    .C1(net1447),
    .X(_06545_));
 sky130_fd_sc_hd__a31o_1 _11633_ (.A1(\core.registers[25][19] ),
    .A2(net1432),
    .A3(net1396),
    .B1(net1481),
    .X(_06546_));
 sky130_fd_sc_hd__a311o_1 _11634_ (.A1(\core.registers[24][19] ),
    .A2(net1432),
    .A3(net1374),
    .B1(_06545_),
    .C1(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__a22o_1 _11635_ (.A1(net1684),
    .A2(\core.registers[26][19] ),
    .B1(\core.registers[27][19] ),
    .B2(net1395),
    .X(_06548_));
 sky130_fd_sc_hd__a22o_1 _11636_ (.A1(net1679),
    .A2(\core.registers[30][19] ),
    .B1(\core.registers[31][19] ),
    .B2(net1384),
    .X(_06549_));
 sky130_fd_sc_hd__a21o_1 _11637_ (.A1(net1442),
    .A2(_06549_),
    .B1(net1466),
    .X(_06550_));
 sky130_fd_sc_hd__a21o_1 _11638_ (.A1(net1432),
    .A2(_06548_),
    .B1(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__a22o_1 _11639_ (.A1(net1680),
    .A2(\core.registers[22][19] ),
    .B1(\core.registers[23][19] ),
    .B2(net1385),
    .X(_06552_));
 sky130_fd_sc_hd__a22o_1 _11640_ (.A1(net1681),
    .A2(\core.registers[18][19] ),
    .B1(\core.registers[19][19] ),
    .B2(net1385),
    .X(_06553_));
 sky130_fd_sc_hd__mux2_1 _11641_ (.A0(_06552_),
    .A1(_06553_),
    .S(net1432),
    .X(_06554_));
 sky130_fd_sc_hd__mux4_1 _11642_ (.A0(\core.registers[16][19] ),
    .A1(\core.registers[17][19] ),
    .A2(\core.registers[20][19] ),
    .A3(\core.registers[21][19] ),
    .S0(net1386),
    .S1(net1442),
    .X(_06555_));
 sky130_fd_sc_hd__a31o_1 _11643_ (.A1(net1484),
    .A2(net1465),
    .A3(_06555_),
    .B1(net1460),
    .X(_06556_));
 sky130_fd_sc_hd__a31o_1 _11644_ (.A1(net1484),
    .A2(net1481),
    .A3(_06554_),
    .B1(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__a31o_1 _11645_ (.A1(net1489),
    .A2(_06547_),
    .A3(_06551_),
    .B1(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__nand2_2 _11646_ (.A(_06543_),
    .B(_06558_),
    .Y(_06559_));
 sky130_fd_sc_hd__o2bb2a_2 _11647_ (.A1_N(net1068),
    .A2_N(net1123),
    .B1(_06559_),
    .B2(_04663_),
    .X(_06560_));
 sky130_fd_sc_hd__inv_2 _11648_ (.A(_06560_),
    .Y(_06561_));
 sky130_fd_sc_hd__mux2_4 _11649_ (.A0(net460),
    .A1(_06561_),
    .S(net1278),
    .X(_06562_));
 sky130_fd_sc_hd__and2_2 _11650_ (.A(_06528_),
    .B(_06562_),
    .X(_06563_));
 sky130_fd_sc_hd__or2_1 _11651_ (.A(_06528_),
    .B(_06562_),
    .X(_06564_));
 sky130_fd_sc_hd__and2b_4 _11652_ (.A_N(_06563_),
    .B(_06564_),
    .X(_06565_));
 sky130_fd_sc_hd__or2_1 _11653_ (.A(\core.registers[1][18] ),
    .B(net1497),
    .X(_06566_));
 sky130_fd_sc_hd__or2_1 _11654_ (.A(\core.registers[6][18] ),
    .B(net1526),
    .X(_06567_));
 sky130_fd_sc_hd__or2_1 _11655_ (.A(\core.registers[17][18] ),
    .B(net1496),
    .X(_06568_));
 sky130_fd_sc_hd__or2_1 _11656_ (.A(\core.registers[28][18] ),
    .B(net1524),
    .X(_06569_));
 sky130_fd_sc_hd__o211a_1 _11657_ (.A1(\core.registers[29][18] ),
    .A2(net1496),
    .B1(_06569_),
    .C1(net1737),
    .X(_06570_));
 sky130_fd_sc_hd__a31o_1 _11658_ (.A1(net1841),
    .A2(net1722),
    .A3(\core.registers[30][18] ),
    .B1(net1749),
    .X(_06571_));
 sky130_fd_sc_hd__a31o_1 _11659_ (.A1(net1841),
    .A2(\core.registers[31][18] ),
    .A3(net1523),
    .B1(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__mux2_1 _11660_ (.A0(\core.registers[8][18] ),
    .A1(\core.registers[9][18] ),
    .S(net1523),
    .X(_06573_));
 sky130_fd_sc_hd__mux2_1 _11661_ (.A0(\core.registers[10][18] ),
    .A1(\core.registers[11][18] ),
    .S(net1527),
    .X(_06574_));
 sky130_fd_sc_hd__mux2_1 _11662_ (.A0(\core.registers[24][18] ),
    .A1(\core.registers[25][18] ),
    .S(net1525),
    .X(_06575_));
 sky130_fd_sc_hd__a221o_1 _11663_ (.A1(net1722),
    .A2(\core.registers[26][18] ),
    .B1(\core.registers[27][18] ),
    .B2(net1524),
    .C1(net1737),
    .X(_06576_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(\core.registers[12][18] ),
    .A1(\core.registers[13][18] ),
    .S(net1527),
    .X(_06577_));
 sky130_fd_sc_hd__mux2_1 _11665_ (.A0(\core.registers[14][18] ),
    .A1(\core.registers[15][18] ),
    .S(net1527),
    .X(_06578_));
 sky130_fd_sc_hd__mux2_1 _11666_ (.A0(_06577_),
    .A1(_06578_),
    .S(net1617),
    .X(_06579_));
 sky130_fd_sc_hd__o221a_1 _11667_ (.A1(_06570_),
    .A2(_06572_),
    .B1(_06579_),
    .B2(net1830),
    .C1(net1833),
    .X(_06580_));
 sky130_fd_sc_hd__mux2_1 _11668_ (.A0(_06573_),
    .A1(_06574_),
    .S(net1617),
    .X(_06581_));
 sky130_fd_sc_hd__o21a_1 _11669_ (.A1(net1841),
    .A2(_06575_),
    .B1(_06576_),
    .X(_06582_));
 sky130_fd_sc_hd__mux2_1 _11670_ (.A0(_06581_),
    .A1(_06582_),
    .S(net1830),
    .X(_06583_));
 sky130_fd_sc_hd__a211o_1 _11671_ (.A1(net1745),
    .A2(_06583_),
    .B1(_06580_),
    .C1(net1632),
    .X(_06584_));
 sky130_fd_sc_hd__o211a_1 _11672_ (.A1(net1722),
    .A2(\core.registers[7][18] ),
    .B1(net1617),
    .C1(_06567_),
    .X(_06585_));
 sky130_fd_sc_hd__mux2_1 _11673_ (.A0(\core.registers[4][18] ),
    .A1(\core.registers[5][18] ),
    .S(net1526),
    .X(_06586_));
 sky130_fd_sc_hd__a211o_1 _11674_ (.A1(net1603),
    .A2(_06586_),
    .B1(_06585_),
    .C1(net1577),
    .X(_06587_));
 sky130_fd_sc_hd__o211a_1 _11675_ (.A1(\core.registers[0][18] ),
    .A2(net1532),
    .B1(_06566_),
    .C1(net1604),
    .X(_06588_));
 sky130_fd_sc_hd__mux2_1 _11676_ (.A0(\core.registers[2][18] ),
    .A1(\core.registers[3][18] ),
    .S(net1532),
    .X(_06589_));
 sky130_fd_sc_hd__a211o_1 _11677_ (.A1(net1618),
    .A2(_06589_),
    .B1(_06588_),
    .C1(net1588),
    .X(_06590_));
 sky130_fd_sc_hd__o211a_1 _11678_ (.A1(\core.registers[16][18] ),
    .A2(net1526),
    .B1(_06568_),
    .C1(net1603),
    .X(_06591_));
 sky130_fd_sc_hd__mux2_1 _11679_ (.A0(\core.registers[18][18] ),
    .A1(\core.registers[19][18] ),
    .S(net1525),
    .X(_06592_));
 sky130_fd_sc_hd__a211o_1 _11680_ (.A1(net1618),
    .A2(_06592_),
    .B1(_06591_),
    .C1(net1588),
    .X(_06593_));
 sky130_fd_sc_hd__mux2_1 _11681_ (.A0(\core.registers[22][18] ),
    .A1(\core.registers[23][18] ),
    .S(net1526),
    .X(_06594_));
 sky130_fd_sc_hd__mux2_1 _11682_ (.A0(\core.registers[20][18] ),
    .A1(\core.registers[21][18] ),
    .S(net1526),
    .X(_06595_));
 sky130_fd_sc_hd__mux2_1 _11683_ (.A0(_06594_),
    .A1(_06595_),
    .S(net1603),
    .X(_06596_));
 sky130_fd_sc_hd__o211a_1 _11684_ (.A1(net1577),
    .A2(_06596_),
    .B1(_06593_),
    .C1(net1572),
    .X(_06597_));
 sky130_fd_sc_hd__a311o_1 _11685_ (.A1(net1568),
    .A2(_06587_),
    .A3(_06590_),
    .B1(_06597_),
    .C1(net1636),
    .X(_06598_));
 sky130_fd_sc_hd__a21o_1 _11686_ (.A1(_06584_),
    .A2(_06598_),
    .B1(net1158),
    .X(_06599_));
 sky130_fd_sc_hd__a21o_4 _11687_ (.A1(net1234),
    .A2(_05377_),
    .B1(net1236),
    .X(_06600_));
 sky130_fd_sc_hd__a22o_1 _11688_ (.A1(\core.pipe1_resultRegister[18] ),
    .A2(net1240),
    .B1(_04520_),
    .B2(\core.pipe1_csrData[18] ),
    .X(_06601_));
 sky130_fd_sc_hd__a21o_1 _11689_ (.A1(net1191),
    .A2(_06600_),
    .B1(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__o211ai_2 _11690_ (.A1(net1154),
    .A2(net1119),
    .B1(_06599_),
    .C1(net1264),
    .Y(_06603_));
 sky130_fd_sc_hd__o21ai_1 _11691_ (.A1(net1192),
    .A2(_06603_),
    .B1(net1161),
    .Y(_06604_));
 sky130_fd_sc_hd__o21a_1 _11692_ (.A1(\core.pipe0_currentInstruction[18] ),
    .A2(net1278),
    .B1(_06604_),
    .X(_06605_));
 sky130_fd_sc_hd__or2_1 _11693_ (.A(\core.registers[13][18] ),
    .B(net1375),
    .X(_06606_));
 sky130_fd_sc_hd__o211a_1 _11694_ (.A1(\core.registers[12][18] ),
    .A2(net1394),
    .B1(_06606_),
    .C1(net1447),
    .X(_06607_));
 sky130_fd_sc_hd__a31o_1 _11695_ (.A1(\core.registers[9][18] ),
    .A2(net1435),
    .A3(net1394),
    .B1(net1482),
    .X(_06608_));
 sky130_fd_sc_hd__a311o_1 _11696_ (.A1(\core.registers[8][18] ),
    .A2(net1435),
    .A3(net1374),
    .B1(_06607_),
    .C1(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__a22o_1 _11697_ (.A1(net1684),
    .A2(\core.registers[10][18] ),
    .B1(\core.registers[11][18] ),
    .B2(net1398),
    .X(_06610_));
 sky130_fd_sc_hd__a22o_1 _11698_ (.A1(net1684),
    .A2(\core.registers[14][18] ),
    .B1(\core.registers[15][18] ),
    .B2(net1398),
    .X(_06611_));
 sky130_fd_sc_hd__a21o_1 _11699_ (.A1(net1447),
    .A2(_06611_),
    .B1(net1469),
    .X(_06612_));
 sky130_fd_sc_hd__a21o_1 _11700_ (.A1(net1435),
    .A2(_06610_),
    .B1(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__a22o_1 _11701_ (.A1(net1685),
    .A2(\core.registers[6][18] ),
    .B1(\core.registers[7][18] ),
    .B2(net1397),
    .X(_06614_));
 sky130_fd_sc_hd__a22o_1 _11702_ (.A1(net1685),
    .A2(\core.registers[2][18] ),
    .B1(\core.registers[3][18] ),
    .B2(net1402),
    .X(_06615_));
 sky130_fd_sc_hd__mux2_1 _11703_ (.A0(_06614_),
    .A1(_06615_),
    .S(net1435),
    .X(_06616_));
 sky130_fd_sc_hd__mux4_1 _11704_ (.A0(\core.registers[0][18] ),
    .A1(\core.registers[1][18] ),
    .A2(\core.registers[4][18] ),
    .A3(\core.registers[5][18] ),
    .S0(net1396),
    .S1(net1447),
    .X(_06617_));
 sky130_fd_sc_hd__a31o_1 _11705_ (.A1(net1486),
    .A2(net1469),
    .A3(_06617_),
    .B1(net1464),
    .X(_06618_));
 sky130_fd_sc_hd__a31o_1 _11706_ (.A1(net1486),
    .A2(net1481),
    .A3(_06616_),
    .B1(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__a31o_1 _11707_ (.A1(net1490),
    .A2(_06609_),
    .A3(_06613_),
    .B1(_06619_),
    .X(_06620_));
 sky130_fd_sc_hd__or2_1 _11708_ (.A(\core.registers[29][18] ),
    .B(net1374),
    .X(_06621_));
 sky130_fd_sc_hd__o211a_1 _11709_ (.A1(\core.registers[28][18] ),
    .A2(net1395),
    .B1(_06621_),
    .C1(net1447),
    .X(_06622_));
 sky130_fd_sc_hd__a31o_1 _11710_ (.A1(\core.registers[25][18] ),
    .A2(net1435),
    .A3(net1396),
    .B1(net1481),
    .X(_06623_));
 sky130_fd_sc_hd__a311o_1 _11711_ (.A1(\core.registers[24][18] ),
    .A2(net1435),
    .A3(net1374),
    .B1(_06622_),
    .C1(_06623_),
    .X(_06624_));
 sky130_fd_sc_hd__a22o_1 _11712_ (.A1(net1684),
    .A2(\core.registers[26][18] ),
    .B1(\core.registers[27][18] ),
    .B2(net1395),
    .X(_06625_));
 sky130_fd_sc_hd__a22o_1 _11713_ (.A1(net1684),
    .A2(\core.registers[30][18] ),
    .B1(\core.registers[31][18] ),
    .B2(net1395),
    .X(_06626_));
 sky130_fd_sc_hd__a21o_1 _11714_ (.A1(net1447),
    .A2(_06626_),
    .B1(net1469),
    .X(_06627_));
 sky130_fd_sc_hd__a21o_1 _11715_ (.A1(net1435),
    .A2(_06625_),
    .B1(_06627_),
    .X(_06628_));
 sky130_fd_sc_hd__a22o_1 _11716_ (.A1(net1685),
    .A2(\core.registers[22][18] ),
    .B1(\core.registers[23][18] ),
    .B2(net1397),
    .X(_06629_));
 sky130_fd_sc_hd__a22o_1 _11717_ (.A1(net1685),
    .A2(\core.registers[18][18] ),
    .B1(\core.registers[19][18] ),
    .B2(net1396),
    .X(_06630_));
 sky130_fd_sc_hd__mux2_1 _11718_ (.A0(_06629_),
    .A1(_06630_),
    .S(net1435),
    .X(_06631_));
 sky130_fd_sc_hd__mux4_1 _11719_ (.A0(\core.registers[16][18] ),
    .A1(\core.registers[17][18] ),
    .A2(\core.registers[20][18] ),
    .A3(\core.registers[21][18] ),
    .S0(net1397),
    .S1(net1447),
    .X(_06632_));
 sky130_fd_sc_hd__a31o_1 _11720_ (.A1(net1486),
    .A2(net1469),
    .A3(_06632_),
    .B1(net1461),
    .X(_06633_));
 sky130_fd_sc_hd__a31o_1 _11721_ (.A1(net1486),
    .A2(net1481),
    .A3(_06631_),
    .B1(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__a31o_1 _11722_ (.A1(net1490),
    .A2(_06624_),
    .A3(_06628_),
    .B1(_06634_),
    .X(_06635_));
 sky130_fd_sc_hd__nand2_2 _11723_ (.A(_06620_),
    .B(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__o2bb2a_2 _11724_ (.A1_N(net1069),
    .A2_N(net1119),
    .B1(_06636_),
    .B2(_04663_),
    .X(_06637_));
 sky130_fd_sc_hd__inv_2 _11725_ (.A(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__mux2_4 _11726_ (.A0(net459),
    .A1(_06638_),
    .S(net1279),
    .X(_06639_));
 sky130_fd_sc_hd__or2_2 _11727_ (.A(_06605_),
    .B(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__clkinv_2 _11728_ (.A(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__and2_4 _11729_ (.A(_06605_),
    .B(_06639_),
    .X(_06642_));
 sky130_fd_sc_hd__nor2_8 _11730_ (.A(_06641_),
    .B(_06642_),
    .Y(_06643_));
 sky130_fd_sc_hd__or4_1 _11731_ (.A(_06410_),
    .B(_06488_),
    .C(_06565_),
    .D(_06643_),
    .X(_06644_));
 sky130_fd_sc_hd__a21o_2 _11732_ (.A1(_06323_),
    .A2(_06330_),
    .B1(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__nand2b_1 _11733_ (.A_N(_06605_),
    .B(_06639_),
    .Y(_06646_));
 sky130_fd_sc_hd__nand2b_1 _11734_ (.A_N(_06370_),
    .B(_06406_),
    .Y(_06647_));
 sky130_fd_sc_hd__nand2b_2 _11735_ (.A_N(_06450_),
    .B(_06484_),
    .Y(_06648_));
 sky130_fd_sc_hd__o21ai_1 _11736_ (.A1(_06410_),
    .A2(_06648_),
    .B1(_06647_),
    .Y(_06649_));
 sky130_fd_sc_hd__nand2b_1 _11737_ (.A_N(_06528_),
    .B(_06562_),
    .Y(_06650_));
 sky130_fd_sc_hd__or3b_1 _11738_ (.A(_06565_),
    .B(_06643_),
    .C_N(_06649_),
    .X(_06651_));
 sky130_fd_sc_hd__o211a_2 _11739_ (.A1(_06565_),
    .A2(_06646_),
    .B1(_06650_),
    .C1(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__or2_4 _11740_ (.A(_04897_),
    .B(_04927_),
    .X(_06653_));
 sky130_fd_sc_hd__clkinv_2 _11741_ (.A(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__and2_4 _11742_ (.A(_04897_),
    .B(_04927_),
    .X(_06655_));
 sky130_fd_sc_hd__nor2_8 _11743_ (.A(_06654_),
    .B(_06655_),
    .Y(_06656_));
 sky130_fd_sc_hd__a21o_1 _11744_ (.A1(_06645_),
    .A2(_06652_),
    .B1(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__a211o_1 _11745_ (.A1(_06645_),
    .A2(_06652_),
    .B1(_06656_),
    .C1(_04854_),
    .X(_06658_));
 sky130_fd_sc_hd__a21o_1 _11746_ (.A1(_04931_),
    .A2(_06658_),
    .B1(_04777_),
    .X(_06659_));
 sky130_fd_sc_hd__and2b_2 _11747_ (.A_N(_04772_),
    .B(_06659_),
    .X(_06660_));
 sky130_fd_sc_hd__xnor2_4 _11748_ (.A(_04697_),
    .B(_06660_),
    .Y(_06661_));
 sky130_fd_sc_hd__a21o_1 _11749_ (.A1(_06323_),
    .A2(_06330_),
    .B1(_06488_),
    .X(_06662_));
 sky130_fd_sc_hd__a21o_1 _11750_ (.A1(_06648_),
    .A2(_06662_),
    .B1(_06410_),
    .X(_06663_));
 sky130_fd_sc_hd__o21ba_2 _11751_ (.A1(_06410_),
    .A2(_06662_),
    .B1_N(_06649_),
    .X(_06664_));
 sky130_fd_sc_hd__xor2_2 _11752_ (.A(_06643_),
    .B(_06664_),
    .X(_06665_));
 sky130_fd_sc_hd__o211a_2 _11753_ (.A1(_06316_),
    .A2(_06318_),
    .B1(_05026_),
    .C1(_05558_),
    .X(_06666_));
 sky130_fd_sc_hd__nor2_1 _11754_ (.A(_06325_),
    .B(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__a21boi_4 _11755_ (.A1(_05111_),
    .A2(_06666_),
    .B1_N(_06326_),
    .Y(_06668_));
 sky130_fd_sc_hd__o21a_1 _11756_ (.A1(_05280_),
    .A2(_06668_),
    .B1(_06327_),
    .X(_06669_));
 sky130_fd_sc_hd__xnor2_2 _11757_ (.A(_05191_),
    .B(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__nand3_1 _11758_ (.A(_04854_),
    .B(_04928_),
    .C(_06657_),
    .Y(_06671_));
 sky130_fd_sc_hd__a21o_1 _11759_ (.A1(_04928_),
    .A2(_06657_),
    .B1(_04854_),
    .X(_06672_));
 sky130_fd_sc_hd__a211oi_1 _11760_ (.A1(_06671_),
    .A2(_06672_),
    .B1(_06665_),
    .C1(_06670_),
    .Y(_06673_));
 sky130_fd_sc_hd__or3b_1 _11761_ (.A(_04776_),
    .B(_04930_),
    .C_N(_06658_),
    .X(_06674_));
 sky130_fd_sc_hd__o21bai_2 _11762_ (.A1(_06316_),
    .A2(_06317_),
    .B1_N(_05551_),
    .Y(_06675_));
 sky130_fd_sc_hd__a21o_1 _11763_ (.A1(_05555_),
    .A2(_06675_),
    .B1(_05455_),
    .X(_06676_));
 sky130_fd_sc_hd__nand3_1 _11764_ (.A(_05368_),
    .B(_05554_),
    .C(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__a21o_1 _11765_ (.A1(_05554_),
    .A2(_06676_),
    .B1(_05368_),
    .X(_06678_));
 sky130_fd_sc_hd__nand3_1 _11766_ (.A(_05455_),
    .B(_05555_),
    .C(_06675_),
    .Y(_06679_));
 sky130_fd_sc_hd__a211o_1 _11767_ (.A1(_05552_),
    .A2(_06316_),
    .B1(_06321_),
    .C1(_05026_),
    .X(_06680_));
 sky130_fd_sc_hd__and2b_1 _11768_ (.A_N(_06666_),
    .B(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__a31o_1 _11769_ (.A1(_05799_),
    .A2(_05883_),
    .A3(_06231_),
    .B1(_06236_),
    .X(_06682_));
 sky130_fd_sc_hd__a21bo_1 _11770_ (.A1(_05714_),
    .A2(_06682_),
    .B1_N(_05716_),
    .X(_06683_));
 sky130_fd_sc_hd__xnor2_2 _11771_ (.A(_05633_),
    .B(_06683_),
    .Y(_06684_));
 sky130_fd_sc_hd__or3b_1 _11772_ (.A(_06316_),
    .B(_06317_),
    .C_N(_05551_),
    .X(_06685_));
 sky130_fd_sc_hd__and2_1 _11773_ (.A(_06675_),
    .B(_06685_),
    .X(_06686_));
 sky130_fd_sc_hd__xnor2_1 _11774_ (.A(_06237_),
    .B(_06314_),
    .Y(_06687_));
 sky130_fd_sc_hd__xnor2_1 _11775_ (.A(_05713_),
    .B(_06682_),
    .Y(_06688_));
 sky130_fd_sc_hd__nand2_1 _11776_ (.A(_05798_),
    .B(_06233_),
    .Y(_06689_));
 sky130_fd_sc_hd__a21o_1 _11777_ (.A1(_05883_),
    .A2(_06231_),
    .B1(_06689_),
    .X(_06690_));
 sky130_fd_sc_hd__and3b_1 _11778_ (.A_N(_06232_),
    .B(_06234_),
    .C(_06690_),
    .X(_06691_));
 sky130_fd_sc_hd__xor2_1 _11779_ (.A(_05883_),
    .B(_06231_),
    .X(_06692_));
 sky130_fd_sc_hd__xnor2_1 _11780_ (.A(_05968_),
    .B(_06230_),
    .Y(_06693_));
 sky130_fd_sc_hd__xnor2_1 _11781_ (.A(_06053_),
    .B(_06229_),
    .Y(_06694_));
 sky130_fd_sc_hd__nand2_8 _11782_ (.A(net932),
    .B(_06227_),
    .Y(_06695_));
 sky130_fd_sc_hd__or2_2 _11783_ (.A(net932),
    .B(_06227_),
    .X(_06696_));
 sky130_fd_sc_hd__and2_4 _11784_ (.A(_06695_),
    .B(_06696_),
    .X(_06697_));
 sky130_fd_sc_hd__nand2_1 _11785_ (.A(_06695_),
    .B(_06696_),
    .Y(_06698_));
 sky130_fd_sc_hd__and4_1 _11786_ (.A(_06137_),
    .B(_06693_),
    .C(_06694_),
    .D(net831),
    .X(_06699_));
 sky130_fd_sc_hd__or4b_1 _11787_ (.A(_06688_),
    .B(_06691_),
    .C(_06692_),
    .D_N(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__or3_4 _11788_ (.A(_06684_),
    .B(_06687_),
    .C(_06700_),
    .X(_06701_));
 sky130_fd_sc_hd__a2111o_1 _11789_ (.A1(_06676_),
    .A2(_06679_),
    .B1(_06681_),
    .C1(_06686_),
    .D1(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__xnor2_1 _11790_ (.A(_05111_),
    .B(_06667_),
    .Y(_06703_));
 sky130_fd_sc_hd__nand3_1 _11791_ (.A(_06323_),
    .B(_06330_),
    .C(_06488_),
    .Y(_06704_));
 sky130_fd_sc_hd__and2_1 _11792_ (.A(_06662_),
    .B(_06704_),
    .X(_06705_));
 sky130_fd_sc_hd__a2111o_2 _11793_ (.A1(_06677_),
    .A2(_06678_),
    .B1(_06702_),
    .C1(_06703_),
    .D1(_06705_),
    .X(_06706_));
 sky130_fd_sc_hd__nand3_1 _11794_ (.A(_06410_),
    .B(_06648_),
    .C(_06662_),
    .Y(_06707_));
 sky130_fd_sc_hd__nand3_1 _11795_ (.A(_06645_),
    .B(_06652_),
    .C(_06656_),
    .Y(_06708_));
 sky130_fd_sc_hd__xnor2_2 _11796_ (.A(_05279_),
    .B(_06668_),
    .Y(_06709_));
 sky130_fd_sc_hd__a221o_1 _11797_ (.A1(_06663_),
    .A2(_06707_),
    .B1(_06708_),
    .B2(_06657_),
    .C1(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__a211o_1 _11798_ (.A1(_06659_),
    .A2(_06674_),
    .B1(_06706_),
    .C1(_06710_),
    .X(_06711_));
 sky130_fd_sc_hd__nand2b_1 _11799_ (.A_N(_04640_),
    .B(_04693_),
    .Y(_06712_));
 sky130_fd_sc_hd__or4_1 _11800_ (.A(_04697_),
    .B(_04777_),
    .C(_04854_),
    .D(_06656_),
    .X(_06713_));
 sky130_fd_sc_hd__a21o_1 _11801_ (.A1(_06645_),
    .A2(_06652_),
    .B1(_06713_),
    .X(_06714_));
 sky130_fd_sc_hd__a21oi_1 _11802_ (.A1(_04776_),
    .A2(_04930_),
    .B1(_04772_),
    .Y(_06715_));
 sky130_fd_sc_hd__o21a_1 _11803_ (.A1(_04697_),
    .A2(_06715_),
    .B1(_06712_),
    .X(_06716_));
 sky130_fd_sc_hd__nand2_2 _11804_ (.A(_06714_),
    .B(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__a22o_1 _11805_ (.A1(\core.pipe1_resultRegister[24] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[24] ),
    .X(_06718_));
 sky130_fd_sc_hd__a21o_4 _11806_ (.A1(net1234),
    .A2(_06142_),
    .B1(net2014),
    .X(_06719_));
 sky130_fd_sc_hd__a21o_4 _11807_ (.A1(net1188),
    .A2(_06719_),
    .B1(_06718_),
    .X(_06720_));
 sky130_fd_sc_hd__or2_1 _11808_ (.A(\core.registers[1][24] ),
    .B(net1494),
    .X(_06721_));
 sky130_fd_sc_hd__or2_1 _11809_ (.A(\core.registers[6][24] ),
    .B(net1518),
    .X(_06722_));
 sky130_fd_sc_hd__or2_1 _11810_ (.A(\core.registers[17][24] ),
    .B(net1494),
    .X(_06723_));
 sky130_fd_sc_hd__or2_1 _11811_ (.A(\core.registers[28][24] ),
    .B(net1505),
    .X(_06724_));
 sky130_fd_sc_hd__o211a_1 _11812_ (.A1(\core.registers[29][24] ),
    .A2(net1493),
    .B1(_06724_),
    .C1(net1735),
    .X(_06725_));
 sky130_fd_sc_hd__a31o_1 _11813_ (.A1(net1838),
    .A2(net1719),
    .A3(\core.registers[30][24] ),
    .B1(net1748),
    .X(_06726_));
 sky130_fd_sc_hd__a31o_1 _11814_ (.A1(net1838),
    .A2(\core.registers[31][24] ),
    .A3(net1505),
    .B1(_06726_),
    .X(_06727_));
 sky130_fd_sc_hd__mux2_1 _11815_ (.A0(\core.registers[8][24] ),
    .A1(\core.registers[9][24] ),
    .S(net1504),
    .X(_06728_));
 sky130_fd_sc_hd__mux2_1 _11816_ (.A0(\core.registers[10][24] ),
    .A1(\core.registers[11][24] ),
    .S(net1504),
    .X(_06729_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(\core.registers[24][24] ),
    .A1(\core.registers[25][24] ),
    .S(net1505),
    .X(_06730_));
 sky130_fd_sc_hd__a221o_1 _11818_ (.A1(net1719),
    .A2(\core.registers[26][24] ),
    .B1(\core.registers[27][24] ),
    .B2(net1508),
    .C1(net1735),
    .X(_06731_));
 sky130_fd_sc_hd__mux2_1 _11819_ (.A0(\core.registers[12][24] ),
    .A1(\core.registers[13][24] ),
    .S(net1504),
    .X(_06732_));
 sky130_fd_sc_hd__mux2_1 _11820_ (.A0(\core.registers[14][24] ),
    .A1(\core.registers[15][24] ),
    .S(net1504),
    .X(_06733_));
 sky130_fd_sc_hd__mux2_1 _11821_ (.A0(_06732_),
    .A1(_06733_),
    .S(net1611),
    .X(_06734_));
 sky130_fd_sc_hd__o221a_1 _11822_ (.A1(_06725_),
    .A2(_06727_),
    .B1(_06734_),
    .B2(net1823),
    .C1(net1832),
    .X(_06735_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(_06728_),
    .A1(_06729_),
    .S(net1611),
    .X(_06736_));
 sky130_fd_sc_hd__o21a_1 _11824_ (.A1(net1838),
    .A2(_06730_),
    .B1(_06731_),
    .X(_06737_));
 sky130_fd_sc_hd__mux2_1 _11825_ (.A0(_06736_),
    .A1(_06737_),
    .S(net1823),
    .X(_06738_));
 sky130_fd_sc_hd__a211o_4 _11826_ (.A1(net1744),
    .A2(_06738_),
    .B1(_06735_),
    .C1(net1631),
    .X(_06739_));
 sky130_fd_sc_hd__o211a_1 _11827_ (.A1(net1725),
    .A2(\core.registers[7][24] ),
    .B1(net1615),
    .C1(_06722_),
    .X(_06740_));
 sky130_fd_sc_hd__mux2_1 _11828_ (.A0(\core.registers[4][24] ),
    .A1(\core.registers[5][24] ),
    .S(net1518),
    .X(_06741_));
 sky130_fd_sc_hd__a211o_1 _11829_ (.A1(net1600),
    .A2(_06741_),
    .B1(_06740_),
    .C1(net1575),
    .X(_06742_));
 sky130_fd_sc_hd__o211a_1 _11830_ (.A1(\core.registers[0][24] ),
    .A2(net1519),
    .B1(_06721_),
    .C1(net1599),
    .X(_06743_));
 sky130_fd_sc_hd__mux2_1 _11831_ (.A0(\core.registers[2][24] ),
    .A1(\core.registers[3][24] ),
    .S(net1518),
    .X(_06744_));
 sky130_fd_sc_hd__a211o_1 _11832_ (.A1(net1615),
    .A2(_06744_),
    .B1(_06743_),
    .C1(net1587),
    .X(_06745_));
 sky130_fd_sc_hd__o211a_1 _11833_ (.A1(\core.registers[16][24] ),
    .A2(net1521),
    .B1(_06723_),
    .C1(net1601),
    .X(_06746_));
 sky130_fd_sc_hd__mux2_1 _11834_ (.A0(\core.registers[18][24] ),
    .A1(\core.registers[19][24] ),
    .S(net1521),
    .X(_06747_));
 sky130_fd_sc_hd__a211o_1 _11835_ (.A1(net1616),
    .A2(_06747_),
    .B1(_06746_),
    .C1(net1586),
    .X(_06748_));
 sky130_fd_sc_hd__mux2_1 _11836_ (.A0(\core.registers[22][24] ),
    .A1(\core.registers[23][24] ),
    .S(net1518),
    .X(_06749_));
 sky130_fd_sc_hd__mux2_1 _11837_ (.A0(\core.registers[20][24] ),
    .A1(\core.registers[21][24] ),
    .S(net1521),
    .X(_06750_));
 sky130_fd_sc_hd__mux2_1 _11838_ (.A0(_06749_),
    .A1(_06750_),
    .S(net1599),
    .X(_06751_));
 sky130_fd_sc_hd__o211a_1 _11839_ (.A1(net1575),
    .A2(_06751_),
    .B1(_06748_),
    .C1(net1571),
    .X(_06752_));
 sky130_fd_sc_hd__a311o_1 _11840_ (.A1(net1567),
    .A2(_06742_),
    .A3(_06745_),
    .B1(_06752_),
    .C1(net1635),
    .X(_06753_));
 sky130_fd_sc_hd__a21o_2 _11841_ (.A1(_06739_),
    .A2(_06753_),
    .B1(net1157),
    .X(_06754_));
 sky130_fd_sc_hd__o211ai_4 _11842_ (.A1(net1153),
    .A2(net1115),
    .B1(_06754_),
    .C1(net1263),
    .Y(_06755_));
 sky130_fd_sc_hd__o21a_1 _11843_ (.A1(net1192),
    .A2(_06755_),
    .B1(net1161),
    .X(_06756_));
 sky130_fd_sc_hd__a21oi_2 _11844_ (.A1(_04415_),
    .A2(net1285),
    .B1(_06756_),
    .Y(_06757_));
 sky130_fd_sc_hd__o22a_1 _11845_ (.A1(net1682),
    .A2(\core.registers[23][24] ),
    .B1(net1391),
    .B2(\core.registers[22][24] ),
    .X(_06758_));
 sky130_fd_sc_hd__or3_1 _11846_ (.A(net1683),
    .B(\core.registers[19][24] ),
    .C(net1446),
    .X(_06759_));
 sky130_fd_sc_hd__o221a_1 _11847_ (.A1(\core.registers[18][24] ),
    .A2(net1331),
    .B1(_06758_),
    .B2(net1434),
    .C1(_06759_),
    .X(_06760_));
 sky130_fd_sc_hd__mux4_1 _11848_ (.A0(\core.registers[16][24] ),
    .A1(\core.registers[17][24] ),
    .A2(\core.registers[20][24] ),
    .A3(\core.registers[21][24] ),
    .S0(net1393),
    .S1(net1446),
    .X(_06761_));
 sky130_fd_sc_hd__mux2_1 _11849_ (.A0(_06760_),
    .A1(_06761_),
    .S(net1467),
    .X(_06762_));
 sky130_fd_sc_hd__o22a_1 _11850_ (.A1(net1682),
    .A2(\core.registers[7][24] ),
    .B1(net1391),
    .B2(\core.registers[6][24] ),
    .X(_06763_));
 sky130_fd_sc_hd__or3_1 _11851_ (.A(net1682),
    .B(\core.registers[3][24] ),
    .C(net1445),
    .X(_06764_));
 sky130_fd_sc_hd__o221a_1 _11852_ (.A1(\core.registers[2][24] ),
    .A2(net1331),
    .B1(_06763_),
    .B2(net1437),
    .C1(_06764_),
    .X(_06765_));
 sky130_fd_sc_hd__mux4_1 _11853_ (.A0(\core.registers[0][24] ),
    .A1(\core.registers[1][24] ),
    .A2(\core.registers[4][24] ),
    .A3(\core.registers[5][24] ),
    .S0(net1391),
    .S1(net1446),
    .X(_06766_));
 sky130_fd_sc_hd__mux2_1 _11854_ (.A0(_06765_),
    .A1(_06766_),
    .S(net1468),
    .X(_06767_));
 sky130_fd_sc_hd__mux2_1 _11855_ (.A0(_06762_),
    .A1(_06767_),
    .S(net1460),
    .X(_06768_));
 sky130_fd_sc_hd__mux2_1 _11856_ (.A0(\core.registers[14][24] ),
    .A1(\core.registers[15][24] ),
    .S(net1379),
    .X(_06769_));
 sky130_fd_sc_hd__mux2_1 _11857_ (.A0(\core.registers[12][24] ),
    .A1(\core.registers[13][24] ),
    .S(net1379),
    .X(_06770_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(_06769_),
    .A1(_06770_),
    .S(net1465),
    .X(_06771_));
 sky130_fd_sc_hd__mux2_1 _11859_ (.A0(\core.registers[28][24] ),
    .A1(\core.registers[29][24] ),
    .S(net1380),
    .X(_06772_));
 sky130_fd_sc_hd__a221o_1 _11860_ (.A1(net1678),
    .A2(\core.registers[30][24] ),
    .B1(\core.registers[31][24] ),
    .B2(net1387),
    .C1(net1704),
    .X(_06773_));
 sky130_fd_sc_hd__o21ai_1 _11861_ (.A1(net1868),
    .A2(_06772_),
    .B1(_06773_),
    .Y(_06774_));
 sky130_fd_sc_hd__nand2_1 _11862_ (.A(net1853),
    .B(_06774_),
    .Y(_06775_));
 sky130_fd_sc_hd__o211a_1 _11863_ (.A1(net1853),
    .A2(_06771_),
    .B1(_06775_),
    .C1(net1862),
    .X(_06776_));
 sky130_fd_sc_hd__a221o_1 _11864_ (.A1(net1678),
    .A2(\core.registers[26][24] ),
    .B1(\core.registers[27][24] ),
    .B2(net1380),
    .C1(net1704),
    .X(_06777_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(\core.registers[24][24] ),
    .A1(\core.registers[25][24] ),
    .S(net1380),
    .X(_06778_));
 sky130_fd_sc_hd__o21ai_1 _11866_ (.A1(net1868),
    .A2(_06778_),
    .B1(_06777_),
    .Y(_06779_));
 sky130_fd_sc_hd__o21a_1 _11867_ (.A1(\core.registers[8][24] ),
    .A2(net1379),
    .B1(net1704),
    .X(_06780_));
 sky130_fd_sc_hd__o21ai_1 _11868_ (.A1(\core.registers[9][24] ),
    .A2(net1373),
    .B1(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__a22o_1 _11869_ (.A1(net1678),
    .A2(\core.registers[10][24] ),
    .B1(\core.registers[11][24] ),
    .B2(net1379),
    .X(_06782_));
 sky130_fd_sc_hd__a21oi_1 _11870_ (.A1(net1868),
    .A2(_06782_),
    .B1(net1853),
    .Y(_06783_));
 sky130_fd_sc_hd__a221o_1 _11871_ (.A1(net1853),
    .A2(_06779_),
    .B1(_06781_),
    .B2(_06783_),
    .C1(net1862),
    .X(_06784_));
 sky130_fd_sc_hd__or3b_4 _11872_ (.A(net1484),
    .B(_06776_),
    .C_N(_06784_),
    .X(_06785_));
 sky130_fd_sc_hd__o21a_1 _11873_ (.A1(net1490),
    .A2(_06768_),
    .B1(_06785_),
    .X(_06786_));
 sky130_fd_sc_hd__a22o_2 _11874_ (.A1(net1068),
    .A2(net1114),
    .B1(_06786_),
    .B2(net1065),
    .X(_06787_));
 sky130_fd_sc_hd__mux2_8 _11875_ (.A0(net466),
    .A1(_06787_),
    .S(net1276),
    .X(_06788_));
 sky130_fd_sc_hd__nor2_2 _11876_ (.A(_06757_),
    .B(_06788_),
    .Y(_06789_));
 sky130_fd_sc_hd__and2_2 _11877_ (.A(_06757_),
    .B(_06788_),
    .X(_06790_));
 sky130_fd_sc_hd__nor2_4 _11878_ (.A(_06789_),
    .B(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__inv_2 _11879_ (.A(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__xnor2_2 _11880_ (.A(_06717_),
    .B(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__o21ai_1 _11881_ (.A1(_06643_),
    .A2(_06664_),
    .B1(_06646_),
    .Y(_06794_));
 sky130_fd_sc_hd__xnor2_1 _11882_ (.A(_06565_),
    .B(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__and4bb_2 _11883_ (.A_N(_06795_),
    .B_N(_06711_),
    .C(_06673_),
    .D(_06793_),
    .X(_06796_));
 sky130_fd_sc_hd__a22o_1 _11884_ (.A1(\core.pipe1_resultRegister[25] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[25] ),
    .X(_06797_));
 sky130_fd_sc_hd__a21o_4 _11885_ (.A1(net1234),
    .A2(_05470_),
    .B1(net2014),
    .X(_06798_));
 sky130_fd_sc_hd__a21o_1 _11886_ (.A1(net1188),
    .A2(_06798_),
    .B1(_06797_),
    .X(_06799_));
 sky130_fd_sc_hd__mux2_1 _11887_ (.A0(\core.registers[8][25] ),
    .A1(\core.registers[9][25] ),
    .S(net1505),
    .X(_06800_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(\core.registers[10][25] ),
    .A1(\core.registers[11][25] ),
    .S(net1505),
    .X(_06801_));
 sky130_fd_sc_hd__mux2_1 _11889_ (.A0(\core.registers[24][25] ),
    .A1(\core.registers[25][25] ),
    .S(net1509),
    .X(_06802_));
 sky130_fd_sc_hd__a221o_1 _11890_ (.A1(net1720),
    .A2(\core.registers[26][25] ),
    .B1(\core.registers[27][25] ),
    .B2(net1509),
    .C1(net1735),
    .X(_06803_));
 sky130_fd_sc_hd__or2_1 _11891_ (.A(\core.registers[28][25] ),
    .B(net1505),
    .X(_06804_));
 sky130_fd_sc_hd__o211a_1 _11892_ (.A1(\core.registers[29][25] ),
    .A2(net1493),
    .B1(_06804_),
    .C1(net1735),
    .X(_06805_));
 sky130_fd_sc_hd__a31o_1 _11893_ (.A1(net1838),
    .A2(net1719),
    .A3(\core.registers[30][25] ),
    .B1(net1748),
    .X(_06806_));
 sky130_fd_sc_hd__a31o_1 _11894_ (.A1(net1839),
    .A2(\core.registers[31][25] ),
    .A3(net1505),
    .B1(_06806_),
    .X(_06807_));
 sky130_fd_sc_hd__or2_1 _11895_ (.A(\core.registers[1][25] ),
    .B(net1495),
    .X(_06808_));
 sky130_fd_sc_hd__or2_1 _11896_ (.A(\core.registers[6][25] ),
    .B(net1511),
    .X(_06809_));
 sky130_fd_sc_hd__or2_1 _11897_ (.A(\core.registers[17][25] ),
    .B(net1493),
    .X(_06810_));
 sky130_fd_sc_hd__mux2_1 _11898_ (.A0(\core.registers[12][25] ),
    .A1(\core.registers[13][25] ),
    .S(net1504),
    .X(_06811_));
 sky130_fd_sc_hd__mux2_1 _11899_ (.A0(\core.registers[14][25] ),
    .A1(\core.registers[15][25] ),
    .S(net1504),
    .X(_06812_));
 sky130_fd_sc_hd__mux2_1 _11900_ (.A0(_06811_),
    .A1(_06812_),
    .S(net1611),
    .X(_06813_));
 sky130_fd_sc_hd__o221a_1 _11901_ (.A1(_06805_),
    .A2(_06807_),
    .B1(_06813_),
    .B2(net1823),
    .C1(net1832),
    .X(_06814_));
 sky130_fd_sc_hd__mux2_1 _11902_ (.A0(_06800_),
    .A1(_06801_),
    .S(net1611),
    .X(_06815_));
 sky130_fd_sc_hd__o21a_1 _11903_ (.A1(net1838),
    .A2(_06802_),
    .B1(_06803_),
    .X(_06816_));
 sky130_fd_sc_hd__mux2_1 _11904_ (.A0(_06815_),
    .A1(_06816_),
    .S(net1823),
    .X(_06817_));
 sky130_fd_sc_hd__a211o_1 _11905_ (.A1(net1744),
    .A2(_06817_),
    .B1(_06814_),
    .C1(net1631),
    .X(_06818_));
 sky130_fd_sc_hd__o211a_1 _11906_ (.A1(net1720),
    .A2(\core.registers[7][25] ),
    .B1(net1613),
    .C1(_06809_),
    .X(_06819_));
 sky130_fd_sc_hd__mux2_1 _11907_ (.A0(\core.registers[4][25] ),
    .A1(\core.registers[5][25] ),
    .S(net1511),
    .X(_06820_));
 sky130_fd_sc_hd__a211o_1 _11908_ (.A1(net1597),
    .A2(_06820_),
    .B1(_06819_),
    .C1(net1576),
    .X(_06821_));
 sky130_fd_sc_hd__o211a_1 _11909_ (.A1(\core.registers[0][25] ),
    .A2(net1511),
    .B1(_06808_),
    .C1(net1597),
    .X(_06822_));
 sky130_fd_sc_hd__mux2_1 _11910_ (.A0(\core.registers[2][25] ),
    .A1(\core.registers[3][25] ),
    .S(net1511),
    .X(_06823_));
 sky130_fd_sc_hd__a211o_1 _11911_ (.A1(net1613),
    .A2(_06823_),
    .B1(_06822_),
    .C1(net1587),
    .X(_06824_));
 sky130_fd_sc_hd__o211a_1 _11912_ (.A1(\core.registers[16][25] ),
    .A2(net1511),
    .B1(_06810_),
    .C1(net1598),
    .X(_06825_));
 sky130_fd_sc_hd__mux2_1 _11913_ (.A0(\core.registers[18][25] ),
    .A1(\core.registers[19][25] ),
    .S(net1511),
    .X(_06826_));
 sky130_fd_sc_hd__a211o_1 _11914_ (.A1(net1613),
    .A2(_06826_),
    .B1(_06825_),
    .C1(net1586),
    .X(_06827_));
 sky130_fd_sc_hd__mux2_1 _11915_ (.A0(\core.registers[22][25] ),
    .A1(\core.registers[23][25] ),
    .S(net1511),
    .X(_06828_));
 sky130_fd_sc_hd__mux2_1 _11916_ (.A0(\core.registers[20][25] ),
    .A1(\core.registers[21][25] ),
    .S(net1507),
    .X(_06829_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(_06828_),
    .A1(_06829_),
    .S(net1597),
    .X(_06830_));
 sky130_fd_sc_hd__o211a_1 _11918_ (.A1(net1576),
    .A2(_06830_),
    .B1(_06827_),
    .C1(net1571),
    .X(_06831_));
 sky130_fd_sc_hd__a311o_1 _11919_ (.A1(net1567),
    .A2(_06821_),
    .A3(_06824_),
    .B1(_06831_),
    .C1(net1635),
    .X(_06832_));
 sky130_fd_sc_hd__a21o_2 _11920_ (.A1(_06818_),
    .A2(_06832_),
    .B1(net1157),
    .X(_06833_));
 sky130_fd_sc_hd__o211ai_4 _11921_ (.A1(net1153),
    .A2(net1111),
    .B1(_06833_),
    .C1(net1263),
    .Y(_06834_));
 sky130_fd_sc_hd__o21ai_1 _11922_ (.A1(net1192),
    .A2(_06834_),
    .B1(net1161),
    .Y(_06835_));
 sky130_fd_sc_hd__o21a_2 _11923_ (.A1(net1822),
    .A2(net1278),
    .B1(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__o22a_1 _11924_ (.A1(net1680),
    .A2(\core.registers[23][25] ),
    .B1(net1385),
    .B2(\core.registers[22][25] ),
    .X(_06837_));
 sky130_fd_sc_hd__or3_1 _11925_ (.A(net1680),
    .B(\core.registers[19][25] ),
    .C(net1442),
    .X(_06838_));
 sky130_fd_sc_hd__o221a_1 _11926_ (.A1(\core.registers[18][25] ),
    .A2(net1331),
    .B1(_06837_),
    .B2(net1431),
    .C1(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__mux4_1 _11927_ (.A0(\core.registers[16][25] ),
    .A1(\core.registers[17][25] ),
    .A2(\core.registers[20][25] ),
    .A3(\core.registers[21][25] ),
    .S0(net1382),
    .S1(net1444),
    .X(_06840_));
 sky130_fd_sc_hd__mux2_1 _11928_ (.A0(_06839_),
    .A1(_06840_),
    .S(net1465),
    .X(_06841_));
 sky130_fd_sc_hd__o22a_1 _11929_ (.A1(net1680),
    .A2(\core.registers[7][25] ),
    .B1(net1385),
    .B2(\core.registers[6][25] ),
    .X(_06842_));
 sky130_fd_sc_hd__or3_1 _11930_ (.A(net1680),
    .B(\core.registers[3][25] ),
    .C(net1442),
    .X(_06843_));
 sky130_fd_sc_hd__o221a_1 _11931_ (.A1(\core.registers[2][25] ),
    .A2(net1333),
    .B1(_06842_),
    .B2(net1432),
    .C1(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__mux4_1 _11932_ (.A0(\core.registers[0][25] ),
    .A1(\core.registers[1][25] ),
    .A2(\core.registers[4][25] ),
    .A3(\core.registers[5][25] ),
    .S0(net1385),
    .S1(net1443),
    .X(_06845_));
 sky130_fd_sc_hd__mux2_1 _11933_ (.A0(_06844_),
    .A1(_06845_),
    .S(net1466),
    .X(_06846_));
 sky130_fd_sc_hd__mux2_1 _11934_ (.A0(_06841_),
    .A1(_06846_),
    .S(net1460),
    .X(_06847_));
 sky130_fd_sc_hd__a221o_1 _11935_ (.A1(net1679),
    .A2(\core.registers[26][25] ),
    .B1(\core.registers[27][25] ),
    .B2(net1383),
    .C1(net1705),
    .X(_06848_));
 sky130_fd_sc_hd__mux2_1 _11936_ (.A0(\core.registers[24][25] ),
    .A1(\core.registers[25][25] ),
    .S(net1383),
    .X(_06849_));
 sky130_fd_sc_hd__o21ai_1 _11937_ (.A1(net1868),
    .A2(_06849_),
    .B1(_06848_),
    .Y(_06850_));
 sky130_fd_sc_hd__a221o_1 _11938_ (.A1(net1678),
    .A2(\core.registers[10][25] ),
    .B1(\core.registers[11][25] ),
    .B2(net1380),
    .C1(net1705),
    .X(_06851_));
 sky130_fd_sc_hd__a21o_1 _11939_ (.A1(\core.registers[8][25] ),
    .A2(net1373),
    .B1(net1868),
    .X(_06852_));
 sky130_fd_sc_hd__a21o_1 _11940_ (.A1(\core.registers[9][25] ),
    .A2(net1380),
    .B1(_06852_),
    .X(_06853_));
 sky130_fd_sc_hd__a21oi_2 _11941_ (.A1(_06851_),
    .A2(_06853_),
    .B1(net1853),
    .Y(_06854_));
 sky130_fd_sc_hd__a211o_1 _11942_ (.A1(net1854),
    .A2(_06850_),
    .B1(_06854_),
    .C1(net1862),
    .X(_06855_));
 sky130_fd_sc_hd__mux2_1 _11943_ (.A0(\core.registers[12][25] ),
    .A1(\core.registers[13][25] ),
    .S(net1379),
    .X(_06856_));
 sky130_fd_sc_hd__mux2_1 _11944_ (.A0(\core.registers[14][25] ),
    .A1(\core.registers[15][25] ),
    .S(net1379),
    .X(_06857_));
 sky130_fd_sc_hd__mux2_1 _11945_ (.A0(_06856_),
    .A1(_06857_),
    .S(net1480),
    .X(_06858_));
 sky130_fd_sc_hd__a221o_1 _11946_ (.A1(net1678),
    .A2(\core.registers[30][25] ),
    .B1(\core.registers[31][25] ),
    .B2(net1380),
    .C1(net1704),
    .X(_06859_));
 sky130_fd_sc_hd__mux2_1 _11947_ (.A0(\core.registers[28][25] ),
    .A1(\core.registers[29][25] ),
    .S(net1380),
    .X(_06860_));
 sky130_fd_sc_hd__o21a_1 _11948_ (.A1(net1868),
    .A2(_06860_),
    .B1(_06859_),
    .X(_06861_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(_06858_),
    .A1(_06861_),
    .S(net1853),
    .X(_06862_));
 sky130_fd_sc_hd__a21oi_1 _11950_ (.A1(net1862),
    .A2(_06862_),
    .B1(net1484),
    .Y(_06863_));
 sky130_fd_sc_hd__o2bb2a_2 _11951_ (.A1_N(_06855_),
    .A2_N(_06863_),
    .B1(net1489),
    .B2(_06847_),
    .X(_06864_));
 sky130_fd_sc_hd__a22o_2 _11952_ (.A1(net1068),
    .A2(net1111),
    .B1(_06864_),
    .B2(net1065),
    .X(_06865_));
 sky130_fd_sc_hd__mux2_8 _11953_ (.A0(net467),
    .A1(_06865_),
    .S(net1276),
    .X(_06866_));
 sky130_fd_sc_hd__nor2_1 _11954_ (.A(_06836_),
    .B(_06866_),
    .Y(_06867_));
 sky130_fd_sc_hd__and2_4 _11955_ (.A(_06836_),
    .B(_06866_),
    .X(_06868_));
 sky130_fd_sc_hd__nor2_4 _11956_ (.A(_06867_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__clkinv_4 _11957_ (.A(_06869_),
    .Y(_06870_));
 sky130_fd_sc_hd__and2b_1 _11958_ (.A_N(_06757_),
    .B(_06788_),
    .X(_06871_));
 sky130_fd_sc_hd__a21oi_2 _11959_ (.A1(_06717_),
    .A2(_06792_),
    .B1(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__xnor2_2 _11960_ (.A(_06870_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__or2_1 _11961_ (.A(_06791_),
    .B(_06869_),
    .X(_06874_));
 sky130_fd_sc_hd__a22o_1 _11962_ (.A1(\core.pipe1_resultRegister[27] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[27] ),
    .X(_06875_));
 sky130_fd_sc_hd__a21o_4 _11963_ (.A1(net1234),
    .A2(_05294_),
    .B1(net1237),
    .X(_06876_));
 sky130_fd_sc_hd__a21o_1 _11964_ (.A1(net1188),
    .A2(_06876_),
    .B1(_06875_),
    .X(_06877_));
 sky130_fd_sc_hd__or2_1 _11965_ (.A(\core.registers[6][27] ),
    .B(net1512),
    .X(_06878_));
 sky130_fd_sc_hd__or2_1 _11966_ (.A(\core.registers[17][27] ),
    .B(net1496),
    .X(_06879_));
 sky130_fd_sc_hd__mux2_1 _11967_ (.A0(\core.registers[28][27] ),
    .A1(\core.registers[29][27] ),
    .S(net1524),
    .X(_06880_));
 sky130_fd_sc_hd__a221o_1 _11968_ (.A1(net1722),
    .A2(\core.registers[30][27] ),
    .B1(\core.registers[31][27] ),
    .B2(net1524),
    .C1(net1737),
    .X(_06881_));
 sky130_fd_sc_hd__o21a_1 _11969_ (.A1(net1839),
    .A2(_06880_),
    .B1(_06881_),
    .X(_06882_));
 sky130_fd_sc_hd__mux2_1 _11970_ (.A0(\core.registers[14][27] ),
    .A1(\core.registers[15][27] ),
    .S(net1524),
    .X(_06883_));
 sky130_fd_sc_hd__mux2_1 _11971_ (.A0(\core.registers[12][27] ),
    .A1(\core.registers[13][27] ),
    .S(net1524),
    .X(_06884_));
 sky130_fd_sc_hd__mux2_1 _11972_ (.A0(_06883_),
    .A1(_06884_),
    .S(net1603),
    .X(_06885_));
 sky130_fd_sc_hd__mux2_1 _11973_ (.A0(_06882_),
    .A1(_06885_),
    .S(net1748),
    .X(_06886_));
 sky130_fd_sc_hd__or2_1 _11974_ (.A(\core.registers[24][27] ),
    .B(net1510),
    .X(_06887_));
 sky130_fd_sc_hd__o211a_1 _11975_ (.A1(\core.registers[25][27] ),
    .A2(net1493),
    .B1(_06887_),
    .C1(net1736),
    .X(_06888_));
 sky130_fd_sc_hd__a31o_1 _11976_ (.A1(net1839),
    .A2(net1720),
    .A3(\core.registers[26][27] ),
    .B1(net1748),
    .X(_06889_));
 sky130_fd_sc_hd__a31o_1 _11977_ (.A1(net1839),
    .A2(\core.registers[27][27] ),
    .A3(net1510),
    .B1(_06889_),
    .X(_06890_));
 sky130_fd_sc_hd__mux2_1 _11978_ (.A0(\core.registers[8][27] ),
    .A1(\core.registers[9][27] ),
    .S(net1524),
    .X(_06891_));
 sky130_fd_sc_hd__mux2_1 _11979_ (.A0(\core.registers[10][27] ),
    .A1(\core.registers[11][27] ),
    .S(net1510),
    .X(_06892_));
 sky130_fd_sc_hd__mux2_1 _11980_ (.A0(_06891_),
    .A1(_06892_),
    .S(net1612),
    .X(_06893_));
 sky130_fd_sc_hd__o221a_1 _11981_ (.A1(_06888_),
    .A2(_06890_),
    .B1(_06893_),
    .B2(net1824),
    .C1(net1744),
    .X(_06894_));
 sky130_fd_sc_hd__a211o_2 _11982_ (.A1(net1832),
    .A2(_06886_),
    .B1(_06894_),
    .C1(net1631),
    .X(_06895_));
 sky130_fd_sc_hd__o211a_1 _11983_ (.A1(net1720),
    .A2(\core.registers[7][27] ),
    .B1(net1612),
    .C1(_06878_),
    .X(_06896_));
 sky130_fd_sc_hd__mux2_1 _11984_ (.A0(\core.registers[4][27] ),
    .A1(\core.registers[5][27] ),
    .S(net1520),
    .X(_06897_));
 sky130_fd_sc_hd__a211o_1 _11985_ (.A1(net1597),
    .A2(_06897_),
    .B1(_06896_),
    .C1(net1576),
    .X(_06898_));
 sky130_fd_sc_hd__mux2_1 _11986_ (.A0(\core.registers[0][27] ),
    .A1(\core.registers[1][27] ),
    .S(net1521),
    .X(_06899_));
 sky130_fd_sc_hd__mux2_1 _11987_ (.A0(\core.registers[2][27] ),
    .A1(\core.registers[3][27] ),
    .S(net1521),
    .X(_06900_));
 sky130_fd_sc_hd__mux2_1 _11988_ (.A0(_06899_),
    .A1(_06900_),
    .S(net1616),
    .X(_06901_));
 sky130_fd_sc_hd__o211a_1 _11989_ (.A1(net1587),
    .A2(_06901_),
    .B1(_06898_),
    .C1(net1567),
    .X(_06902_));
 sky130_fd_sc_hd__o211a_1 _11990_ (.A1(\core.registers[16][27] ),
    .A2(net1525),
    .B1(_06879_),
    .C1(net1603),
    .X(_06903_));
 sky130_fd_sc_hd__mux2_1 _11991_ (.A0(\core.registers[18][27] ),
    .A1(\core.registers[19][27] ),
    .S(net1525),
    .X(_06904_));
 sky130_fd_sc_hd__a211o_1 _11992_ (.A1(net1617),
    .A2(_06904_),
    .B1(_06903_),
    .C1(net1587),
    .X(_06905_));
 sky130_fd_sc_hd__mux2_1 _11993_ (.A0(\core.registers[22][27] ),
    .A1(\core.registers[23][27] ),
    .S(net1525),
    .X(_06906_));
 sky130_fd_sc_hd__mux2_1 _11994_ (.A0(\core.registers[20][27] ),
    .A1(\core.registers[21][27] ),
    .S(net1525),
    .X(_06907_));
 sky130_fd_sc_hd__mux2_1 _11995_ (.A0(_06906_),
    .A1(_06907_),
    .S(net1603),
    .X(_06908_));
 sky130_fd_sc_hd__o211a_1 _11996_ (.A1(net1576),
    .A2(_06908_),
    .B1(_06905_),
    .C1(net1571),
    .X(_06909_));
 sky130_fd_sc_hd__o31a_1 _11997_ (.A1(net1635),
    .A2(_06902_),
    .A3(_06909_),
    .B1(_06895_),
    .X(_06910_));
 sky130_fd_sc_hd__o21a_1 _11998_ (.A1(net1157),
    .A2(_06910_),
    .B1(net1263),
    .X(_06911_));
 sky130_fd_sc_hd__o21ai_1 _11999_ (.A1(net1153),
    .A2(net1107),
    .B1(_06911_),
    .Y(_06912_));
 sky130_fd_sc_hd__o21ai_1 _12000_ (.A1(net1193),
    .A2(_06912_),
    .B1(net1162),
    .Y(_06913_));
 sky130_fd_sc_hd__o21a_1 _12001_ (.A1(net1820),
    .A2(net1278),
    .B1(_06913_),
    .X(_06914_));
 sky130_fd_sc_hd__o22a_1 _12002_ (.A1(net1685),
    .A2(\core.registers[23][27] ),
    .B1(net1396),
    .B2(\core.registers[22][27] ),
    .X(_06915_));
 sky130_fd_sc_hd__or3_1 _12003_ (.A(net1680),
    .B(\core.registers[19][27] ),
    .C(net1442),
    .X(_06916_));
 sky130_fd_sc_hd__o221a_1 _12004_ (.A1(\core.registers[18][27] ),
    .A2(net1331),
    .B1(_06915_),
    .B2(net1432),
    .C1(_06916_),
    .X(_06917_));
 sky130_fd_sc_hd__mux4_1 _12005_ (.A0(\core.registers[16][27] ),
    .A1(\core.registers[17][27] ),
    .A2(\core.registers[20][27] ),
    .A3(\core.registers[21][27] ),
    .S0(net1396),
    .S1(net1447),
    .X(_06918_));
 sky130_fd_sc_hd__mux2_1 _12006_ (.A0(_06917_),
    .A1(_06918_),
    .S(net1465),
    .X(_06919_));
 sky130_fd_sc_hd__o22a_1 _12007_ (.A1(net1681),
    .A2(\core.registers[7][27] ),
    .B1(net1392),
    .B2(\core.registers[6][27] ),
    .X(_06920_));
 sky130_fd_sc_hd__or3_1 _12008_ (.A(net1683),
    .B(\core.registers[3][27] ),
    .C(net1443),
    .X(_06921_));
 sky130_fd_sc_hd__o221a_1 _12009_ (.A1(\core.registers[2][27] ),
    .A2(net1331),
    .B1(_06920_),
    .B2(net1433),
    .C1(_06921_),
    .X(_06922_));
 sky130_fd_sc_hd__mux4_1 _12010_ (.A0(\core.registers[0][27] ),
    .A1(\core.registers[1][27] ),
    .A2(\core.registers[4][27] ),
    .A3(\core.registers[5][27] ),
    .S0(net1392),
    .S1(net1443),
    .X(_06923_));
 sky130_fd_sc_hd__mux2_1 _12011_ (.A0(_06922_),
    .A1(_06923_),
    .S(net1468),
    .X(_06924_));
 sky130_fd_sc_hd__mux2_1 _12012_ (.A0(_06919_),
    .A1(_06924_),
    .S(net1460),
    .X(_06925_));
 sky130_fd_sc_hd__mux2_1 _12013_ (.A0(\core.registers[24][27] ),
    .A1(\core.registers[25][27] ),
    .S(net1384),
    .X(_06926_));
 sky130_fd_sc_hd__a221o_1 _12014_ (.A1(net1679),
    .A2(\core.registers[26][27] ),
    .B1(\core.registers[27][27] ),
    .B2(net1384),
    .C1(net1705),
    .X(_06927_));
 sky130_fd_sc_hd__o21ai_1 _12015_ (.A1(net1869),
    .A2(_06926_),
    .B1(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__a221o_1 _12016_ (.A1(net1679),
    .A2(\core.registers[10][27] ),
    .B1(\core.registers[11][27] ),
    .B2(net1384),
    .C1(net1705),
    .X(_06929_));
 sky130_fd_sc_hd__a21o_1 _12017_ (.A1(\core.registers[8][27] ),
    .A2(net1374),
    .B1(net1870),
    .X(_06930_));
 sky130_fd_sc_hd__a21o_1 _12018_ (.A1(\core.registers[9][27] ),
    .A2(net1395),
    .B1(_06930_),
    .X(_06931_));
 sky130_fd_sc_hd__a21oi_1 _12019_ (.A1(_06929_),
    .A2(_06931_),
    .B1(net1854),
    .Y(_06932_));
 sky130_fd_sc_hd__a211o_1 _12020_ (.A1(net1854),
    .A2(_06928_),
    .B1(_06932_),
    .C1(net1862),
    .X(_06933_));
 sky130_fd_sc_hd__mux2_1 _12021_ (.A0(\core.registers[12][27] ),
    .A1(\core.registers[13][27] ),
    .S(net1395),
    .X(_06934_));
 sky130_fd_sc_hd__mux2_1 _12022_ (.A0(\core.registers[14][27] ),
    .A1(\core.registers[15][27] ),
    .S(net1395),
    .X(_06935_));
 sky130_fd_sc_hd__mux2_1 _12023_ (.A0(_06934_),
    .A1(_06935_),
    .S(net1481),
    .X(_06936_));
 sky130_fd_sc_hd__a221o_1 _12024_ (.A1(net1684),
    .A2(\core.registers[30][27] ),
    .B1(\core.registers[31][27] ),
    .B2(net1395),
    .C1(net1706),
    .X(_06937_));
 sky130_fd_sc_hd__mux2_1 _12025_ (.A0(\core.registers[28][27] ),
    .A1(\core.registers[29][27] ),
    .S(net1395),
    .X(_06938_));
 sky130_fd_sc_hd__o21a_1 _12026_ (.A1(net1870),
    .A2(_06938_),
    .B1(_06937_),
    .X(_06939_));
 sky130_fd_sc_hd__mux2_1 _12027_ (.A0(_06936_),
    .A1(_06939_),
    .S(net1855),
    .X(_06940_));
 sky130_fd_sc_hd__a21oi_1 _12028_ (.A1(net1863),
    .A2(_06940_),
    .B1(_04642_),
    .Y(_06941_));
 sky130_fd_sc_hd__a2bb2o_2 _12029_ (.A1_N(net1489),
    .A2_N(_06925_),
    .B1(_06933_),
    .B2(_06941_),
    .X(_06942_));
 sky130_fd_sc_hd__o2bb2a_2 _12030_ (.A1_N(net1068),
    .A2_N(net1107),
    .B1(_06942_),
    .B2(_04663_),
    .X(_06943_));
 sky130_fd_sc_hd__inv_2 _12031_ (.A(_06943_),
    .Y(_06944_));
 sky130_fd_sc_hd__mux2_8 _12032_ (.A0(net469),
    .A1(_06944_),
    .S(net1277),
    .X(_06945_));
 sky130_fd_sc_hd__inv_2 _12033_ (.A(_06945_),
    .Y(_06946_));
 sky130_fd_sc_hd__nor2_1 _12034_ (.A(_06914_),
    .B(_06945_),
    .Y(_06947_));
 sky130_fd_sc_hd__nand2_1 _12035_ (.A(_06914_),
    .B(_06945_),
    .Y(_06948_));
 sky130_fd_sc_hd__and2b_4 _12036_ (.A_N(_06947_),
    .B(_06948_),
    .X(_06949_));
 sky130_fd_sc_hd__inv_2 _12037_ (.A(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__a22o_2 _12038_ (.A1(\core.pipe1_resultRegister[26] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[26] ),
    .X(_06951_));
 sky130_fd_sc_hd__a21o_4 _12039_ (.A1(net1234),
    .A2(_05382_),
    .B1(net2014),
    .X(_06952_));
 sky130_fd_sc_hd__a21o_2 _12040_ (.A1(net1188),
    .A2(_06952_),
    .B1(_06951_),
    .X(_06953_));
 sky130_fd_sc_hd__or2_1 _12041_ (.A(\core.registers[1][26] ),
    .B(net1503),
    .X(_06954_));
 sky130_fd_sc_hd__or2_1 _12042_ (.A(\core.registers[6][26] ),
    .B(net1533),
    .X(_06955_));
 sky130_fd_sc_hd__or2_1 _12043_ (.A(\core.registers[17][26] ),
    .B(net1497),
    .X(_06956_));
 sky130_fd_sc_hd__or2_1 _12044_ (.A(\core.registers[29][26] ),
    .B(net1496),
    .X(_06957_));
 sky130_fd_sc_hd__o211a_1 _12045_ (.A1(\core.registers[28][26] ),
    .A2(net1523),
    .B1(_06957_),
    .C1(net1737),
    .X(_06958_));
 sky130_fd_sc_hd__a31o_1 _12046_ (.A1(net1841),
    .A2(net1722),
    .A3(\core.registers[30][26] ),
    .B1(net1749),
    .X(_06959_));
 sky130_fd_sc_hd__a31o_1 _12047_ (.A1(net1841),
    .A2(\core.registers[31][26] ),
    .A3(net1523),
    .B1(_06959_),
    .X(_06960_));
 sky130_fd_sc_hd__mux2_1 _12048_ (.A0(\core.registers[8][26] ),
    .A1(\core.registers[9][26] ),
    .S(net1523),
    .X(_06961_));
 sky130_fd_sc_hd__mux2_1 _12049_ (.A0(\core.registers[10][26] ),
    .A1(\core.registers[11][26] ),
    .S(net1523),
    .X(_06962_));
 sky130_fd_sc_hd__mux2_1 _12050_ (.A0(\core.registers[24][26] ),
    .A1(\core.registers[25][26] ),
    .S(net1523),
    .X(_06963_));
 sky130_fd_sc_hd__a221o_1 _12051_ (.A1(net1722),
    .A2(\core.registers[26][26] ),
    .B1(\core.registers[27][26] ),
    .B2(net1523),
    .C1(net1737),
    .X(_06964_));
 sky130_fd_sc_hd__mux2_1 _12052_ (.A0(\core.registers[12][26] ),
    .A1(\core.registers[13][26] ),
    .S(net1523),
    .X(_06965_));
 sky130_fd_sc_hd__mux2_1 _12053_ (.A0(\core.registers[14][26] ),
    .A1(\core.registers[15][26] ),
    .S(net1523),
    .X(_06966_));
 sky130_fd_sc_hd__mux2_1 _12054_ (.A0(_06965_),
    .A1(_06966_),
    .S(net1617),
    .X(_06967_));
 sky130_fd_sc_hd__o221a_1 _12055_ (.A1(_06958_),
    .A2(_06960_),
    .B1(_06967_),
    .B2(net1825),
    .C1(net1833),
    .X(_06968_));
 sky130_fd_sc_hd__mux2_1 _12056_ (.A0(_06961_),
    .A1(_06962_),
    .S(net1617),
    .X(_06969_));
 sky130_fd_sc_hd__o21a_1 _12057_ (.A1(net1841),
    .A2(_06963_),
    .B1(_06964_),
    .X(_06970_));
 sky130_fd_sc_hd__mux2_1 _12058_ (.A0(_06969_),
    .A1(_06970_),
    .S(net1825),
    .X(_06971_));
 sky130_fd_sc_hd__a211o_2 _12059_ (.A1(net1745),
    .A2(_06971_),
    .B1(_06968_),
    .C1(net1632),
    .X(_06972_));
 sky130_fd_sc_hd__o211a_1 _12060_ (.A1(net1723),
    .A2(\core.registers[7][26] ),
    .B1(net1619),
    .C1(_06955_),
    .X(_06973_));
 sky130_fd_sc_hd__mux2_1 _12061_ (.A0(\core.registers[4][26] ),
    .A1(\core.registers[5][26] ),
    .S(net1530),
    .X(_06974_));
 sky130_fd_sc_hd__a211o_1 _12062_ (.A1(net1602),
    .A2(_06974_),
    .B1(_06973_),
    .C1(net1578),
    .X(_06975_));
 sky130_fd_sc_hd__o211a_1 _12063_ (.A1(\core.registers[0][26] ),
    .A2(net1533),
    .B1(_06954_),
    .C1(net1604),
    .X(_06976_));
 sky130_fd_sc_hd__mux2_1 _12064_ (.A0(\core.registers[2][26] ),
    .A1(\core.registers[3][26] ),
    .S(net1533),
    .X(_06977_));
 sky130_fd_sc_hd__a211o_1 _12065_ (.A1(net1618),
    .A2(_06977_),
    .B1(_06976_),
    .C1(net1589),
    .X(_06978_));
 sky130_fd_sc_hd__o211a_1 _12066_ (.A1(\core.registers[16][26] ),
    .A2(net1530),
    .B1(_06956_),
    .C1(net1602),
    .X(_06979_));
 sky130_fd_sc_hd__mux2_1 _12067_ (.A0(\core.registers[18][26] ),
    .A1(\core.registers[19][26] ),
    .S(net1530),
    .X(_06980_));
 sky130_fd_sc_hd__a211o_1 _12068_ (.A1(net1618),
    .A2(_06980_),
    .B1(_06979_),
    .C1(net1589),
    .X(_06981_));
 sky130_fd_sc_hd__mux2_1 _12069_ (.A0(\core.registers[22][26] ),
    .A1(\core.registers[23][26] ),
    .S(net1530),
    .X(_06982_));
 sky130_fd_sc_hd__mux2_1 _12070_ (.A0(\core.registers[20][26] ),
    .A1(\core.registers[21][26] ),
    .S(net1530),
    .X(_06983_));
 sky130_fd_sc_hd__mux2_1 _12071_ (.A0(_06982_),
    .A1(_06983_),
    .S(net1602),
    .X(_06984_));
 sky130_fd_sc_hd__o211a_1 _12072_ (.A1(net1578),
    .A2(_06984_),
    .B1(_06981_),
    .C1(net1572),
    .X(_06985_));
 sky130_fd_sc_hd__a311o_1 _12073_ (.A1(net1568),
    .A2(_06975_),
    .A3(_06978_),
    .B1(_06985_),
    .C1(net1636),
    .X(_06986_));
 sky130_fd_sc_hd__a21o_2 _12074_ (.A1(_06972_),
    .A2(_06986_),
    .B1(net1158),
    .X(_06987_));
 sky130_fd_sc_hd__o211ai_4 _12075_ (.A1(net1154),
    .A2(net1103),
    .B1(_06987_),
    .C1(net1264),
    .Y(_06988_));
 sky130_fd_sc_hd__o21ai_2 _12076_ (.A1(net1193),
    .A2(_06988_),
    .B1(net1162),
    .Y(_06989_));
 sky130_fd_sc_hd__o21a_1 _12077_ (.A1(net1821),
    .A2(net1278),
    .B1(_06989_),
    .X(_06990_));
 sky130_fd_sc_hd__o22a_1 _12078_ (.A1(net1687),
    .A2(\core.registers[23][26] ),
    .B1(net1403),
    .B2(\core.registers[22][26] ),
    .X(_06991_));
 sky130_fd_sc_hd__or3_1 _12079_ (.A(net1687),
    .B(\core.registers[19][26] ),
    .C(net1448),
    .X(_06992_));
 sky130_fd_sc_hd__o221a_1 _12080_ (.A1(\core.registers[18][26] ),
    .A2(net1332),
    .B1(_06991_),
    .B2(net1436),
    .C1(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__mux4_1 _12081_ (.A0(\core.registers[16][26] ),
    .A1(\core.registers[17][26] ),
    .A2(\core.registers[20][26] ),
    .A3(\core.registers[21][26] ),
    .S0(net1403),
    .S1(net1448),
    .X(_06994_));
 sky130_fd_sc_hd__mux2_1 _12082_ (.A0(_06993_),
    .A1(_06994_),
    .S(net1470),
    .X(_06995_));
 sky130_fd_sc_hd__o22a_1 _12083_ (.A1(net1687),
    .A2(\core.registers[7][26] ),
    .B1(net1402),
    .B2(\core.registers[6][26] ),
    .X(_06996_));
 sky130_fd_sc_hd__or3_1 _12084_ (.A(net1687),
    .B(\core.registers[3][26] ),
    .C(net1448),
    .X(_06997_));
 sky130_fd_sc_hd__o221a_1 _12085_ (.A1(\core.registers[2][26] ),
    .A2(net1333),
    .B1(_06996_),
    .B2(net1436),
    .C1(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__mux4_1 _12086_ (.A0(\core.registers[0][26] ),
    .A1(\core.registers[1][26] ),
    .A2(\core.registers[4][26] ),
    .A3(\core.registers[5][26] ),
    .S0(net1402),
    .S1(net1448),
    .X(_06999_));
 sky130_fd_sc_hd__mux2_1 _12087_ (.A0(_06998_),
    .A1(_06999_),
    .S(net1469),
    .X(_07000_));
 sky130_fd_sc_hd__mux2_1 _12088_ (.A0(_06995_),
    .A1(_07000_),
    .S(net1461),
    .X(_07001_));
 sky130_fd_sc_hd__mux2_1 _12089_ (.A0(\core.registers[14][26] ),
    .A1(\core.registers[15][26] ),
    .S(net1394),
    .X(_07002_));
 sky130_fd_sc_hd__mux2_1 _12090_ (.A0(\core.registers[12][26] ),
    .A1(\core.registers[13][26] ),
    .S(net1394),
    .X(_07003_));
 sky130_fd_sc_hd__mux2_1 _12091_ (.A0(_07002_),
    .A1(_07003_),
    .S(net1469),
    .X(_07004_));
 sky130_fd_sc_hd__mux2_1 _12092_ (.A0(\core.registers[28][26] ),
    .A1(\core.registers[29][26] ),
    .S(net1394),
    .X(_07005_));
 sky130_fd_sc_hd__a221o_1 _12093_ (.A1(net1684),
    .A2(\core.registers[30][26] ),
    .B1(\core.registers[31][26] ),
    .B2(net1394),
    .C1(net1706),
    .X(_07006_));
 sky130_fd_sc_hd__o21ai_1 _12094_ (.A1(net1870),
    .A2(_07005_),
    .B1(_07006_),
    .Y(_07007_));
 sky130_fd_sc_hd__nand2_1 _12095_ (.A(net1855),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__o211a_1 _12096_ (.A1(net1855),
    .A2(_07004_),
    .B1(_07008_),
    .C1(net1863),
    .X(_07009_));
 sky130_fd_sc_hd__mux2_1 _12097_ (.A0(\core.registers[24][26] ),
    .A1(\core.registers[25][26] ),
    .S(net1394),
    .X(_07010_));
 sky130_fd_sc_hd__a221o_1 _12098_ (.A1(net1684),
    .A2(\core.registers[26][26] ),
    .B1(\core.registers[27][26] ),
    .B2(net1394),
    .C1(net1706),
    .X(_07011_));
 sky130_fd_sc_hd__o21ai_1 _12099_ (.A1(net1870),
    .A2(_07010_),
    .B1(_07011_),
    .Y(_07012_));
 sky130_fd_sc_hd__o21a_1 _12100_ (.A1(\core.registers[8][26] ),
    .A2(net1394),
    .B1(net1706),
    .X(_07013_));
 sky130_fd_sc_hd__o21ai_1 _12101_ (.A1(\core.registers[9][26] ),
    .A2(net1374),
    .B1(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__a22o_1 _12102_ (.A1(net1684),
    .A2(\core.registers[10][26] ),
    .B1(\core.registers[11][26] ),
    .B2(net1394),
    .X(_07015_));
 sky130_fd_sc_hd__a21oi_1 _12103_ (.A1(net1870),
    .A2(_07015_),
    .B1(net1855),
    .Y(_07016_));
 sky130_fd_sc_hd__a221o_1 _12104_ (.A1(net1855),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07016_),
    .C1(net1863),
    .X(_07017_));
 sky130_fd_sc_hd__or3b_2 _12105_ (.A(net1486),
    .B(_07009_),
    .C_N(_07017_),
    .X(_07018_));
 sky130_fd_sc_hd__o21a_2 _12106_ (.A1(_04641_),
    .A2(_07001_),
    .B1(_07018_),
    .X(_07019_));
 sky130_fd_sc_hd__a22o_4 _12107_ (.A1(net1069),
    .A2(net1103),
    .B1(_07019_),
    .B2(net1065),
    .X(_07020_));
 sky130_fd_sc_hd__mux2_8 _12108_ (.A0(net468),
    .A1(_07020_),
    .S(net1276),
    .X(_07021_));
 sky130_fd_sc_hd__nor2_2 _12109_ (.A(_06990_),
    .B(_07021_),
    .Y(_07022_));
 sky130_fd_sc_hd__nand2_2 _12110_ (.A(_06990_),
    .B(_07021_),
    .Y(_07023_));
 sky130_fd_sc_hd__nand2b_4 _12111_ (.A_N(_07022_),
    .B(_07023_),
    .Y(_07024_));
 sky130_fd_sc_hd__or3b_1 _12112_ (.A(_06874_),
    .B(_06949_),
    .C_N(_07024_),
    .X(_07025_));
 sky130_fd_sc_hd__a21o_2 _12113_ (.A1(_06714_),
    .A2(_06716_),
    .B1(_07025_),
    .X(_07026_));
 sky130_fd_sc_hd__nand2b_1 _12114_ (.A_N(_06990_),
    .B(_07021_),
    .Y(_07027_));
 sky130_fd_sc_hd__and2b_1 _12115_ (.A_N(_06836_),
    .B(_06866_),
    .X(_07028_));
 sky130_fd_sc_hd__a21o_1 _12116_ (.A1(_06870_),
    .A2(_06871_),
    .B1(_07028_),
    .X(_07029_));
 sky130_fd_sc_hd__nand2_1 _12117_ (.A(_07024_),
    .B(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__a21o_1 _12118_ (.A1(_07027_),
    .A2(_07030_),
    .B1(_06949_),
    .X(_07031_));
 sky130_fd_sc_hd__o21a_1 _12119_ (.A1(_06914_),
    .A2(_06946_),
    .B1(_07031_),
    .X(_07032_));
 sky130_fd_sc_hd__a221o_1 _12120_ (.A1(net1719),
    .A2(\core.registers[26][28] ),
    .B1(\core.registers[27][28] ),
    .B2(net1516),
    .C1(net1736),
    .X(_07033_));
 sky130_fd_sc_hd__mux2_1 _12121_ (.A0(\core.registers[24][28] ),
    .A1(\core.registers[25][28] ),
    .S(net1516),
    .X(_07034_));
 sky130_fd_sc_hd__o21ai_1 _12122_ (.A1(net1843),
    .A2(_07034_),
    .B1(_07033_),
    .Y(_07035_));
 sky130_fd_sc_hd__a221o_1 _12123_ (.A1(net1721),
    .A2(\core.registers[30][28] ),
    .B1(\core.registers[31][28] ),
    .B2(net1520),
    .C1(net1736),
    .X(_07036_));
 sky130_fd_sc_hd__mux2_1 _12124_ (.A0(\core.registers[28][28] ),
    .A1(\core.registers[29][28] ),
    .S(net1520),
    .X(_07037_));
 sky130_fd_sc_hd__o21a_1 _12125_ (.A1(net1843),
    .A2(_07037_),
    .B1(_07036_),
    .X(_07038_));
 sky130_fd_sc_hd__mux2_1 _12126_ (.A0(\core.registers[12][28] ),
    .A1(\core.registers[13][28] ),
    .S(net1514),
    .X(_07039_));
 sky130_fd_sc_hd__mux2_1 _12127_ (.A0(\core.registers[14][28] ),
    .A1(\core.registers[15][28] ),
    .S(net1514),
    .X(_07040_));
 sky130_fd_sc_hd__mux2_1 _12128_ (.A0(_07039_),
    .A1(_07040_),
    .S(net1614),
    .X(_07041_));
 sky130_fd_sc_hd__mux2_1 _12129_ (.A0(_07038_),
    .A1(_07041_),
    .S(net1748),
    .X(_07042_));
 sky130_fd_sc_hd__or2_1 _12130_ (.A(\core.registers[6][28] ),
    .B(net1518),
    .X(_07043_));
 sky130_fd_sc_hd__or2_1 _12131_ (.A(\core.registers[17][28] ),
    .B(net1494),
    .X(_07044_));
 sky130_fd_sc_hd__mux2_1 _12132_ (.A0(\core.registers[8][28] ),
    .A1(\core.registers[9][28] ),
    .S(net1514),
    .X(_07045_));
 sky130_fd_sc_hd__mux2_1 _12133_ (.A0(\core.registers[10][28] ),
    .A1(\core.registers[11][28] ),
    .S(net1514),
    .X(_07046_));
 sky130_fd_sc_hd__mux2_1 _12134_ (.A0(_07045_),
    .A1(_07046_),
    .S(net1614),
    .X(_07047_));
 sky130_fd_sc_hd__or2_1 _12135_ (.A(net1824),
    .B(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__a21oi_1 _12136_ (.A1(net1824),
    .A2(_07035_),
    .B1(net1833),
    .Y(_07049_));
 sky130_fd_sc_hd__a221o_1 _12137_ (.A1(net1832),
    .A2(_07042_),
    .B1(_07048_),
    .B2(_07049_),
    .C1(net1631),
    .X(_07050_));
 sky130_fd_sc_hd__o211a_1 _12138_ (.A1(net1721),
    .A2(\core.registers[7][28] ),
    .B1(net1615),
    .C1(_07043_),
    .X(_07051_));
 sky130_fd_sc_hd__mux2_1 _12139_ (.A0(\core.registers[4][28] ),
    .A1(\core.registers[5][28] ),
    .S(net1518),
    .X(_07052_));
 sky130_fd_sc_hd__a211o_1 _12140_ (.A1(net1599),
    .A2(_07052_),
    .B1(_07051_),
    .C1(net1575),
    .X(_07053_));
 sky130_fd_sc_hd__mux2_1 _12141_ (.A0(\core.registers[0][28] ),
    .A1(\core.registers[1][28] ),
    .S(net1519),
    .X(_07054_));
 sky130_fd_sc_hd__mux2_1 _12142_ (.A0(\core.registers[2][28] ),
    .A1(\core.registers[3][28] ),
    .S(net1519),
    .X(_07055_));
 sky130_fd_sc_hd__mux2_1 _12143_ (.A0(_07054_),
    .A1(_07055_),
    .S(net1615),
    .X(_07056_));
 sky130_fd_sc_hd__o211a_1 _12144_ (.A1(net1587),
    .A2(_07056_),
    .B1(_07053_),
    .C1(net1567),
    .X(_07057_));
 sky130_fd_sc_hd__o211a_1 _12145_ (.A1(\core.registers[16][28] ),
    .A2(net1517),
    .B1(_07044_),
    .C1(net1599),
    .X(_07058_));
 sky130_fd_sc_hd__mux2_1 _12146_ (.A0(\core.registers[18][28] ),
    .A1(\core.registers[19][28] ),
    .S(net1517),
    .X(_07059_));
 sky130_fd_sc_hd__a211o_1 _12147_ (.A1(net1614),
    .A2(_07059_),
    .B1(_07058_),
    .C1(net1586),
    .X(_07060_));
 sky130_fd_sc_hd__mux2_1 _12148_ (.A0(\core.registers[22][28] ),
    .A1(\core.registers[23][28] ),
    .S(net1519),
    .X(_07061_));
 sky130_fd_sc_hd__mux2_1 _12149_ (.A0(\core.registers[20][28] ),
    .A1(\core.registers[21][28] ),
    .S(net1515),
    .X(_07062_));
 sky130_fd_sc_hd__mux2_1 _12150_ (.A0(_07061_),
    .A1(_07062_),
    .S(net1599),
    .X(_07063_));
 sky130_fd_sc_hd__o211a_1 _12151_ (.A1(net1576),
    .A2(_07063_),
    .B1(_07060_),
    .C1(net1571),
    .X(_07064_));
 sky130_fd_sc_hd__o31a_1 _12152_ (.A1(net1635),
    .A2(_07057_),
    .A3(_07064_),
    .B1(_07050_),
    .X(_07065_));
 sky130_fd_sc_hd__o21a_1 _12153_ (.A1(net1157),
    .A2(_07065_),
    .B1(net1263),
    .X(_07066_));
 sky130_fd_sc_hd__a21o_4 _12154_ (.A1(net1235),
    .A2(_04953_),
    .B1(net1237),
    .X(_07067_));
 sky130_fd_sc_hd__a22o_1 _12155_ (.A1(\core.pipe1_resultRegister[28] ),
    .A2(net1238),
    .B1(net1267),
    .B2(\core.pipe1_csrData[28] ),
    .X(_07068_));
 sky130_fd_sc_hd__a21o_1 _12156_ (.A1(net1188),
    .A2(_07067_),
    .B1(_07068_),
    .X(_07069_));
 sky130_fd_sc_hd__o21ai_4 _12157_ (.A1(net1153),
    .A2(net1099),
    .B1(_07066_),
    .Y(_07070_));
 sky130_fd_sc_hd__o21ai_1 _12158_ (.A1(net1193),
    .A2(_07070_),
    .B1(net1161),
    .Y(_07071_));
 sky130_fd_sc_hd__o21a_2 _12159_ (.A1(net1819),
    .A2(net1279),
    .B1(_07071_),
    .X(_07072_));
 sky130_fd_sc_hd__and3_1 _12160_ (.A(\core.pipe0_currentInstruction[15] ),
    .B(\core.registers[23][28] ),
    .C(net1666),
    .X(_07073_));
 sky130_fd_sc_hd__mux2_1 _12161_ (.A0(\core.registers[4][28] ),
    .A1(\core.registers[5][28] ),
    .S(net1390),
    .X(_07074_));
 sky130_fd_sc_hd__mux2_1 _12162_ (.A0(\core.registers[6][28] ),
    .A1(\core.registers[7][28] ),
    .S(net1390),
    .X(_07075_));
 sky130_fd_sc_hd__mux2_1 _12163_ (.A0(_07074_),
    .A1(_07075_),
    .S(net1478),
    .X(_07076_));
 sky130_fd_sc_hd__mux2_1 _12164_ (.A0(\core.registers[2][28] ),
    .A1(\core.registers[3][28] ),
    .S(net1391),
    .X(_07077_));
 sky130_fd_sc_hd__mux2_1 _12165_ (.A0(\core.registers[0][28] ),
    .A1(\core.registers[1][28] ),
    .S(net1391),
    .X(_07078_));
 sky130_fd_sc_hd__or2_1 _12166_ (.A(net1479),
    .B(_07078_),
    .X(_07079_));
 sky130_fd_sc_hd__o211a_1 _12167_ (.A1(net1467),
    .A2(_07077_),
    .B1(_07079_),
    .C1(net1434),
    .X(_07080_));
 sky130_fd_sc_hd__a211o_1 _12168_ (.A1(net1446),
    .A2(_07076_),
    .B1(_07080_),
    .C1(net1490),
    .X(_07081_));
 sky130_fd_sc_hd__mux2_1 _12169_ (.A0(\core.registers[10][28] ),
    .A1(\core.registers[11][28] ),
    .S(net1388),
    .X(_07082_));
 sky130_fd_sc_hd__mux2_1 _12170_ (.A0(\core.registers[8][28] ),
    .A1(\core.registers[9][28] ),
    .S(net1388),
    .X(_07083_));
 sky130_fd_sc_hd__or2_1 _12171_ (.A(net1478),
    .B(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__o211a_1 _12172_ (.A1(net1467),
    .A2(_07082_),
    .B1(_07084_),
    .C1(net1434),
    .X(_07085_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(\core.registers[12][28] ),
    .A1(\core.registers[13][28] ),
    .S(net1388),
    .X(_07086_));
 sky130_fd_sc_hd__mux2_1 _12174_ (.A0(\core.registers[14][28] ),
    .A1(\core.registers[15][28] ),
    .S(net1388),
    .X(_07087_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(_07086_),
    .A1(_07087_),
    .S(net1478),
    .X(_07088_));
 sky130_fd_sc_hd__a211o_1 _12176_ (.A1(net1445),
    .A2(_07088_),
    .B1(_07085_),
    .C1(net1485),
    .X(_07089_));
 sky130_fd_sc_hd__a211o_1 _12177_ (.A1(net1682),
    .A2(\core.registers[22][28] ),
    .B1(net1468),
    .C1(_07073_),
    .X(_07090_));
 sky130_fd_sc_hd__mux2_1 _12178_ (.A0(\core.registers[20][28] ),
    .A1(\core.registers[21][28] ),
    .S(net1389),
    .X(_07091_));
 sky130_fd_sc_hd__o211a_1 _12179_ (.A1(net1478),
    .A2(_07091_),
    .B1(_07090_),
    .C1(net1445),
    .X(_07092_));
 sky130_fd_sc_hd__mux2_1 _12180_ (.A0(\core.registers[16][28] ),
    .A1(\core.registers[17][28] ),
    .S(net1390),
    .X(_07093_));
 sky130_fd_sc_hd__or2_1 _12181_ (.A(net1479),
    .B(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__mux2_1 _12182_ (.A0(\core.registers[18][28] ),
    .A1(\core.registers[19][28] ),
    .S(net1390),
    .X(_07095_));
 sky130_fd_sc_hd__o211a_1 _12183_ (.A1(net1467),
    .A2(_07095_),
    .B1(_07094_),
    .C1(net1434),
    .X(_07096_));
 sky130_fd_sc_hd__mux2_1 _12184_ (.A0(\core.registers[28][28] ),
    .A1(\core.registers[29][28] ),
    .S(net1392),
    .X(_07097_));
 sky130_fd_sc_hd__mux2_1 _12185_ (.A0(\core.registers[30][28] ),
    .A1(\core.registers[31][28] ),
    .S(net1392),
    .X(_07098_));
 sky130_fd_sc_hd__mux2_1 _12186_ (.A0(_07097_),
    .A1(_07098_),
    .S(net1479),
    .X(_07099_));
 sky130_fd_sc_hd__mux2_1 _12187_ (.A0(\core.registers[26][28] ),
    .A1(\core.registers[27][28] ),
    .S(net1389),
    .X(_07100_));
 sky130_fd_sc_hd__mux2_1 _12188_ (.A0(\core.registers[24][28] ),
    .A1(\core.registers[25][28] ),
    .S(net1389),
    .X(_07101_));
 sky130_fd_sc_hd__or2_1 _12189_ (.A(net1478),
    .B(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__o211a_1 _12190_ (.A1(net1467),
    .A2(_07100_),
    .B1(_07102_),
    .C1(net1433),
    .X(_07103_));
 sky130_fd_sc_hd__a211o_1 _12191_ (.A1(net1444),
    .A2(_07099_),
    .B1(_07103_),
    .C1(net1485),
    .X(_07104_));
 sky130_fd_sc_hd__o311a_1 _12192_ (.A1(net1489),
    .A2(_07092_),
    .A3(_07096_),
    .B1(_07104_),
    .C1(net1464),
    .X(_07105_));
 sky130_fd_sc_hd__a31o_1 _12193_ (.A1(net1460),
    .A2(_07081_),
    .A3(_07089_),
    .B1(_07105_),
    .X(_07106_));
 sky130_fd_sc_hd__a22o_2 _12194_ (.A1(net1068),
    .A2(net1099),
    .B1(_07106_),
    .B2(net1065),
    .X(_07107_));
 sky130_fd_sc_hd__mux2_8 _12195_ (.A0(net470),
    .A1(_07107_),
    .S(net1276),
    .X(_07108_));
 sky130_fd_sc_hd__inv_2 _12196_ (.A(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__nor2_2 _12197_ (.A(_07072_),
    .B(_07108_),
    .Y(_07110_));
 sky130_fd_sc_hd__nand2_2 _12198_ (.A(_07072_),
    .B(_07108_),
    .Y(_07111_));
 sky130_fd_sc_hd__nand2b_2 _12199_ (.A_N(_07110_),
    .B(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__clkinv_4 _12200_ (.A(_07112_),
    .Y(_07113_));
 sky130_fd_sc_hd__a21o_2 _12201_ (.A1(_07026_),
    .A2(_07032_),
    .B1(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__nand3_1 _12202_ (.A(_07026_),
    .B(_07032_),
    .C(_07113_),
    .Y(_07115_));
 sky130_fd_sc_hd__and2_1 _12203_ (.A(_07114_),
    .B(_07115_),
    .X(_07116_));
 sky130_fd_sc_hd__a21oi_1 _12204_ (.A1(_06714_),
    .A2(_06716_),
    .B1(_06874_),
    .Y(_07117_));
 sky130_fd_sc_hd__o21ai_2 _12205_ (.A1(_07029_),
    .A2(_07117_),
    .B1(_07024_),
    .Y(_07118_));
 sky130_fd_sc_hd__or3_1 _12206_ (.A(_07024_),
    .B(_07029_),
    .C(_07117_),
    .X(_07119_));
 sky130_fd_sc_hd__nand2_2 _12207_ (.A(_07118_),
    .B(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__a22o_2 _12208_ (.A1(\core.pipe1_resultRegister[29] ),
    .A2(net1239),
    .B1(net1268),
    .B2(\core.pipe1_csrData[29] ),
    .X(_07121_));
 sky130_fd_sc_hd__a21o_1 _12209_ (.A1(net1235),
    .A2(_05036_),
    .B1(net1237),
    .X(_07122_));
 sky130_fd_sc_hd__a21o_4 _12210_ (.A1(net1190),
    .A2(_07122_),
    .B1(_07121_),
    .X(_07123_));
 sky130_fd_sc_hd__or2_1 _12211_ (.A(\core.registers[1][29] ),
    .B(net1501),
    .X(_07124_));
 sky130_fd_sc_hd__or2_1 _12212_ (.A(\core.registers[6][29] ),
    .B(net1562),
    .X(_07125_));
 sky130_fd_sc_hd__or2_1 _12213_ (.A(\core.registers[17][29] ),
    .B(net1502),
    .X(_07126_));
 sky130_fd_sc_hd__or2_1 _12214_ (.A(\core.registers[28][29] ),
    .B(net1547),
    .X(_07127_));
 sky130_fd_sc_hd__o211a_1 _12215_ (.A1(\core.registers[29][29] ),
    .A2(net1502),
    .B1(_07127_),
    .C1(net1740),
    .X(_07128_));
 sky130_fd_sc_hd__a31o_1 _12216_ (.A1(net1845),
    .A2(net1732),
    .A3(\core.registers[30][29] ),
    .B1(net1750),
    .X(_07129_));
 sky130_fd_sc_hd__a31o_1 _12217_ (.A1(net1845),
    .A2(\core.registers[31][29] ),
    .A3(net1547),
    .B1(_07129_),
    .X(_07130_));
 sky130_fd_sc_hd__mux2_1 _12218_ (.A0(\core.registers[8][29] ),
    .A1(\core.registers[9][29] ),
    .S(net1551),
    .X(_07131_));
 sky130_fd_sc_hd__mux2_1 _12219_ (.A0(\core.registers[10][29] ),
    .A1(\core.registers[11][29] ),
    .S(net1552),
    .X(_07132_));
 sky130_fd_sc_hd__mux2_1 _12220_ (.A0(\core.registers[24][29] ),
    .A1(\core.registers[25][29] ),
    .S(net1551),
    .X(_07133_));
 sky130_fd_sc_hd__a221o_1 _12221_ (.A1(net1731),
    .A2(\core.registers[26][29] ),
    .B1(\core.registers[27][29] ),
    .B2(net1551),
    .C1(net1740),
    .X(_07134_));
 sky130_fd_sc_hd__mux2_1 _12222_ (.A0(\core.registers[12][29] ),
    .A1(\core.registers[13][29] ),
    .S(net1548),
    .X(_07135_));
 sky130_fd_sc_hd__mux2_1 _12223_ (.A0(\core.registers[14][29] ),
    .A1(\core.registers[15][29] ),
    .S(net1547),
    .X(_07136_));
 sky130_fd_sc_hd__mux2_1 _12224_ (.A0(_07135_),
    .A1(_07136_),
    .S(net1626),
    .X(_07137_));
 sky130_fd_sc_hd__o221a_1 _12225_ (.A1(_07128_),
    .A2(_07130_),
    .B1(_07137_),
    .B2(net1826),
    .C1(net1834),
    .X(_07138_));
 sky130_fd_sc_hd__mux2_1 _12226_ (.A0(_07131_),
    .A1(_07132_),
    .S(net1624),
    .X(_07139_));
 sky130_fd_sc_hd__o21a_1 _12227_ (.A1(net1845),
    .A2(_07133_),
    .B1(_07134_),
    .X(_07140_));
 sky130_fd_sc_hd__mux2_1 _12228_ (.A0(_07139_),
    .A1(_07140_),
    .S(net1826),
    .X(_07141_));
 sky130_fd_sc_hd__a211o_2 _12229_ (.A1(net1747),
    .A2(_07141_),
    .B1(_07138_),
    .C1(net1634),
    .X(_07142_));
 sky130_fd_sc_hd__o211a_1 _12230_ (.A1(net1733),
    .A2(\core.registers[7][29] ),
    .B1(net1628),
    .C1(_07125_),
    .X(_07143_));
 sky130_fd_sc_hd__mux2_1 _12231_ (.A0(\core.registers[4][29] ),
    .A1(\core.registers[5][29] ),
    .S(net1563),
    .X(_07144_));
 sky130_fd_sc_hd__a211o_1 _12232_ (.A1(net1608),
    .A2(_07144_),
    .B1(_07143_),
    .C1(net1582),
    .X(_07145_));
 sky130_fd_sc_hd__o211a_1 _12233_ (.A1(\core.registers[0][29] ),
    .A2(net1563),
    .B1(_07124_),
    .C1(net1607),
    .X(_07146_));
 sky130_fd_sc_hd__mux2_1 _12234_ (.A0(\core.registers[2][29] ),
    .A1(\core.registers[3][29] ),
    .S(net1563),
    .X(_07147_));
 sky130_fd_sc_hd__a211o_1 _12235_ (.A1(net1627),
    .A2(_07147_),
    .B1(_07146_),
    .C1(net1593),
    .X(_07148_));
 sky130_fd_sc_hd__o211a_1 _12236_ (.A1(\core.registers[16][29] ),
    .A2(net1562),
    .B1(_07126_),
    .C1(net1608),
    .X(_07149_));
 sky130_fd_sc_hd__mux2_1 _12237_ (.A0(\core.registers[18][29] ),
    .A1(\core.registers[19][29] ),
    .S(net1562),
    .X(_07150_));
 sky130_fd_sc_hd__a211o_1 _12238_ (.A1(net1628),
    .A2(_07150_),
    .B1(_07149_),
    .C1(net1593),
    .X(_07151_));
 sky130_fd_sc_hd__mux2_1 _12239_ (.A0(\core.registers[22][29] ),
    .A1(\core.registers[23][29] ),
    .S(net1562),
    .X(_07152_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(\core.registers[20][29] ),
    .A1(\core.registers[21][29] ),
    .S(net1562),
    .X(_07153_));
 sky130_fd_sc_hd__mux2_1 _12241_ (.A0(_07152_),
    .A1(_07153_),
    .S(net1608),
    .X(_07154_));
 sky130_fd_sc_hd__o211a_1 _12242_ (.A1(net1582),
    .A2(_07154_),
    .B1(_07151_),
    .C1(net1574),
    .X(_07155_));
 sky130_fd_sc_hd__a311o_2 _12243_ (.A1(net1569),
    .A2(_07145_),
    .A3(_07148_),
    .B1(_07155_),
    .C1(net1638),
    .X(_07156_));
 sky130_fd_sc_hd__a21o_2 _12244_ (.A1(_07142_),
    .A2(_07156_),
    .B1(net1160),
    .X(_07157_));
 sky130_fd_sc_hd__o211ai_4 _12245_ (.A1(net1155),
    .A2(net1095),
    .B1(_07157_),
    .C1(net1266),
    .Y(_07158_));
 sky130_fd_sc_hd__o21a_2 _12246_ (.A1(net1193),
    .A2(_07158_),
    .B1(net1162),
    .X(_07159_));
 sky130_fd_sc_hd__a21oi_4 _12247_ (.A1(_04414_),
    .A2(net1286),
    .B1(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__o22a_1 _12248_ (.A1(net1700),
    .A2(\core.registers[23][29] ),
    .B1(net1429),
    .B2(\core.registers[22][29] ),
    .X(_07161_));
 sky130_fd_sc_hd__or3_1 _12249_ (.A(net1700),
    .B(\core.registers[19][29] ),
    .C(net1457),
    .X(_07162_));
 sky130_fd_sc_hd__o221a_1 _12250_ (.A1(\core.registers[18][29] ),
    .A2(net1336),
    .B1(_07161_),
    .B2(net1440),
    .C1(_07162_),
    .X(_07163_));
 sky130_fd_sc_hd__mux4_1 _12251_ (.A0(\core.registers[16][29] ),
    .A1(\core.registers[17][29] ),
    .A2(\core.registers[20][29] ),
    .A3(\core.registers[21][29] ),
    .S0(net1428),
    .S1(net1457),
    .X(_07164_));
 sky130_fd_sc_hd__mux2_1 _12252_ (.A0(_07163_),
    .A1(_07164_),
    .S(net1475),
    .X(_07165_));
 sky130_fd_sc_hd__o22a_1 _12253_ (.A1(net1700),
    .A2(\core.registers[7][29] ),
    .B1(net1428),
    .B2(\core.registers[6][29] ),
    .X(_07166_));
 sky130_fd_sc_hd__or3_1 _12254_ (.A(net1702),
    .B(\core.registers[3][29] ),
    .C(net1458),
    .X(_07167_));
 sky130_fd_sc_hd__o221a_1 _12255_ (.A1(\core.registers[2][29] ),
    .A2(net1336),
    .B1(_07166_),
    .B2(net1441),
    .C1(_07167_),
    .X(_07168_));
 sky130_fd_sc_hd__mux4_1 _12256_ (.A0(\core.registers[0][29] ),
    .A1(\core.registers[1][29] ),
    .A2(\core.registers[4][29] ),
    .A3(\core.registers[5][29] ),
    .S0(net1428),
    .S1(net1457),
    .X(_07169_));
 sky130_fd_sc_hd__mux2_1 _12257_ (.A0(_07168_),
    .A1(_07169_),
    .S(net1475),
    .X(_07170_));
 sky130_fd_sc_hd__mux2_2 _12258_ (.A0(_07165_),
    .A1(_07170_),
    .S(net1462),
    .X(_07171_));
 sky130_fd_sc_hd__mux2_1 _12259_ (.A0(\core.registers[14][29] ),
    .A1(\core.registers[15][29] ),
    .S(net1415),
    .X(_07172_));
 sky130_fd_sc_hd__mux2_1 _12260_ (.A0(\core.registers[12][29] ),
    .A1(\core.registers[13][29] ),
    .S(net1416),
    .X(_07173_));
 sky130_fd_sc_hd__mux2_1 _12261_ (.A0(_07172_),
    .A1(_07173_),
    .S(net1474),
    .X(_07174_));
 sky130_fd_sc_hd__mux2_1 _12262_ (.A0(\core.registers[28][29] ),
    .A1(\core.registers[29][29] ),
    .S(net1415),
    .X(_07175_));
 sky130_fd_sc_hd__a221o_1 _12263_ (.A1(net1695),
    .A2(\core.registers[30][29] ),
    .B1(\core.registers[31][29] ),
    .B2(net1415),
    .C1(net1713),
    .X(_07176_));
 sky130_fd_sc_hd__o21ai_1 _12264_ (.A1(net1875),
    .A2(_07175_),
    .B1(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__nand2_1 _12265_ (.A(net1858),
    .B(_07177_),
    .Y(_07178_));
 sky130_fd_sc_hd__o211a_1 _12266_ (.A1(net1858),
    .A2(_07174_),
    .B1(_07178_),
    .C1(net1864),
    .X(_07179_));
 sky130_fd_sc_hd__a221o_1 _12267_ (.A1(net1698),
    .A2(\core.registers[26][29] ),
    .B1(\core.registers[27][29] ),
    .B2(net1419),
    .C1(net1709),
    .X(_07180_));
 sky130_fd_sc_hd__mux2_1 _12268_ (.A0(\core.registers[24][29] ),
    .A1(\core.registers[25][29] ),
    .S(net1419),
    .X(_07181_));
 sky130_fd_sc_hd__o21ai_1 _12269_ (.A1(net1875),
    .A2(_07181_),
    .B1(_07180_),
    .Y(_07182_));
 sky130_fd_sc_hd__o21a_1 _12270_ (.A1(\core.registers[8][29] ),
    .A2(net1421),
    .B1(net1713),
    .X(_07183_));
 sky130_fd_sc_hd__o21ai_1 _12271_ (.A1(\core.registers[9][29] ),
    .A2(net1376),
    .B1(_07183_),
    .Y(_07184_));
 sky130_fd_sc_hd__a22o_1 _12272_ (.A1(net1698),
    .A2(\core.registers[10][29] ),
    .B1(\core.registers[11][29] ),
    .B2(net1421),
    .X(_07185_));
 sky130_fd_sc_hd__a21oi_1 _12273_ (.A1(net1875),
    .A2(_07185_),
    .B1(net1858),
    .Y(_07186_));
 sky130_fd_sc_hd__a221o_1 _12274_ (.A1(net1858),
    .A2(_07182_),
    .B1(_07184_),
    .B2(_07186_),
    .C1(net1864),
    .X(_07187_));
 sky130_fd_sc_hd__or3b_4 _12275_ (.A(net1487),
    .B(_07179_),
    .C_N(_07187_),
    .X(_07188_));
 sky130_fd_sc_hd__o21a_2 _12276_ (.A1(net1491),
    .A2(_07171_),
    .B1(_07188_),
    .X(_07189_));
 sky130_fd_sc_hd__a22o_4 _12277_ (.A1(net1070),
    .A2(net1095),
    .B1(_07189_),
    .B2(net1066),
    .X(_07190_));
 sky130_fd_sc_hd__mux2_8 _12278_ (.A0(net471),
    .A1(_07190_),
    .S(net1277),
    .X(_07191_));
 sky130_fd_sc_hd__clkinv_2 _12279_ (.A(_07191_),
    .Y(_07192_));
 sky130_fd_sc_hd__nor2_4 _12280_ (.A(_07160_),
    .B(_07191_),
    .Y(_07193_));
 sky130_fd_sc_hd__inv_2 _12281_ (.A(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__and2_4 _12282_ (.A(_07160_),
    .B(_07191_),
    .X(_07195_));
 sky130_fd_sc_hd__nor2_8 _12283_ (.A(_07193_),
    .B(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__or2_1 _12284_ (.A(_07072_),
    .B(_07109_),
    .X(_07197_));
 sky130_fd_sc_hd__a21oi_2 _12285_ (.A1(_07114_),
    .A2(_07197_),
    .B1(_07196_),
    .Y(_07198_));
 sky130_fd_sc_hd__and3_2 _12286_ (.A(_07114_),
    .B(_07196_),
    .C(_07197_),
    .X(_07199_));
 sky130_fd_sc_hd__a21oi_1 _12287_ (.A1(_07027_),
    .A2(_07118_),
    .B1(_06950_),
    .Y(_07200_));
 sky130_fd_sc_hd__and3_1 _12288_ (.A(_06950_),
    .B(_07027_),
    .C(_07118_),
    .X(_07201_));
 sky130_fd_sc_hd__o2111ai_4 _12289_ (.A1(_07198_),
    .A2(_07199_),
    .B1(_06661_),
    .C1(_06796_),
    .D1(_07120_),
    .Y(_07202_));
 sky130_fd_sc_hd__or4_2 _12290_ (.A(_06873_),
    .B(_07116_),
    .C(_07200_),
    .D(_07201_),
    .X(_07203_));
 sky130_fd_sc_hd__a22o_1 _12291_ (.A1(\core.pipe1_resultRegister[31] ),
    .A2(net1240),
    .B1(net1268),
    .B2(\core.pipe1_csrData[31] ),
    .X(_07204_));
 sky130_fd_sc_hd__a31o_1 _12292_ (.A1(_04566_),
    .A2(_04571_),
    .A3(net1233),
    .B1(net2014),
    .X(_07205_));
 sky130_fd_sc_hd__a21o_2 _12293_ (.A1(net1189),
    .A2(_07205_),
    .B1(_07204_),
    .X(_07206_));
 sky130_fd_sc_hd__or2_1 _12294_ (.A(\core.registers[6][31] ),
    .B(net1563),
    .X(_07207_));
 sky130_fd_sc_hd__or2_1 _12295_ (.A(\core.registers[17][31] ),
    .B(net1501),
    .X(_07208_));
 sky130_fd_sc_hd__mux2_1 _12296_ (.A0(\core.registers[28][31] ),
    .A1(\core.registers[29][31] ),
    .S(net1557),
    .X(_07209_));
 sky130_fd_sc_hd__a221o_1 _12297_ (.A1(net1732),
    .A2(\core.registers[30][31] ),
    .B1(\core.registers[31][31] ),
    .B2(net1557),
    .C1(net1741),
    .X(_07210_));
 sky130_fd_sc_hd__o21a_1 _12298_ (.A1(net1847),
    .A2(_07209_),
    .B1(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__mux2_1 _12299_ (.A0(\core.registers[14][31] ),
    .A1(\core.registers[15][31] ),
    .S(net1558),
    .X(_07212_));
 sky130_fd_sc_hd__mux2_1 _12300_ (.A0(\core.registers[12][31] ),
    .A1(\core.registers[13][31] ),
    .S(net1558),
    .X(_07213_));
 sky130_fd_sc_hd__mux2_1 _12301_ (.A0(_07212_),
    .A1(_07213_),
    .S(net1609),
    .X(_07214_));
 sky130_fd_sc_hd__mux2_1 _12302_ (.A0(_07211_),
    .A1(_07214_),
    .S(net1751),
    .X(_07215_));
 sky130_fd_sc_hd__or2_1 _12303_ (.A(\core.registers[24][31] ),
    .B(net1560),
    .X(_07216_));
 sky130_fd_sc_hd__o211a_1 _12304_ (.A1(\core.registers[25][31] ),
    .A2(net1501),
    .B1(_07216_),
    .C1(net1741),
    .X(_07217_));
 sky130_fd_sc_hd__a31o_1 _12305_ (.A1(net1847),
    .A2(net1731),
    .A3(\core.registers[26][31] ),
    .B1(net1751),
    .X(_07218_));
 sky130_fd_sc_hd__a31o_1 _12306_ (.A1(net1847),
    .A2(\core.registers[27][31] ),
    .A3(net1558),
    .B1(_07218_),
    .X(_07219_));
 sky130_fd_sc_hd__mux2_1 _12307_ (.A0(\core.registers[8][31] ),
    .A1(\core.registers[9][31] ),
    .S(net1560),
    .X(_07220_));
 sky130_fd_sc_hd__mux2_1 _12308_ (.A0(\core.registers[10][31] ),
    .A1(\core.registers[11][31] ),
    .S(net1560),
    .X(_07221_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(_07220_),
    .A1(_07221_),
    .S(net1627),
    .X(_07222_));
 sky130_fd_sc_hd__o221a_1 _12310_ (.A1(_07217_),
    .A2(_07219_),
    .B1(_07222_),
    .B2(net1827),
    .C1(net1747),
    .X(_07223_));
 sky130_fd_sc_hd__a211o_2 _12311_ (.A1(net1835),
    .A2(_07215_),
    .B1(_07223_),
    .C1(net1633),
    .X(_07224_));
 sky130_fd_sc_hd__o211a_1 _12312_ (.A1(net1734),
    .A2(\core.registers[7][31] ),
    .B1(net1627),
    .C1(_07207_),
    .X(_07225_));
 sky130_fd_sc_hd__mux2_1 _12313_ (.A0(\core.registers[4][31] ),
    .A1(\core.registers[5][31] ),
    .S(net1563),
    .X(_07226_));
 sky130_fd_sc_hd__a211o_1 _12314_ (.A1(net1608),
    .A2(_07226_),
    .B1(_07225_),
    .C1(net1582),
    .X(_07227_));
 sky130_fd_sc_hd__mux2_1 _12315_ (.A0(\core.registers[0][31] ),
    .A1(\core.registers[1][31] ),
    .S(net1562),
    .X(_07228_));
 sky130_fd_sc_hd__mux2_1 _12316_ (.A0(\core.registers[2][31] ),
    .A1(\core.registers[3][31] ),
    .S(net1562),
    .X(_07229_));
 sky130_fd_sc_hd__mux2_1 _12317_ (.A0(_07228_),
    .A1(_07229_),
    .S(net1628),
    .X(_07230_));
 sky130_fd_sc_hd__o211a_2 _12318_ (.A1(net1593),
    .A2(_07230_),
    .B1(_07227_),
    .C1(net1569),
    .X(_07231_));
 sky130_fd_sc_hd__o211a_1 _12319_ (.A1(\core.registers[16][31] ),
    .A2(net1561),
    .B1(_07208_),
    .C1(net1607),
    .X(_07232_));
 sky130_fd_sc_hd__mux2_1 _12320_ (.A0(\core.registers[18][31] ),
    .A1(\core.registers[19][31] ),
    .S(net1561),
    .X(_07233_));
 sky130_fd_sc_hd__a211o_1 _12321_ (.A1(net1627),
    .A2(_07233_),
    .B1(_07232_),
    .C1(net1592),
    .X(_07234_));
 sky130_fd_sc_hd__mux2_1 _12322_ (.A0(\core.registers[22][31] ),
    .A1(\core.registers[23][31] ),
    .S(net1561),
    .X(_07235_));
 sky130_fd_sc_hd__mux2_1 _12323_ (.A0(\core.registers[20][31] ),
    .A1(\core.registers[21][31] ),
    .S(net1561),
    .X(_07236_));
 sky130_fd_sc_hd__mux2_1 _12324_ (.A0(_07235_),
    .A1(_07236_),
    .S(net1607),
    .X(_07237_));
 sky130_fd_sc_hd__o211a_1 _12325_ (.A1(net1581),
    .A2(_07237_),
    .B1(_07234_),
    .C1(net1574),
    .X(_07238_));
 sky130_fd_sc_hd__o31a_4 _12326_ (.A1(net1638),
    .A2(_07231_),
    .A3(_07238_),
    .B1(_07224_),
    .X(_07239_));
 sky130_fd_sc_hd__o21a_1 _12327_ (.A1(net1156),
    .A2(net1091),
    .B1(net1265),
    .X(_07240_));
 sky130_fd_sc_hd__o21ai_4 _12328_ (.A1(net1159),
    .A2(_07239_),
    .B1(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__a21oi_1 _12329_ (.A1(net1279),
    .A2(_04484_),
    .B1(net1815),
    .Y(_07242_));
 sky130_fd_sc_hd__a31o_1 _12330_ (.A1(net1279),
    .A2(_04484_),
    .A3(_07241_),
    .B1(_07242_),
    .X(_07243_));
 sky130_fd_sc_hd__o22a_1 _12331_ (.A1(net1699),
    .A2(\core.registers[23][31] ),
    .B1(net1427),
    .B2(\core.registers[22][31] ),
    .X(_07244_));
 sky130_fd_sc_hd__or3_1 _12332_ (.A(net1699),
    .B(\core.registers[19][31] ),
    .C(net1455),
    .X(_07245_));
 sky130_fd_sc_hd__o221a_1 _12333_ (.A1(\core.registers[18][31] ),
    .A2(net1335),
    .B1(_07244_),
    .B2(net1440),
    .C1(_07245_),
    .X(_07246_));
 sky130_fd_sc_hd__mux4_1 _12334_ (.A0(\core.registers[16][31] ),
    .A1(\core.registers[17][31] ),
    .A2(\core.registers[20][31] ),
    .A3(\core.registers[21][31] ),
    .S0(net1427),
    .S1(net1456),
    .X(_07247_));
 sky130_fd_sc_hd__mux2_1 _12335_ (.A0(_07246_),
    .A1(_07247_),
    .S(net1475),
    .X(_07248_));
 sky130_fd_sc_hd__o22a_1 _12336_ (.A1(net1700),
    .A2(\core.registers[7][31] ),
    .B1(net1428),
    .B2(\core.registers[6][31] ),
    .X(_07249_));
 sky130_fd_sc_hd__or3_1 _12337_ (.A(net1700),
    .B(\core.registers[3][31] ),
    .C(net1457),
    .X(_07250_));
 sky130_fd_sc_hd__o221a_1 _12338_ (.A1(\core.registers[2][31] ),
    .A2(net1335),
    .B1(_07249_),
    .B2(net1440),
    .C1(_07250_),
    .X(_07251_));
 sky130_fd_sc_hd__mux4_1 _12339_ (.A0(\core.registers[0][31] ),
    .A1(\core.registers[1][31] ),
    .A2(\core.registers[4][31] ),
    .A3(\core.registers[5][31] ),
    .S0(net1428),
    .S1(net1458),
    .X(_07252_));
 sky130_fd_sc_hd__mux2_2 _12340_ (.A0(_07251_),
    .A1(_07252_),
    .S(net1475),
    .X(_07253_));
 sky130_fd_sc_hd__mux2_2 _12341_ (.A0(_07248_),
    .A1(_07253_),
    .S(net1463),
    .X(_07254_));
 sky130_fd_sc_hd__nor2_1 _12342_ (.A(net1492),
    .B(_07254_),
    .Y(_07255_));
 sky130_fd_sc_hd__mux2_1 _12343_ (.A0(\core.registers[14][31] ),
    .A1(\core.registers[15][31] ),
    .S(net1423),
    .X(_07256_));
 sky130_fd_sc_hd__mux2_1 _12344_ (.A0(\core.registers[12][31] ),
    .A1(\core.registers[13][31] ),
    .S(net1424),
    .X(_07257_));
 sky130_fd_sc_hd__mux2_1 _12345_ (.A0(_07256_),
    .A1(_07257_),
    .S(net1474),
    .X(_07258_));
 sky130_fd_sc_hd__mux2_1 _12346_ (.A0(\core.registers[28][31] ),
    .A1(\core.registers[29][31] ),
    .S(net1423),
    .X(_07259_));
 sky130_fd_sc_hd__a221o_1 _12347_ (.A1(net1696),
    .A2(\core.registers[30][31] ),
    .B1(\core.registers[31][31] ),
    .B2(net1423),
    .C1(net1712),
    .X(_07260_));
 sky130_fd_sc_hd__o21ai_1 _12348_ (.A1(net1876),
    .A2(_07259_),
    .B1(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__o21ai_1 _12349_ (.A1(net1859),
    .A2(_07258_),
    .B1(net1865),
    .Y(_07262_));
 sky130_fd_sc_hd__a21o_1 _12350_ (.A1(net1860),
    .A2(_07261_),
    .B1(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__a221o_1 _12351_ (.A1(net1699),
    .A2(\core.registers[26][31] ),
    .B1(\core.registers[27][31] ),
    .B2(net1426),
    .C1(net1711),
    .X(_07264_));
 sky130_fd_sc_hd__mux2_1 _12352_ (.A0(\core.registers[24][31] ),
    .A1(\core.registers[25][31] ),
    .S(net1426),
    .X(_07265_));
 sky130_fd_sc_hd__o21ai_1 _12353_ (.A1(net1876),
    .A2(_07265_),
    .B1(_07264_),
    .Y(_07266_));
 sky130_fd_sc_hd__o21a_1 _12354_ (.A1(\core.registers[8][31] ),
    .A2(net1426),
    .B1(net1711),
    .X(_07267_));
 sky130_fd_sc_hd__o21ai_1 _12355_ (.A1(\core.registers[9][31] ),
    .A2(net1378),
    .B1(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__a22o_1 _12356_ (.A1(net1697),
    .A2(\core.registers[10][31] ),
    .B1(\core.registers[11][31] ),
    .B2(net1426),
    .X(_07269_));
 sky130_fd_sc_hd__a21oi_1 _12357_ (.A1(net1876),
    .A2(_07269_),
    .B1(net1859),
    .Y(_07270_));
 sky130_fd_sc_hd__a221o_1 _12358_ (.A1(net1859),
    .A2(_07266_),
    .B1(_07268_),
    .B2(_07270_),
    .C1(net1864),
    .X(_07271_));
 sky130_fd_sc_hd__a31o_4 _12359_ (.A1(net1491),
    .A2(_07263_),
    .A3(_07271_),
    .B1(_07255_),
    .X(_07272_));
 sky130_fd_sc_hd__o2bb2a_4 _12360_ (.A1_N(net1071),
    .A2_N(net1091),
    .B1(_07272_),
    .B2(_04663_),
    .X(_07273_));
 sky130_fd_sc_hd__inv_2 _12361_ (.A(_07273_),
    .Y(_07274_));
 sky130_fd_sc_hd__mux2_8 _12362_ (.A0(net474),
    .A1(_07274_),
    .S(net1277),
    .X(_07275_));
 sky130_fd_sc_hd__or2_2 _12363_ (.A(_07243_),
    .B(_07275_),
    .X(_07276_));
 sky130_fd_sc_hd__inv_2 _12364_ (.A(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__a22o_1 _12365_ (.A1(\core.pipe1_resultRegister[30] ),
    .A2(net1240),
    .B1(net1268),
    .B2(\core.pipe1_csrData[30] ),
    .X(_07278_));
 sky130_fd_sc_hd__a21o_1 _12366_ (.A1(net1235),
    .A2(_05202_),
    .B1(net1237),
    .X(_07279_));
 sky130_fd_sc_hd__a21o_2 _12367_ (.A1(net1190),
    .A2(_07279_),
    .B1(_07278_),
    .X(_07280_));
 sky130_fd_sc_hd__mux2_1 _12368_ (.A0(\core.registers[24][30] ),
    .A1(\core.registers[25][30] ),
    .S(net1548),
    .X(_07281_));
 sky130_fd_sc_hd__a221o_1 _12369_ (.A1(net1731),
    .A2(\core.registers[26][30] ),
    .B1(\core.registers[27][30] ),
    .B2(net1548),
    .C1(net1740),
    .X(_07282_));
 sky130_fd_sc_hd__o21ai_1 _12370_ (.A1(net1845),
    .A2(_07281_),
    .B1(_07282_),
    .Y(_07283_));
 sky130_fd_sc_hd__a221o_1 _12371_ (.A1(net1732),
    .A2(\core.registers[30][30] ),
    .B1(\core.registers[31][30] ),
    .B2(net1547),
    .C1(net1740),
    .X(_07284_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(\core.registers[28][30] ),
    .A1(\core.registers[29][30] ),
    .S(net1547),
    .X(_07285_));
 sky130_fd_sc_hd__o21a_1 _12373_ (.A1(net1844),
    .A2(_07285_),
    .B1(_07284_),
    .X(_07286_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(\core.registers[12][30] ),
    .A1(\core.registers[13][30] ),
    .S(net1547),
    .X(_07287_));
 sky130_fd_sc_hd__mux2_1 _12375_ (.A0(\core.registers[14][30] ),
    .A1(\core.registers[15][30] ),
    .S(net1547),
    .X(_07288_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(_07287_),
    .A1(_07288_),
    .S(net1626),
    .X(_07289_));
 sky130_fd_sc_hd__mux2_1 _12377_ (.A0(_07286_),
    .A1(_07289_),
    .S(net1750),
    .X(_07290_));
 sky130_fd_sc_hd__or2_1 _12378_ (.A(\core.registers[6][30] ),
    .B(net1553),
    .X(_07291_));
 sky130_fd_sc_hd__or2_1 _12379_ (.A(\core.registers[22][30] ),
    .B(net1553),
    .X(_07292_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(\core.registers[8][30] ),
    .A1(\core.registers[9][30] ),
    .S(net1551),
    .X(_07293_));
 sky130_fd_sc_hd__mux2_1 _12381_ (.A0(\core.registers[10][30] ),
    .A1(\core.registers[11][30] ),
    .S(net1551),
    .X(_07294_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(_07293_),
    .A1(_07294_),
    .S(net1624),
    .X(_07295_));
 sky130_fd_sc_hd__or2_1 _12383_ (.A(net1826),
    .B(_07295_),
    .X(_07296_));
 sky130_fd_sc_hd__a21oi_1 _12384_ (.A1(net1826),
    .A2(_07283_),
    .B1(net1834),
    .Y(_07297_));
 sky130_fd_sc_hd__a221o_2 _12385_ (.A1(net1834),
    .A2(_07290_),
    .B1(_07296_),
    .B2(_07297_),
    .C1(net1634),
    .X(_07298_));
 sky130_fd_sc_hd__o211a_1 _12386_ (.A1(net1731),
    .A2(\core.registers[7][30] ),
    .B1(net1624),
    .C1(_07291_),
    .X(_07299_));
 sky130_fd_sc_hd__mux2_1 _12387_ (.A0(\core.registers[4][30] ),
    .A1(\core.registers[5][30] ),
    .S(net1560),
    .X(_07300_));
 sky130_fd_sc_hd__a211o_1 _12388_ (.A1(net1610),
    .A2(_07300_),
    .B1(_07299_),
    .C1(net1581),
    .X(_07301_));
 sky130_fd_sc_hd__mux2_1 _12389_ (.A0(\core.registers[0][30] ),
    .A1(\core.registers[1][30] ),
    .S(net1560),
    .X(_07302_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(\core.registers[2][30] ),
    .A1(\core.registers[3][30] ),
    .S(net1553),
    .X(_07303_));
 sky130_fd_sc_hd__mux2_1 _12391_ (.A0(_07302_),
    .A1(_07303_),
    .S(net1624),
    .X(_07304_));
 sky130_fd_sc_hd__o211a_1 _12392_ (.A1(net1592),
    .A2(_07304_),
    .B1(_07301_),
    .C1(net1570),
    .X(_07305_));
 sky130_fd_sc_hd__mux2_1 _12393_ (.A0(\core.registers[16][30] ),
    .A1(\core.registers[17][30] ),
    .S(net1553),
    .X(_07306_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(\core.registers[18][30] ),
    .A1(\core.registers[19][30] ),
    .S(net1553),
    .X(_07307_));
 sky130_fd_sc_hd__mux2_1 _12395_ (.A0(_07306_),
    .A1(_07307_),
    .S(net1625),
    .X(_07308_));
 sky130_fd_sc_hd__o211a_1 _12396_ (.A1(net1731),
    .A2(\core.registers[23][30] ),
    .B1(net1625),
    .C1(_07292_),
    .X(_07309_));
 sky130_fd_sc_hd__mux2_1 _12397_ (.A0(\core.registers[20][30] ),
    .A1(\core.registers[21][30] ),
    .S(net1553),
    .X(_07310_));
 sky130_fd_sc_hd__a211o_1 _12398_ (.A1(net1610),
    .A2(_07310_),
    .B1(_07309_),
    .C1(net1581),
    .X(_07311_));
 sky130_fd_sc_hd__o211a_1 _12399_ (.A1(net1592),
    .A2(_07308_),
    .B1(_07311_),
    .C1(net1574),
    .X(_07312_));
 sky130_fd_sc_hd__o31a_4 _12400_ (.A1(net1638),
    .A2(_07305_),
    .A3(_07312_),
    .B1(_07298_),
    .X(_07313_));
 sky130_fd_sc_hd__o21a_1 _12401_ (.A1(net1160),
    .A2(_07313_),
    .B1(net1265),
    .X(_07314_));
 sky130_fd_sc_hd__o21ai_4 _12402_ (.A1(net1156),
    .A2(net1087),
    .B1(_07314_),
    .Y(_07315_));
 sky130_fd_sc_hd__o21ai_1 _12403_ (.A1(net1193),
    .A2(_07315_),
    .B1(net1162),
    .Y(_07316_));
 sky130_fd_sc_hd__o21a_1 _12404_ (.A1(net1817),
    .A2(net1279),
    .B1(_07316_),
    .X(_07317_));
 sky130_fd_sc_hd__o22a_1 _12405_ (.A1(net1697),
    .A2(\core.registers[23][30] ),
    .B1(net1420),
    .B2(\core.registers[22][30] ),
    .X(_07318_));
 sky130_fd_sc_hd__or3_1 _12406_ (.A(net1697),
    .B(\core.registers[19][30] ),
    .C(net1455),
    .X(_07319_));
 sky130_fd_sc_hd__o221a_1 _12407_ (.A1(\core.registers[18][30] ),
    .A2(net1335),
    .B1(_07318_),
    .B2(net1441),
    .C1(_07319_),
    .X(_07320_));
 sky130_fd_sc_hd__mux4_1 _12408_ (.A0(\core.registers[16][30] ),
    .A1(\core.registers[17][30] ),
    .A2(\core.registers[20][30] ),
    .A3(\core.registers[21][30] ),
    .S0(net1420),
    .S1(net1455),
    .X(_07321_));
 sky130_fd_sc_hd__mux2_1 _12409_ (.A0(_07320_),
    .A1(_07321_),
    .S(net1476),
    .X(_07322_));
 sky130_fd_sc_hd__o22a_1 _12410_ (.A1(net1697),
    .A2(\core.registers[7][30] ),
    .B1(net1420),
    .B2(\core.registers[6][30] ),
    .X(_07323_));
 sky130_fd_sc_hd__or3_1 _12411_ (.A(net1697),
    .B(\core.registers[3][30] ),
    .C(net1456),
    .X(_07324_));
 sky130_fd_sc_hd__o221a_1 _12412_ (.A1(\core.registers[2][30] ),
    .A2(net1335),
    .B1(_07323_),
    .B2(net1441),
    .C1(_07324_),
    .X(_07325_));
 sky130_fd_sc_hd__mux4_1 _12413_ (.A0(\core.registers[0][30] ),
    .A1(\core.registers[1][30] ),
    .A2(\core.registers[4][30] ),
    .A3(\core.registers[5][30] ),
    .S0(net1426),
    .S1(net1456),
    .X(_07326_));
 sky130_fd_sc_hd__mux2_1 _12414_ (.A0(_07325_),
    .A1(_07326_),
    .S(net1476),
    .X(_07327_));
 sky130_fd_sc_hd__mux2_2 _12415_ (.A0(_07322_),
    .A1(_07327_),
    .S(net1463),
    .X(_07328_));
 sky130_fd_sc_hd__a221o_1 _12416_ (.A1(net1695),
    .A2(\core.registers[26][30] ),
    .B1(\core.registers[27][30] ),
    .B2(net1416),
    .C1(net1709),
    .X(_07329_));
 sky130_fd_sc_hd__mux2_1 _12417_ (.A0(\core.registers[24][30] ),
    .A1(\core.registers[25][30] ),
    .S(net1416),
    .X(_07330_));
 sky130_fd_sc_hd__o21ai_1 _12418_ (.A1(net1875),
    .A2(_07330_),
    .B1(_07329_),
    .Y(_07331_));
 sky130_fd_sc_hd__a221o_1 _12419_ (.A1(net1698),
    .A2(\core.registers[10][30] ),
    .B1(\core.registers[11][30] ),
    .B2(net1419),
    .C1(net1709),
    .X(_07332_));
 sky130_fd_sc_hd__a21o_1 _12420_ (.A1(\core.registers[8][30] ),
    .A2(net1376),
    .B1(net1875),
    .X(_07333_));
 sky130_fd_sc_hd__a21o_1 _12421_ (.A1(\core.registers[9][30] ),
    .A2(net1419),
    .B1(_07333_),
    .X(_07334_));
 sky130_fd_sc_hd__a21oi_1 _12422_ (.A1(_07332_),
    .A2(_07334_),
    .B1(net1859),
    .Y(_07335_));
 sky130_fd_sc_hd__a211o_1 _12423_ (.A1(net1859),
    .A2(_07331_),
    .B1(_07335_),
    .C1(net1864),
    .X(_07336_));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(\core.registers[12][30] ),
    .A1(\core.registers[13][30] ),
    .S(net1415),
    .X(_07337_));
 sky130_fd_sc_hd__mux2_1 _12425_ (.A0(\core.registers[14][30] ),
    .A1(\core.registers[15][30] ),
    .S(net1415),
    .X(_07338_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(_07337_),
    .A1(_07338_),
    .S(net1483),
    .X(_07339_));
 sky130_fd_sc_hd__a221o_1 _12427_ (.A1(net1695),
    .A2(\core.registers[30][30] ),
    .B1(\core.registers[31][30] ),
    .B2(net1415),
    .C1(net1710),
    .X(_07340_));
 sky130_fd_sc_hd__mux2_1 _12428_ (.A0(\core.registers[28][30] ),
    .A1(\core.registers[29][30] ),
    .S(net1415),
    .X(_07341_));
 sky130_fd_sc_hd__o21a_1 _12429_ (.A1(net1874),
    .A2(_07341_),
    .B1(_07340_),
    .X(_07342_));
 sky130_fd_sc_hd__mux2_1 _12430_ (.A0(_07339_),
    .A1(_07342_),
    .S(net1857),
    .X(_07343_));
 sky130_fd_sc_hd__a21oi_2 _12431_ (.A1(net1864),
    .A2(_07343_),
    .B1(net1487),
    .Y(_07344_));
 sky130_fd_sc_hd__o2bb2a_4 _12432_ (.A1_N(_07336_),
    .A2_N(_07344_),
    .B1(net1491),
    .B2(_07328_),
    .X(_07345_));
 sky130_fd_sc_hd__a22o_4 _12433_ (.A1(net1071),
    .A2(net1087),
    .B1(_07345_),
    .B2(net1066),
    .X(_07346_));
 sky130_fd_sc_hd__mux2_8 _12434_ (.A0(net473),
    .A1(_07346_),
    .S(net1276),
    .X(_07347_));
 sky130_fd_sc_hd__nor2_2 _12435_ (.A(_07317_),
    .B(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__and2_4 _12436_ (.A(_07317_),
    .B(_07347_),
    .X(_07349_));
 sky130_fd_sc_hd__nor2_8 _12437_ (.A(_07348_),
    .B(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__inv_2 _12438_ (.A(_07350_),
    .Y(_07351_));
 sky130_fd_sc_hd__a2111o_4 _12439_ (.A1(_07026_),
    .A2(_07032_),
    .B1(_07113_),
    .C1(_07196_),
    .D1(_07350_),
    .X(_07352_));
 sky130_fd_sc_hd__and2_2 _12440_ (.A(_07243_),
    .B(_07275_),
    .X(_07353_));
 sky130_fd_sc_hd__o32a_1 _12441_ (.A1(_07072_),
    .A2(_07109_),
    .A3(_07196_),
    .B1(_07192_),
    .B2(_07160_),
    .X(_07354_));
 sky130_fd_sc_hd__or2_1 _12442_ (.A(_07350_),
    .B(_07354_),
    .X(_07355_));
 sky130_fd_sc_hd__nand2b_1 _12443_ (.A_N(_07317_),
    .B(_07347_),
    .Y(_07356_));
 sky130_fd_sc_hd__and2_1 _12444_ (.A(_07355_),
    .B(_07356_),
    .X(_07357_));
 sky130_fd_sc_hd__nand2b_1 _12445_ (.A_N(_07353_),
    .B(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__inv_2 _12446_ (.A(_07358_),
    .Y(_07359_));
 sky130_fd_sc_hd__nor2_4 _12447_ (.A(_07277_),
    .B(_07353_),
    .Y(_07360_));
 sky130_fd_sc_hd__a21o_1 _12448_ (.A1(_07352_),
    .A2(_07359_),
    .B1(_07277_),
    .X(_07361_));
 sky130_fd_sc_hd__and3_1 _12449_ (.A(_07276_),
    .B(_07352_),
    .C(_07359_),
    .X(_07362_));
 sky130_fd_sc_hd__and2_1 _12450_ (.A(_07352_),
    .B(_07355_),
    .X(_07363_));
 sky130_fd_sc_hd__a21oi_1 _12451_ (.A1(_07352_),
    .A2(_07357_),
    .B1(_07360_),
    .Y(_07364_));
 sky130_fd_sc_hd__o211ai_2 _12452_ (.A1(_07114_),
    .A2(_07196_),
    .B1(_07350_),
    .C1(_07354_),
    .Y(_07365_));
 sky130_fd_sc_hd__a211o_1 _12453_ (.A1(_07363_),
    .A2(_07365_),
    .B1(_07364_),
    .C1(_07362_),
    .X(_07366_));
 sky130_fd_sc_hd__nor3_1 _12454_ (.A(_07202_),
    .B(_07203_),
    .C(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__o21ai_4 _12455_ (.A1(net1880),
    .A2(net1882),
    .B1(net1665),
    .Y(_07368_));
 sky130_fd_sc_hd__o21a_4 _12456_ (.A1(net1880),
    .A2(net1881),
    .B1(net1666),
    .X(_07369_));
 sky130_fd_sc_hd__nand2_2 _12457_ (.A(net1878),
    .B(net1666),
    .Y(_07370_));
 sky130_fd_sc_hd__and2_1 _12458_ (.A(net1372),
    .B(_07370_),
    .X(_07371_));
 sky130_fd_sc_hd__nand2_1 _12459_ (.A(net1372),
    .B(_07370_),
    .Y(_07372_));
 sky130_fd_sc_hd__a31o_1 _12460_ (.A1(_07276_),
    .A2(_07352_),
    .A3(_07357_),
    .B1(_07353_),
    .X(_07373_));
 sky130_fd_sc_hd__nor2_8 _12461_ (.A(_04423_),
    .B(_04477_),
    .Y(_07374_));
 sky130_fd_sc_hd__nand2_1 _12462_ (.A(net1878),
    .B(_04476_),
    .Y(_07375_));
 sky130_fd_sc_hd__nor2_1 _12463_ (.A(_07373_),
    .B(net1325),
    .Y(_07376_));
 sky130_fd_sc_hd__and3_4 _12464_ (.A(net1880),
    .B(net1881),
    .C(net1666),
    .X(_07377_));
 sky130_fd_sc_hd__and2_4 _12465_ (.A(net1878),
    .B(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__nand2_8 _12466_ (.A(net1878),
    .B(_07377_),
    .Y(_07379_));
 sky130_fd_sc_hd__nor3_4 _12467_ (.A(_04423_),
    .B(net1881),
    .C(_04463_),
    .Y(_07380_));
 sky130_fd_sc_hd__or3_4 _12468_ (.A(_04423_),
    .B(net1881),
    .C(_04463_),
    .X(_07381_));
 sky130_fd_sc_hd__mux2_1 _12469_ (.A0(net1321),
    .A1(net1318),
    .S(_07361_),
    .X(_07382_));
 sky130_fd_sc_hd__nor2_4 _12470_ (.A(_07369_),
    .B(_07370_),
    .Y(_07383_));
 sky130_fd_sc_hd__or2_4 _12471_ (.A(_07369_),
    .B(_07370_),
    .X(_07384_));
 sky130_fd_sc_hd__a211o_1 _12472_ (.A1(_07373_),
    .A2(net1316),
    .B1(_07382_),
    .C1(_07376_),
    .X(_07385_));
 sky130_fd_sc_hd__nor2_4 _12473_ (.A(net1878),
    .B(_04477_),
    .Y(_07386_));
 sky130_fd_sc_hd__nand2_1 _12474_ (.A(_04423_),
    .B(_04476_),
    .Y(_07387_));
 sky130_fd_sc_hd__o31a_1 _12475_ (.A1(_07202_),
    .A2(_07203_),
    .A3(_07366_),
    .B1(net1313),
    .X(_07388_));
 sky130_fd_sc_hd__a211o_1 _12476_ (.A1(_07367_),
    .A2(net1330),
    .B1(_07385_),
    .C1(_07388_),
    .X(_07389_));
 sky130_fd_sc_hd__o211a_1 _12477_ (.A1(net1878),
    .A2(_04463_),
    .B1(_04461_),
    .C1(_04449_),
    .X(_07390_));
 sky130_fd_sc_hd__inv_2 _12478_ (.A(net1260),
    .Y(_07391_));
 sky130_fd_sc_hd__and2_2 _12479_ (.A(net801),
    .B(net1260),
    .X(_07392_));
 sky130_fd_sc_hd__and3_4 _12480_ (.A(_04449_),
    .B(_04451_),
    .C(_04455_),
    .X(_07393_));
 sky130_fd_sc_hd__and2_4 _12481_ (.A(net1329),
    .B(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__nand2_1 _12482_ (.A(net1329),
    .B(_07393_),
    .Y(_07395_));
 sky130_fd_sc_hd__a21oi_4 _12483_ (.A1(net2015),
    .A2(net1259),
    .B1(net1229),
    .Y(_07396_));
 sky130_fd_sc_hd__a21o_2 _12484_ (.A1(net2015),
    .A2(net1259),
    .B1(net1229),
    .X(_07397_));
 sky130_fd_sc_hd__nor2_1 _12485_ (.A(net1295),
    .B(net1230),
    .Y(_07398_));
 sky130_fd_sc_hd__nand2_8 _12486_ (.A(net1290),
    .B(net1226),
    .Y(_07399_));
 sky130_fd_sc_hd__a21oi_4 _12487_ (.A1(net799),
    .A2(net1259),
    .B1(net1183),
    .Y(_07400_));
 sky130_fd_sc_hd__a21o_4 _12488_ (.A1(net799),
    .A2(net1259),
    .B1(net1182),
    .X(_07401_));
 sky130_fd_sc_hd__and2_4 _12489_ (.A(net1665),
    .B(_04450_),
    .X(_07402_));
 sky130_fd_sc_hd__nand2_8 _12490_ (.A(net1665),
    .B(_04450_),
    .Y(_07403_));
 sky130_fd_sc_hd__a32o_2 _12491_ (.A1(\core.pipe0_currentInstruction[8] ),
    .A2(net801),
    .A3(net1261),
    .B1(net1183),
    .B2(net1849),
    .X(_07404_));
 sky130_fd_sc_hd__xnor2_1 _12492_ (.A(net461),
    .B(_07402_),
    .Y(_07405_));
 sky130_fd_sc_hd__or2_2 _12493_ (.A(_07394_),
    .B(_07405_),
    .X(_07406_));
 sky130_fd_sc_hd__o21ai_4 _12494_ (.A1(_06132_),
    .A2(net1228),
    .B1(_07406_),
    .Y(_07407_));
 sky130_fd_sc_hd__nand2_1 _12495_ (.A(_07404_),
    .B(_07407_),
    .Y(_07408_));
 sky130_fd_sc_hd__xnor2_2 _12496_ (.A(_07404_),
    .B(_07407_),
    .Y(_07409_));
 sky130_fd_sc_hd__a211o_2 _12497_ (.A1(_04454_),
    .A2(_06225_),
    .B1(net1228),
    .C1(net1730),
    .X(_07410_));
 sky130_fd_sc_hd__xnor2_1 _12498_ (.A(_07409_),
    .B(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__a21oi_2 _12499_ (.A1(_07403_),
    .A2(_07411_),
    .B1(net797),
    .Y(_07412_));
 sky130_fd_sc_hd__and4_4 _12500_ (.A(\core.pipe0_currentInstruction[6] ),
    .B(\core.pipe0_currentInstruction[5] ),
    .C(\core.pipe0_currentInstruction[4] ),
    .D(_04461_),
    .X(_07413_));
 sky130_fd_sc_hd__or4_1 _12501_ (.A(\core.pipe0_currentInstruction[10] ),
    .B(\core.pipe0_currentInstruction[9] ),
    .C(\core.pipe0_currentInstruction[8] ),
    .D(\core.pipe0_currentInstruction[7] ),
    .X(_07414_));
 sky130_fd_sc_hd__or3_4 _12502_ (.A(\core.pipe0_currentInstruction[13] ),
    .B(\core.pipe0_currentInstruction[11] ),
    .C(_07414_),
    .X(_07415_));
 sky130_fd_sc_hd__or4b_4 _12503_ (.A(net1879),
    .B(_07415_),
    .C(net1882),
    .D_N(_07413_),
    .X(_07416_));
 sky130_fd_sc_hd__or3_1 _12504_ (.A(net1866),
    .B(net1873),
    .C(\core.pipe0_currentInstruction[15] ),
    .X(_07417_));
 sky130_fd_sc_hd__or4_1 _12505_ (.A(net1821),
    .B(net1822),
    .C(net1856),
    .D(\core.pipe0_currentInstruction[18] ),
    .X(_07418_));
 sky130_fd_sc_hd__or4_4 _12506_ (.A(net1829),
    .B(net1831),
    .C(_07417_),
    .D(_07418_),
    .X(_07419_));
 sky130_fd_sc_hd__or4b_1 _12507_ (.A(_04414_),
    .B(net1820),
    .C(net1837),
    .D_N(net1819),
    .X(_07420_));
 sky130_fd_sc_hd__or4b_2 _12508_ (.A(net1816),
    .B(_07420_),
    .C(net1817),
    .D_N(_04608_),
    .X(_07421_));
 sky130_fd_sc_hd__nor3_4 _12509_ (.A(_07416_),
    .B(_07419_),
    .C(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__or4b_2 _12510_ (.A(net1879),
    .B(_07415_),
    .C(net1882),
    .D_N(_07413_),
    .X(_07423_));
 sky130_fd_sc_hd__or2_2 _12511_ (.A(\core.pipe0_currentInstruction[18] ),
    .B(_07417_),
    .X(_07424_));
 sky130_fd_sc_hd__or4_1 _12512_ (.A(net1816),
    .B(net1818),
    .C(_04414_),
    .D(net1837),
    .X(_07425_));
 sky130_fd_sc_hd__or4_1 _12513_ (.A(net1821),
    .B(net1822),
    .C(net1829),
    .D(net1831),
    .X(_07426_));
 sky130_fd_sc_hd__or4_1 _12514_ (.A(net1743),
    .B(net1851),
    .C(net1856),
    .D(_07426_),
    .X(_07427_));
 sky130_fd_sc_hd__or4b_2 _12515_ (.A(net1820),
    .B(_07425_),
    .C(_07427_),
    .D_N(net1819),
    .X(_07428_));
 sky130_fd_sc_hd__nor3_4 _12516_ (.A(_07423_),
    .B(_07424_),
    .C(_07428_),
    .Y(_07429_));
 sky130_fd_sc_hd__or3_1 _12517_ (.A(net1816),
    .B(net1817),
    .C(_04414_),
    .X(_07430_));
 sky130_fd_sc_hd__or4b_1 _12518_ (.A(net1851),
    .B(net1861),
    .C(_07430_),
    .D_N(net1819),
    .X(_07431_));
 sky130_fd_sc_hd__or4_1 _12519_ (.A(net1820),
    .B(net1837),
    .C(net1743),
    .D(_07424_),
    .X(_07432_));
 sky130_fd_sc_hd__or4_4 _12520_ (.A(_07416_),
    .B(_07426_),
    .C(_07431_),
    .D(_07432_),
    .X(_07433_));
 sky130_fd_sc_hd__a211oi_2 _12521_ (.A1(\core.fetchProgramCounter[1] ),
    .A2(net797),
    .B1(_07412_),
    .C1(net1180),
    .Y(_07434_));
 sky130_fd_sc_hd__nor2_1 _12522_ (.A(\core.csr.trapReturnVector[1] ),
    .B(_07433_),
    .Y(_07435_));
 sky130_fd_sc_hd__o31a_2 _12523_ (.A1(net782),
    .A2(_07434_),
    .A3(_07435_),
    .B1(net1774),
    .X(_07436_));
 sky130_fd_sc_hd__a211oi_4 _12524_ (.A1(net1762),
    .A2(_04412_),
    .B1(net1980),
    .C1(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__nor2_8 _12525_ (.A(net793),
    .B(_07422_),
    .Y(_07438_));
 sky130_fd_sc_hd__or2_4 _12526_ (.A(net793),
    .B(_07422_),
    .X(_07439_));
 sky130_fd_sc_hd__and3_1 _12527_ (.A(\core.fetchProgramCounter[0] ),
    .B(net767),
    .C(net787),
    .X(_07440_));
 sky130_fd_sc_hd__a31o_1 _12528_ (.A1(\core.csr.trapReturnVector[0] ),
    .A2(net767),
    .A3(_07422_),
    .B1(net1762),
    .X(_07441_));
 sky130_fd_sc_hd__o21a_1 _12529_ (.A1(_07440_),
    .A2(_07441_),
    .B1(net1931),
    .X(_07442_));
 sky130_fd_sc_hd__o21a_4 _12530_ (.A1(net1774),
    .A2(\core.fetchProgramCounter[0] ),
    .B1(_07442_),
    .X(_07443_));
 sky130_fd_sc_hd__nor2_4 _12531_ (.A(\core.csr.instruction_memoryAddress[1] ),
    .B(\core.csr.instruction_memoryAddress[0] ),
    .Y(_07444_));
 sky130_fd_sc_hd__or2_1 _12532_ (.A(\core.csr.instruction_memoryAddress[1] ),
    .B(\core.csr.instruction_memoryAddress[0] ),
    .X(_07445_));
 sky130_fd_sc_hd__or2_2 _12533_ (.A(_07412_),
    .B(net1645),
    .X(_07446_));
 sky130_fd_sc_hd__and3_1 _12534_ (.A(\core.csr.traps.mie.currentValue[20] ),
    .B(net1797),
    .C(net181),
    .X(_07447_));
 sky130_fd_sc_hd__and3_1 _12535_ (.A(\core.csr.traps.mie.currentValue[23] ),
    .B(net1797),
    .C(net184),
    .X(_07448_));
 sky130_fd_sc_hd__and3_1 _12536_ (.A(\core.csr.traps.mie.currentValue[21] ),
    .B(net1797),
    .C(net182),
    .X(_07449_));
 sky130_fd_sc_hd__and3_2 _12537_ (.A(\core.csr.traps.mie.currentValue[24] ),
    .B(net1797),
    .C(net185),
    .X(_07450_));
 sky130_fd_sc_hd__and3_1 _12538_ (.A(\core.csr.traps.mie.currentValue[30] ),
    .B(net1797),
    .C(net176),
    .X(_07451_));
 sky130_fd_sc_hd__and3_1 _12539_ (.A(\core.csr.traps.mie.currentValue[27] ),
    .B(net1797),
    .C(net173),
    .X(_07452_));
 sky130_fd_sc_hd__and3_2 _12540_ (.A(\core.csr.traps.mie.currentValue[17] ),
    .B(net1798),
    .C(net178),
    .X(_07453_));
 sky130_fd_sc_hd__and3_1 _12541_ (.A(\core.csr.traps.mie.currentValue[29] ),
    .B(net1797),
    .C(net175),
    .X(_07454_));
 sky130_fd_sc_hd__and3_1 _12542_ (.A(\core.csr.traps.mie.currentValue[28] ),
    .B(net1797),
    .C(net174),
    .X(_07455_));
 sky130_fd_sc_hd__and3_4 _12543_ (.A(\core.csr.traps.mie.currentValue[16] ),
    .B(net1798),
    .C(net171),
    .X(_07456_));
 sky130_fd_sc_hd__and3_1 _12544_ (.A(\core.csr.traps.mie.currentValue[25] ),
    .B(net1798),
    .C(net186),
    .X(_07457_));
 sky130_fd_sc_hd__and3_1 _12545_ (.A(\core.csr.traps.mie.currentValue[22] ),
    .B(net1797),
    .C(net183),
    .X(_07458_));
 sky130_fd_sc_hd__and3_1 _12546_ (.A(\core.csr.traps.mie.currentValue[26] ),
    .B(net1798),
    .C(net172),
    .X(_07459_));
 sky130_fd_sc_hd__and3_1 _12547_ (.A(\core.csr.traps.mie.currentValue[31] ),
    .B(net1798),
    .C(net177),
    .X(_07460_));
 sky130_fd_sc_hd__and3_1 _12548_ (.A(\core.csr.traps.mie.currentValue[18] ),
    .B(net1798),
    .C(net179),
    .X(_07461_));
 sky130_fd_sc_hd__and3_1 _12549_ (.A(\core.csr.traps.mie.currentValue[19] ),
    .B(net1797),
    .C(net180),
    .X(_07462_));
 sky130_fd_sc_hd__or4_4 _12550_ (.A(_07447_),
    .B(_07455_),
    .C(_07457_),
    .D(_07459_),
    .X(_07463_));
 sky130_fd_sc_hd__or4_2 _12551_ (.A(_07449_),
    .B(_07451_),
    .C(_07456_),
    .D(_07458_),
    .X(_07464_));
 sky130_fd_sc_hd__or4_1 _12552_ (.A(_07450_),
    .B(_07452_),
    .C(_07453_),
    .D(_07461_),
    .X(_07465_));
 sky130_fd_sc_hd__or4_1 _12553_ (.A(_07448_),
    .B(_07454_),
    .C(_07460_),
    .D(_07462_),
    .X(_07466_));
 sky130_fd_sc_hd__or3_4 _12554_ (.A(_07464_),
    .B(_07465_),
    .C(_07466_),
    .X(_07467_));
 sky130_fd_sc_hd__nor2_8 _12555_ (.A(_07463_),
    .B(_07467_),
    .Y(_07468_));
 sky130_fd_sc_hd__or3b_1 _12556_ (.A(_07437_),
    .B(_07443_),
    .C_N(_07468_),
    .X(_07469_));
 sky130_fd_sc_hd__nor2_1 _12557_ (.A(_07446_),
    .B(_07469_),
    .Y(_07470_));
 sky130_fd_sc_hd__nand2_1 _12558_ (.A(_04465_),
    .B(net1241),
    .Y(_07471_));
 sky130_fd_sc_hd__and2_2 _12559_ (.A(_06137_),
    .B(_06695_),
    .X(_07472_));
 sky130_fd_sc_hd__nor2_4 _12560_ (.A(_06137_),
    .B(_06695_),
    .Y(_07473_));
 sky130_fd_sc_hd__nor2_8 _12561_ (.A(_07472_),
    .B(_07473_),
    .Y(_07474_));
 sky130_fd_sc_hd__inv_6 _12562_ (.A(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__nor2_1 _12563_ (.A(_06697_),
    .B(net817),
    .Y(_07476_));
 sky130_fd_sc_hd__or2_4 _12564_ (.A(_06697_),
    .B(net817),
    .X(_07477_));
 sky130_fd_sc_hd__nor2_8 _12565_ (.A(_04482_),
    .B(net1372),
    .Y(_07478_));
 sky130_fd_sc_hd__nand2_2 _12566_ (.A(net1241),
    .B(_07369_),
    .Y(_07479_));
 sky130_fd_sc_hd__mux2_1 _12567_ (.A0(_04477_),
    .A1(_07479_),
    .S(_06136_),
    .X(_07480_));
 sky130_fd_sc_hd__o22a_4 _12568_ (.A1(net1176),
    .A2(net813),
    .B1(_07480_),
    .B2(net830),
    .X(_07481_));
 sky130_fd_sc_hd__nor3_1 _12569_ (.A(_04468_),
    .B(_07446_),
    .C(_07481_),
    .Y(_07482_));
 sky130_fd_sc_hd__a21o_1 _12570_ (.A1(net1326),
    .A2(net1325),
    .B1(_04473_),
    .X(_07483_));
 sky130_fd_sc_hd__o311a_1 _12571_ (.A1(net1821),
    .A2(net1822),
    .A3(_04471_),
    .B1(_07483_),
    .C1(net1666),
    .X(_07484_));
 sky130_fd_sc_hd__nand2_1 _12572_ (.A(\core.pipe0_currentInstruction[5] ),
    .B(\core.pipe0_currentInstruction[4] ),
    .Y(_07485_));
 sky130_fd_sc_hd__a21o_2 _12573_ (.A1(\core.pipe0_currentInstruction[6] ),
    .A2(net1662),
    .B1(_07485_),
    .X(_07486_));
 sky130_fd_sc_hd__nor3_2 _12574_ (.A(_04462_),
    .B(_07484_),
    .C(_07486_),
    .Y(_07487_));
 sky130_fd_sc_hd__inv_2 _12575_ (.A(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__nor2_1 _12576_ (.A(_04478_),
    .B(_07487_),
    .Y(_07489_));
 sky130_fd_sc_hd__or2_2 _12577_ (.A(_04478_),
    .B(_07487_),
    .X(_07490_));
 sky130_fd_sc_hd__and3_1 _12578_ (.A(_04480_),
    .B(net1184),
    .C(net1083),
    .X(_07491_));
 sky130_fd_sc_hd__and4_4 _12579_ (.A(_04447_),
    .B(_04452_),
    .C(_04457_),
    .D(net1329),
    .X(_07492_));
 sky130_fd_sc_hd__nor2_4 _12580_ (.A(_04456_),
    .B(_07486_),
    .Y(_07493_));
 sky130_fd_sc_hd__or2_2 _12581_ (.A(net1289),
    .B(_07493_),
    .X(_07494_));
 sky130_fd_sc_hd__or4_1 _12582_ (.A(net1668),
    .B(_04467_),
    .C(net1260),
    .D(_07413_),
    .X(_07495_));
 sky130_fd_sc_hd__nor4b_2 _12583_ (.A(_07492_),
    .B(_07494_),
    .C(_07495_),
    .D_N(_07491_),
    .Y(_07496_));
 sky130_fd_sc_hd__or3_1 _12584_ (.A(net1763),
    .B(net1837),
    .C(net1849),
    .X(_07497_));
 sky130_fd_sc_hd__or4_4 _12585_ (.A(_04471_),
    .B(_07416_),
    .C(_07419_),
    .D(_07497_),
    .X(_07498_));
 sky130_fd_sc_hd__inv_2 _12586_ (.A(_07498_),
    .Y(_07499_));
 sky130_fd_sc_hd__nor2_1 _12587_ (.A(_07446_),
    .B(_07498_),
    .Y(_07500_));
 sky130_fd_sc_hd__or4_1 _12588_ (.A(_04471_),
    .B(_07424_),
    .C(_07426_),
    .D(_07497_),
    .X(_07501_));
 sky130_fd_sc_hd__or3_1 _12589_ (.A(_07482_),
    .B(net1019),
    .C(_07500_),
    .X(_07502_));
 sky130_fd_sc_hd__nor2_2 _12590_ (.A(_04482_),
    .B(_07481_),
    .Y(_07503_));
 sky130_fd_sc_hd__or2_4 _12591_ (.A(_04482_),
    .B(_07481_),
    .X(_07504_));
 sky130_fd_sc_hd__or4b_4 _12592_ (.A(_07499_),
    .B(_07502_),
    .C(net811),
    .D_N(_07470_),
    .X(\core.csr.inTrap ));
 sky130_fd_sc_hd__or2_4 _12593_ (.A(\coreWBInterface.state[1] ),
    .B(\coreWBInterface.state[0] ),
    .X(_07505_));
 sky130_fd_sc_hd__and2_1 _12594_ (.A(net1815),
    .B(net792),
    .X(_07506_));
 sky130_fd_sc_hd__nand2_2 _12595_ (.A(net1815),
    .B(net792),
    .Y(_07507_));
 sky130_fd_sc_hd__o21a_1 _12596_ (.A1(net461),
    .A2(_07403_),
    .B1(net472),
    .X(_07508_));
 sky130_fd_sc_hd__and2_2 _12597_ (.A(net475),
    .B(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__and3_1 _12598_ (.A(net477),
    .B(net476),
    .C(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__and2_2 _12599_ (.A(net478),
    .B(_07510_),
    .X(_07511_));
 sky130_fd_sc_hd__and3_1 _12600_ (.A(net480),
    .B(net479),
    .C(_07511_),
    .X(_07512_));
 sky130_fd_sc_hd__and2_2 _12601_ (.A(net481),
    .B(_07512_),
    .X(_07513_));
 sky130_fd_sc_hd__and3_1 _12602_ (.A(net452),
    .B(net451),
    .C(_07513_),
    .X(_07514_));
 sky130_fd_sc_hd__and2_2 _12603_ (.A(net453),
    .B(_07514_),
    .X(_07515_));
 sky130_fd_sc_hd__and3_1 _12604_ (.A(net455),
    .B(net454),
    .C(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__and2_2 _12605_ (.A(net456),
    .B(_07516_),
    .X(_07517_));
 sky130_fd_sc_hd__and3_1 _12606_ (.A(net458),
    .B(net457),
    .C(_07517_),
    .X(_07518_));
 sky130_fd_sc_hd__and2_4 _12607_ (.A(net459),
    .B(_07518_),
    .X(_07519_));
 sky130_fd_sc_hd__and3_1 _12608_ (.A(net462),
    .B(net460),
    .C(_07519_),
    .X(_07520_));
 sky130_fd_sc_hd__and2_2 _12609_ (.A(net463),
    .B(_07520_),
    .X(_07521_));
 sky130_fd_sc_hd__and3_1 _12610_ (.A(net465),
    .B(net464),
    .C(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__and2_2 _12611_ (.A(net466),
    .B(_07522_),
    .X(_07523_));
 sky130_fd_sc_hd__and3_1 _12612_ (.A(net468),
    .B(net467),
    .C(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__and2_1 _12613_ (.A(net469),
    .B(_07524_),
    .X(_07525_));
 sky130_fd_sc_hd__and3_1 _12614_ (.A(net471),
    .B(net470),
    .C(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__nand2_2 _12615_ (.A(net473),
    .B(_07526_),
    .Y(_07527_));
 sky130_fd_sc_hd__or2_1 _12616_ (.A(net473),
    .B(_07526_),
    .X(_07528_));
 sky130_fd_sc_hd__nand2_2 _12617_ (.A(_07527_),
    .B(_07528_),
    .Y(_07529_));
 sky130_fd_sc_hd__o2bb2a_1 _12618_ (.A1_N(_07396_),
    .A2_N(_07529_),
    .B1(_07346_),
    .B2(net1226),
    .X(_07530_));
 sky130_fd_sc_hd__a21oi_4 _12619_ (.A1(net799),
    .A2(net1259),
    .B1(net1295),
    .Y(_07531_));
 sky130_fd_sc_hd__a21o_4 _12620_ (.A1(net800),
    .A2(net1260),
    .B1(net1296),
    .X(_07532_));
 sky130_fd_sc_hd__o22a_1 _12621_ (.A1(net1291),
    .A2(_07530_),
    .B1(net790),
    .B2(net473),
    .X(_07533_));
 sky130_fd_sc_hd__nand2_1 _12622_ (.A(net786),
    .B(_07533_),
    .Y(_07534_));
 sky130_fd_sc_hd__a21oi_1 _12623_ (.A1(net470),
    .A2(_07525_),
    .B1(net471),
    .Y(_07535_));
 sky130_fd_sc_hd__or2_2 _12624_ (.A(_07526_),
    .B(_07535_),
    .X(_07536_));
 sky130_fd_sc_hd__o2bb2a_1 _12625_ (.A1_N(_07396_),
    .A2_N(_07536_),
    .B1(_07190_),
    .B2(net1227),
    .X(_07537_));
 sky130_fd_sc_hd__o22a_1 _12626_ (.A1(net471),
    .A2(net790),
    .B1(_07537_),
    .B2(net1291),
    .X(_07538_));
 sky130_fd_sc_hd__nand2_1 _12627_ (.A(_07506_),
    .B(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__or2_1 _12628_ (.A(_07506_),
    .B(_07538_),
    .X(_07540_));
 sky130_fd_sc_hd__nand2_1 _12629_ (.A(_07539_),
    .B(_07540_),
    .Y(_07541_));
 sky130_fd_sc_hd__xnor2_2 _12630_ (.A(net479),
    .B(_07511_),
    .Y(_07542_));
 sky130_fd_sc_hd__a211o_1 _12631_ (.A1(net801),
    .A2(net1261),
    .B1(net1231),
    .C1(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__nand2_1 _12632_ (.A(_05628_),
    .B(net1231),
    .Y(_07544_));
 sky130_fd_sc_hd__a21oi_2 _12633_ (.A1(_07543_),
    .A2(_07544_),
    .B1(net1296),
    .Y(_07545_));
 sky130_fd_sc_hd__nor2_2 _12634_ (.A(_04406_),
    .B(_07531_),
    .Y(_07546_));
 sky130_fd_sc_hd__o211a_1 _12635_ (.A1(_07545_),
    .A2(_07546_),
    .B1(net1820),
    .C1(net795),
    .X(_07547_));
 sky130_fd_sc_hd__o211ai_1 _12636_ (.A1(_07545_),
    .A2(_07546_),
    .B1(net1820),
    .C1(net795),
    .Y(_07548_));
 sky130_fd_sc_hd__a211oi_2 _12637_ (.A1(net1820),
    .A2(net795),
    .B1(_07545_),
    .C1(_07546_),
    .Y(_07549_));
 sky130_fd_sc_hd__nor2_1 _12638_ (.A(net478),
    .B(_07510_),
    .Y(_07550_));
 sky130_fd_sc_hd__or2_2 _12639_ (.A(_07511_),
    .B(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__a211o_1 _12640_ (.A1(net800),
    .A2(net1261),
    .B1(net1231),
    .C1(_07551_),
    .X(_07552_));
 sky130_fd_sc_hd__nand2_1 _12641_ (.A(_05709_),
    .B(net1231),
    .Y(_07553_));
 sky130_fd_sc_hd__a21oi_2 _12642_ (.A1(_07552_),
    .A2(_07553_),
    .B1(net1296),
    .Y(_07554_));
 sky130_fd_sc_hd__and2_1 _12643_ (.A(net478),
    .B(net789),
    .X(_07555_));
 sky130_fd_sc_hd__o211a_2 _12644_ (.A1(_07554_),
    .A2(_07555_),
    .B1(net1821),
    .C1(net795),
    .X(_07556_));
 sky130_fd_sc_hd__nand2b_1 _12645_ (.A_N(_07549_),
    .B(_07556_),
    .Y(_07557_));
 sky130_fd_sc_hd__a21oi_1 _12646_ (.A1(net476),
    .A2(_07509_),
    .B1(net477),
    .Y(_07558_));
 sky130_fd_sc_hd__or2_1 _12647_ (.A(_07510_),
    .B(_07558_),
    .X(_07559_));
 sky130_fd_sc_hd__a211o_1 _12648_ (.A1(net800),
    .A2(net1261),
    .B1(net1231),
    .C1(_07559_),
    .X(_07560_));
 sky130_fd_sc_hd__nand2_1 _12649_ (.A(_05794_),
    .B(net1231),
    .Y(_07561_));
 sky130_fd_sc_hd__a21oi_2 _12650_ (.A1(_07560_),
    .A2(_07561_),
    .B1(net1296),
    .Y(_07562_));
 sky130_fd_sc_hd__and2_1 _12651_ (.A(net477),
    .B(net789),
    .X(_07563_));
 sky130_fd_sc_hd__and2_1 _12652_ (.A(\core.pipe0_currentInstruction[25] ),
    .B(net796),
    .X(_07564_));
 sky130_fd_sc_hd__nor3_2 _12653_ (.A(_07562_),
    .B(_07563_),
    .C(_07564_),
    .Y(_07565_));
 sky130_fd_sc_hd__a22oi_4 _12654_ (.A1(\core.pipe0_currentInstruction[10] ),
    .A2(_07392_),
    .B1(net1183),
    .B2(net1831),
    .Y(_07566_));
 sky130_fd_sc_hd__nor2_1 _12655_ (.A(net475),
    .B(_07508_),
    .Y(_07567_));
 sky130_fd_sc_hd__or2_1 _12656_ (.A(_07509_),
    .B(_07567_),
    .X(_07568_));
 sky130_fd_sc_hd__a211o_1 _12657_ (.A1(net800),
    .A2(net1261),
    .B1(net1231),
    .C1(_07568_),
    .X(_07569_));
 sky130_fd_sc_hd__nand2_1 _12658_ (.A(_05962_),
    .B(net1232),
    .Y(_07570_));
 sky130_fd_sc_hd__a21o_1 _12659_ (.A1(_07569_),
    .A2(_07570_),
    .B1(net1296),
    .X(_07571_));
 sky130_fd_sc_hd__nand2_1 _12660_ (.A(net475),
    .B(net789),
    .Y(_07572_));
 sky130_fd_sc_hd__a21oi_2 _12661_ (.A1(_07571_),
    .A2(_07572_),
    .B1(_07566_),
    .Y(_07573_));
 sky130_fd_sc_hd__and3_2 _12662_ (.A(_07566_),
    .B(_07571_),
    .C(_07572_),
    .X(_07574_));
 sky130_fd_sc_hd__o2bb2a_1 _12663_ (.A1_N(\core.pipe0_currentInstruction[9] ),
    .A2_N(_07392_),
    .B1(net1184),
    .B2(net1746),
    .X(_07575_));
 sky130_fd_sc_hd__nor3_1 _12664_ (.A(net472),
    .B(net461),
    .C(_07403_),
    .Y(_07576_));
 sky130_fd_sc_hd__nor2_1 _12665_ (.A(_07508_),
    .B(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__inv_2 _12666_ (.A(_07577_),
    .Y(_07578_));
 sky130_fd_sc_hd__a211o_1 _12667_ (.A1(net800),
    .A2(net1260),
    .B1(net1231),
    .C1(_07578_),
    .X(_07579_));
 sky130_fd_sc_hd__or2_1 _12668_ (.A(_06046_),
    .B(net1228),
    .X(_07580_));
 sky130_fd_sc_hd__a21o_1 _12669_ (.A1(_07579_),
    .A2(_07580_),
    .B1(net1297),
    .X(_07581_));
 sky130_fd_sc_hd__nand2_1 _12670_ (.A(net472),
    .B(net789),
    .Y(_07582_));
 sky130_fd_sc_hd__a21oi_1 _12671_ (.A1(_07581_),
    .A2(_07582_),
    .B1(_07575_),
    .Y(_07583_));
 sky130_fd_sc_hd__a21o_1 _12672_ (.A1(_07581_),
    .A2(_07582_),
    .B1(_07575_),
    .X(_07584_));
 sky130_fd_sc_hd__o21ai_2 _12673_ (.A1(_07409_),
    .A2(_07410_),
    .B1(_07408_),
    .Y(_07585_));
 sky130_fd_sc_hd__nand3_1 _12674_ (.A(_07575_),
    .B(_07581_),
    .C(_07582_),
    .Y(_07586_));
 sky130_fd_sc_hd__and3_1 _12675_ (.A(_07584_),
    .B(_07585_),
    .C(_07586_),
    .X(_07587_));
 sky130_fd_sc_hd__nor2_1 _12676_ (.A(_07583_),
    .B(_07587_),
    .Y(_07588_));
 sky130_fd_sc_hd__a211o_1 _12677_ (.A1(_07585_),
    .A2(_07586_),
    .B1(_07573_),
    .C1(_07583_),
    .X(_07589_));
 sky130_fd_sc_hd__and2b_1 _12678_ (.A_N(_07574_),
    .B(_07589_),
    .X(_07590_));
 sky130_fd_sc_hd__o2bb2a_2 _12679_ (.A1_N(\core.pipe0_currentInstruction[11] ),
    .A2_N(_07392_),
    .B1(net1185),
    .B2(net1752),
    .X(_07591_));
 sky130_fd_sc_hd__xnor2_1 _12680_ (.A(net476),
    .B(_07509_),
    .Y(_07592_));
 sky130_fd_sc_hd__a211o_1 _12681_ (.A1(net801),
    .A2(net1260),
    .B1(net1231),
    .C1(_07592_),
    .X(_07593_));
 sky130_fd_sc_hd__nand2_1 _12682_ (.A(_05878_),
    .B(net1231),
    .Y(_07594_));
 sky130_fd_sc_hd__a21o_1 _12683_ (.A1(_07593_),
    .A2(_07594_),
    .B1(net1297),
    .X(_07595_));
 sky130_fd_sc_hd__nand2_2 _12684_ (.A(net476),
    .B(net789),
    .Y(_07596_));
 sky130_fd_sc_hd__a21oi_4 _12685_ (.A1(_07595_),
    .A2(_07596_),
    .B1(_07591_),
    .Y(_07597_));
 sky130_fd_sc_hd__and3_1 _12686_ (.A(_07591_),
    .B(_07595_),
    .C(_07596_),
    .X(_07598_));
 sky130_fd_sc_hd__nor2_1 _12687_ (.A(_07597_),
    .B(_07598_),
    .Y(_07599_));
 sky130_fd_sc_hd__and2_1 _12688_ (.A(_07590_),
    .B(_07599_),
    .X(_07600_));
 sky130_fd_sc_hd__o21a_1 _12689_ (.A1(_07562_),
    .A2(_07563_),
    .B1(_07564_),
    .X(_07601_));
 sky130_fd_sc_hd__nor2_1 _12690_ (.A(_07597_),
    .B(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__nor2_1 _12691_ (.A(_07565_),
    .B(_07601_),
    .Y(_07603_));
 sky130_fd_sc_hd__or4_1 _12692_ (.A(_07565_),
    .B(_07597_),
    .C(_07598_),
    .D(_07601_),
    .X(_07604_));
 sky130_fd_sc_hd__nor2_1 _12693_ (.A(_07565_),
    .B(_07602_),
    .Y(_07605_));
 sky130_fd_sc_hd__a21o_1 _12694_ (.A1(_07600_),
    .A2(_07603_),
    .B1(_07605_),
    .X(_07606_));
 sky130_fd_sc_hd__a211oi_2 _12695_ (.A1(net1821),
    .A2(net795),
    .B1(_07554_),
    .C1(_07555_),
    .Y(_07607_));
 sky130_fd_sc_hd__nor2_1 _12696_ (.A(_07547_),
    .B(_07549_),
    .Y(_07608_));
 sky130_fd_sc_hd__nor2_2 _12697_ (.A(_07556_),
    .B(_07607_),
    .Y(_07609_));
 sky130_fd_sc_hd__or4_1 _12698_ (.A(_07547_),
    .B(_07549_),
    .C(_07556_),
    .D(_07607_),
    .X(_07610_));
 sky130_fd_sc_hd__or4b_4 _12699_ (.A(_07574_),
    .B(_07604_),
    .C(_07610_),
    .D_N(_07589_),
    .X(_07611_));
 sky130_fd_sc_hd__o311a_2 _12700_ (.A1(_07565_),
    .A2(_07602_),
    .A3(_07610_),
    .B1(_07557_),
    .C1(_07548_),
    .X(_07612_));
 sky130_fd_sc_hd__nand2_1 _12701_ (.A(_07611_),
    .B(_07612_),
    .Y(_07613_));
 sky130_fd_sc_hd__nor2_1 _12702_ (.A(net456),
    .B(_07516_),
    .Y(_07614_));
 sky130_fd_sc_hd__or2_1 _12703_ (.A(_07517_),
    .B(_07614_),
    .X(_07615_));
 sky130_fd_sc_hd__a211o_1 _12704_ (.A1(net799),
    .A2(net1259),
    .B1(net1229),
    .C1(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__nand2_1 _12705_ (.A(_05186_),
    .B(net1230),
    .Y(_07617_));
 sky130_fd_sc_hd__a21oi_2 _12706_ (.A1(_07616_),
    .A2(_07617_),
    .B1(net1294),
    .Y(_07618_));
 sky130_fd_sc_hd__and2_1 _12707_ (.A(net456),
    .B(net789),
    .X(_07619_));
 sky130_fd_sc_hd__or2_4 _12708_ (.A(net1815),
    .B(net1297),
    .X(_07620_));
 sky130_fd_sc_hd__and2_4 _12709_ (.A(net794),
    .B(_07620_),
    .X(_07621_));
 sky130_fd_sc_hd__nand2_4 _12710_ (.A(net793),
    .B(_07620_),
    .Y(_07622_));
 sky130_fd_sc_hd__nand2_1 _12711_ (.A(net1688),
    .B(net1295),
    .Y(_07623_));
 sky130_fd_sc_hd__o211a_1 _12712_ (.A1(_07618_),
    .A2(_07619_),
    .B1(_07621_),
    .C1(_07623_),
    .X(_07624_));
 sky130_fd_sc_hd__a211oi_2 _12713_ (.A1(_07621_),
    .A2(_07623_),
    .B1(_07618_),
    .C1(_07619_),
    .Y(_07625_));
 sky130_fd_sc_hd__a211o_1 _12714_ (.A1(_07621_),
    .A2(_07623_),
    .B1(_07618_),
    .C1(_07619_),
    .X(_07626_));
 sky130_fd_sc_hd__nor2_1 _12715_ (.A(_07624_),
    .B(_07625_),
    .Y(_07627_));
 sky130_fd_sc_hd__nand2_1 _12716_ (.A(_04423_),
    .B(net1295),
    .Y(_07628_));
 sky130_fd_sc_hd__a21oi_1 _12717_ (.A1(net454),
    .A2(_07515_),
    .B1(net455),
    .Y(_07629_));
 sky130_fd_sc_hd__or2_1 _12718_ (.A(_07516_),
    .B(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__a211o_1 _12719_ (.A1(net801),
    .A2(net1262),
    .B1(net1230),
    .C1(_07630_),
    .X(_07631_));
 sky130_fd_sc_hd__nand2_1 _12720_ (.A(_05275_),
    .B(net1230),
    .Y(_07632_));
 sky130_fd_sc_hd__a21oi_2 _12721_ (.A1(_07631_),
    .A2(_07632_),
    .B1(net1295),
    .Y(_07633_));
 sky130_fd_sc_hd__and2_1 _12722_ (.A(net455),
    .B(net789),
    .X(_07634_));
 sky130_fd_sc_hd__o211a_2 _12723_ (.A1(_07633_),
    .A2(_07634_),
    .B1(_07621_),
    .C1(_07628_),
    .X(_07635_));
 sky130_fd_sc_hd__a211oi_2 _12724_ (.A1(_07621_),
    .A2(_07628_),
    .B1(_07633_),
    .C1(_07634_),
    .Y(_07636_));
 sky130_fd_sc_hd__or2_1 _12725_ (.A(_07635_),
    .B(_07636_),
    .X(_07637_));
 sky130_fd_sc_hd__or4_4 _12726_ (.A(_07624_),
    .B(_07625_),
    .C(_07635_),
    .D(_07636_),
    .X(_07638_));
 sky130_fd_sc_hd__o211ai_4 _12727_ (.A1(net1881),
    .A2(net1290),
    .B1(net794),
    .C1(_07620_),
    .Y(_07639_));
 sky130_fd_sc_hd__nor2_1 _12728_ (.A(net453),
    .B(_07514_),
    .Y(_07640_));
 sky130_fd_sc_hd__or2_1 _12729_ (.A(_07515_),
    .B(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__a211o_1 _12730_ (.A1(net801),
    .A2(net1262),
    .B1(net1230),
    .C1(_07641_),
    .X(_07642_));
 sky130_fd_sc_hd__nand2_1 _12731_ (.A(_05022_),
    .B(net1230),
    .Y(_07643_));
 sky130_fd_sc_hd__a21o_1 _12732_ (.A1(_07642_),
    .A2(_07643_),
    .B1(net1295),
    .X(_07644_));
 sky130_fd_sc_hd__nand2_1 _12733_ (.A(net453),
    .B(net789),
    .Y(_07645_));
 sky130_fd_sc_hd__a21oi_1 _12734_ (.A1(_07644_),
    .A2(_07645_),
    .B1(_07639_),
    .Y(_07646_));
 sky130_fd_sc_hd__a21o_2 _12735_ (.A1(_07644_),
    .A2(_07645_),
    .B1(_07639_),
    .X(_07647_));
 sky130_fd_sc_hd__and3_1 _12736_ (.A(_07639_),
    .B(_07644_),
    .C(_07645_),
    .X(_07648_));
 sky130_fd_sc_hd__nor2_1 _12737_ (.A(_07646_),
    .B(_07648_),
    .Y(_07649_));
 sky130_fd_sc_hd__nor2_1 _12738_ (.A(_05107_),
    .B(net1228),
    .Y(_07650_));
 sky130_fd_sc_hd__inv_2 _12739_ (.A(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__xnor2_1 _12740_ (.A(net454),
    .B(_07515_),
    .Y(_07652_));
 sky130_fd_sc_hd__inv_2 _12741_ (.A(_07652_),
    .Y(_07653_));
 sky130_fd_sc_hd__a211o_1 _12742_ (.A1(net799),
    .A2(net1259),
    .B1(net1229),
    .C1(_07653_),
    .X(_07654_));
 sky130_fd_sc_hd__a21o_2 _12743_ (.A1(_07651_),
    .A2(_07654_),
    .B1(net1295),
    .X(_07655_));
 sky130_fd_sc_hd__or2_4 _12744_ (.A(net454),
    .B(_07531_),
    .X(_07656_));
 sky130_fd_sc_hd__o211a_2 _12745_ (.A1(net1880),
    .A2(_04454_),
    .B1(net794),
    .C1(_07620_),
    .X(_07657_));
 sky130_fd_sc_hd__a21oi_4 _12746_ (.A1(_07655_),
    .A2(_07656_),
    .B1(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__nand3_4 _12747_ (.A(_07655_),
    .B(_07656_),
    .C(_07657_),
    .Y(_07659_));
 sky130_fd_sc_hd__and2b_1 _12748_ (.A_N(_07658_),
    .B(_07659_),
    .X(_07660_));
 sky130_fd_sc_hd__or4b_1 _12749_ (.A(_07646_),
    .B(_07648_),
    .C(_07658_),
    .D_N(_07659_),
    .X(_07661_));
 sky130_fd_sc_hd__nor2_1 _12750_ (.A(_07638_),
    .B(_07661_),
    .Y(_07662_));
 sky130_fd_sc_hd__a22o_2 _12751_ (.A1(\core.pipe0_currentInstruction[7] ),
    .A2(_07392_),
    .B1(net1183),
    .B2(_07620_),
    .X(_07663_));
 sky130_fd_sc_hd__nand2_1 _12752_ (.A(net1725),
    .B(net1296),
    .Y(_07664_));
 sky130_fd_sc_hd__a21oi_1 _12753_ (.A1(net451),
    .A2(_07513_),
    .B1(net452),
    .Y(_07665_));
 sky130_fd_sc_hd__or2_1 _12754_ (.A(_07514_),
    .B(_07665_),
    .X(_07666_));
 sky130_fd_sc_hd__a211o_1 _12755_ (.A1(net800),
    .A2(net1260),
    .B1(net1232),
    .C1(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__nand2_1 _12756_ (.A(_05330_),
    .B(net1232),
    .Y(_07668_));
 sky130_fd_sc_hd__a21oi_1 _12757_ (.A1(_07667_),
    .A2(_07668_),
    .B1(net1296),
    .Y(_07669_));
 sky130_fd_sc_hd__and2_1 _12758_ (.A(net452),
    .B(net789),
    .X(_07670_));
 sky130_fd_sc_hd__o211a_1 _12759_ (.A1(_07669_),
    .A2(_07670_),
    .B1(_07663_),
    .C1(_07664_),
    .X(_07671_));
 sky130_fd_sc_hd__a211o_1 _12760_ (.A1(_07663_),
    .A2(_07664_),
    .B1(_07669_),
    .C1(_07670_),
    .X(_07672_));
 sky130_fd_sc_hd__and2b_1 _12761_ (.A_N(_07671_),
    .B(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__xnor2_1 _12762_ (.A(net451),
    .B(_07513_),
    .Y(_07674_));
 sky130_fd_sc_hd__a211o_1 _12763_ (.A1(net800),
    .A2(net1260),
    .B1(net1232),
    .C1(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__nand2_2 _12764_ (.A(_05451_),
    .B(net1232),
    .Y(_07676_));
 sky130_fd_sc_hd__a21oi_4 _12765_ (.A1(_07675_),
    .A2(_07676_),
    .B1(net1296),
    .Y(_07677_));
 sky130_fd_sc_hd__and2_2 _12766_ (.A(net451),
    .B(_07532_),
    .X(_07678_));
 sky130_fd_sc_hd__or2_1 _12767_ (.A(_07677_),
    .B(_07678_),
    .X(_07679_));
 sky130_fd_sc_hd__o211ai_4 _12768_ (.A1(_07677_),
    .A2(_07678_),
    .B1(net1817),
    .C1(net794),
    .Y(_07680_));
 sky130_fd_sc_hd__a211o_1 _12769_ (.A1(net1817),
    .A2(net794),
    .B1(_07677_),
    .C1(_07678_),
    .X(_07681_));
 sky130_fd_sc_hd__nand2_1 _12770_ (.A(_07680_),
    .B(_07681_),
    .Y(_07682_));
 sky130_fd_sc_hd__nand4b_2 _12771_ (.A_N(_07671_),
    .B(_07672_),
    .C(_07680_),
    .D(_07681_),
    .Y(_07683_));
 sky130_fd_sc_hd__a21oi_1 _12772_ (.A1(net479),
    .A2(_07511_),
    .B1(net480),
    .Y(_07684_));
 sky130_fd_sc_hd__or2_1 _12773_ (.A(_07512_),
    .B(_07684_),
    .X(_07685_));
 sky130_fd_sc_hd__a211o_1 _12774_ (.A1(net800),
    .A2(net1260),
    .B1(net1232),
    .C1(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__nand2_1 _12775_ (.A(_06310_),
    .B(net1232),
    .Y(_07687_));
 sky130_fd_sc_hd__a21oi_2 _12776_ (.A1(_07686_),
    .A2(_07687_),
    .B1(net1296),
    .Y(_07688_));
 sky130_fd_sc_hd__and2_1 _12777_ (.A(net480),
    .B(_07532_),
    .X(_07689_));
 sky130_fd_sc_hd__o211a_2 _12778_ (.A1(_07688_),
    .A2(_07689_),
    .B1(net1819),
    .C1(net795),
    .X(_07690_));
 sky130_fd_sc_hd__a211oi_2 _12779_ (.A1(net1819),
    .A2(net795),
    .B1(_07688_),
    .C1(_07689_),
    .Y(_07691_));
 sky130_fd_sc_hd__nor2_1 _12780_ (.A(_07690_),
    .B(_07691_),
    .Y(_07692_));
 sky130_fd_sc_hd__nor2_1 _12781_ (.A(net481),
    .B(_07512_),
    .Y(_07693_));
 sky130_fd_sc_hd__or2_1 _12782_ (.A(_07513_),
    .B(_07693_),
    .X(_07694_));
 sky130_fd_sc_hd__a211o_1 _12783_ (.A1(net800),
    .A2(net1260),
    .B1(net1232),
    .C1(_07694_),
    .X(_07695_));
 sky130_fd_sc_hd__nand2_1 _12784_ (.A(_05547_),
    .B(net1232),
    .Y(_07696_));
 sky130_fd_sc_hd__a21oi_2 _12785_ (.A1(_07695_),
    .A2(_07696_),
    .B1(net1295),
    .Y(_07697_));
 sky130_fd_sc_hd__and2_1 _12786_ (.A(net481),
    .B(_07532_),
    .X(_07698_));
 sky130_fd_sc_hd__a211oi_2 _12787_ (.A1(\core.pipe0_currentInstruction[29] ),
    .A2(net796),
    .B1(_07697_),
    .C1(_07698_),
    .Y(_07699_));
 sky130_fd_sc_hd__o211a_1 _12788_ (.A1(_07697_),
    .A2(_07698_),
    .B1(\core.pipe0_currentInstruction[29] ),
    .C1(net796),
    .X(_07700_));
 sky130_fd_sc_hd__nor2_1 _12789_ (.A(_07699_),
    .B(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__or4_2 _12790_ (.A(_07690_),
    .B(_07691_),
    .C(_07699_),
    .D(_07700_),
    .X(_07702_));
 sky130_fd_sc_hd__or4_4 _12791_ (.A(_07638_),
    .B(_07661_),
    .C(_07683_),
    .D(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__a21o_4 _12792_ (.A1(_07611_),
    .A2(_07612_),
    .B1(_07703_),
    .X(_07704_));
 sky130_fd_sc_hd__a211oi_4 _12793_ (.A1(_07647_),
    .A2(_07659_),
    .B1(_07658_),
    .C1(_07638_),
    .Y(_07705_));
 sky130_fd_sc_hd__a21o_1 _12794_ (.A1(_07626_),
    .A2(_07635_),
    .B1(_07624_),
    .X(_07706_));
 sky130_fd_sc_hd__o21ba_1 _12795_ (.A1(_07690_),
    .A2(_07700_),
    .B1_N(_07699_),
    .X(_07707_));
 sky130_fd_sc_hd__a41o_1 _12796_ (.A1(net1817),
    .A2(net2013),
    .A3(_07672_),
    .A4(_07679_),
    .B1(_07671_),
    .X(_07708_));
 sky130_fd_sc_hd__a41o_2 _12797_ (.A1(_07673_),
    .A2(_07680_),
    .A3(_07681_),
    .A4(_07707_),
    .B1(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__a211oi_4 _12798_ (.A1(_07662_),
    .A2(_07709_),
    .B1(_07706_),
    .C1(_07705_),
    .Y(_07710_));
 sky130_fd_sc_hd__nor2_1 _12799_ (.A(net463),
    .B(_07520_),
    .Y(_07711_));
 sky130_fd_sc_hd__or2_1 _12800_ (.A(_07521_),
    .B(_07711_),
    .X(_07712_));
 sky130_fd_sc_hd__o2bb2a_1 _12801_ (.A1_N(_07396_),
    .A2_N(_07712_),
    .B1(_04849_),
    .B2(net1226),
    .X(_07713_));
 sky130_fd_sc_hd__o22a_4 _12802_ (.A1(net463),
    .A2(net790),
    .B1(_07713_),
    .B2(net1291),
    .X(_07714_));
 sky130_fd_sc_hd__xnor2_4 _12803_ (.A(net785),
    .B(_07714_),
    .Y(_07715_));
 sky130_fd_sc_hd__xnor2_1 _12804_ (.A(net464),
    .B(_07521_),
    .Y(_07716_));
 sky130_fd_sc_hd__o2bb2a_1 _12805_ (.A1_N(_07396_),
    .A2_N(_07716_),
    .B1(_04770_),
    .B2(net1226),
    .X(_07717_));
 sky130_fd_sc_hd__o22a_1 _12806_ (.A1(net464),
    .A2(net790),
    .B1(_07717_),
    .B2(net1291),
    .X(_07718_));
 sky130_fd_sc_hd__nand2_1 _12807_ (.A(net785),
    .B(_07718_),
    .Y(_07719_));
 sky130_fd_sc_hd__or2_1 _12808_ (.A(net785),
    .B(_07718_),
    .X(_07720_));
 sky130_fd_sc_hd__and2_2 _12809_ (.A(_07719_),
    .B(_07720_),
    .X(_07721_));
 sky130_fd_sc_hd__a21oi_1 _12810_ (.A1(net460),
    .A2(_07519_),
    .B1(net462),
    .Y(_07722_));
 sky130_fd_sc_hd__or2_1 _12811_ (.A(_07520_),
    .B(_07722_),
    .X(_07723_));
 sky130_fd_sc_hd__o2bb2a_1 _12812_ (.A1_N(_07396_),
    .A2_N(_07723_),
    .B1(_04926_),
    .B2(net1226),
    .X(_07724_));
 sky130_fd_sc_hd__o22a_4 _12813_ (.A1(net462),
    .A2(net790),
    .B1(_07724_),
    .B2(net1291),
    .X(_07725_));
 sky130_fd_sc_hd__nand2_1 _12814_ (.A(net785),
    .B(_07725_),
    .Y(_07726_));
 sky130_fd_sc_hd__xnor2_4 _12815_ (.A(net785),
    .B(_07725_),
    .Y(_07727_));
 sky130_fd_sc_hd__a21oi_1 _12816_ (.A1(net464),
    .A2(_07521_),
    .B1(net465),
    .Y(_07728_));
 sky130_fd_sc_hd__or2_1 _12817_ (.A(_07522_),
    .B(_07728_),
    .X(_07729_));
 sky130_fd_sc_hd__o2bb2a_1 _12818_ (.A1_N(_07396_),
    .A2_N(_07729_),
    .B1(_04692_),
    .B2(net1226),
    .X(_07730_));
 sky130_fd_sc_hd__o22a_2 _12819_ (.A1(net465),
    .A2(net790),
    .B1(_07730_),
    .B2(net1291),
    .X(_07731_));
 sky130_fd_sc_hd__xnor2_2 _12820_ (.A(net785),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__nor3_1 _12821_ (.A(_07715_),
    .B(_07727_),
    .C(_07732_),
    .Y(_07733_));
 sky130_fd_sc_hd__nand2_2 _12822_ (.A(_07721_),
    .B(_07733_),
    .Y(_07734_));
 sky130_fd_sc_hd__nand2_1 _12823_ (.A(_06560_),
    .B(net1229),
    .Y(_07735_));
 sky130_fd_sc_hd__xor2_2 _12824_ (.A(net460),
    .B(_07519_),
    .X(_07736_));
 sky130_fd_sc_hd__a211o_1 _12825_ (.A1(net2015),
    .A2(net1259),
    .B1(net1229),
    .C1(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__a21oi_4 _12826_ (.A1(_07735_),
    .A2(_07737_),
    .B1(net1294),
    .Y(_07738_));
 sky130_fd_sc_hd__nor2_2 _12827_ (.A(net460),
    .B(net791),
    .Y(_07739_));
 sky130_fd_sc_hd__nor2_2 _12828_ (.A(net1855),
    .B(net1290),
    .Y(_07740_));
 sky130_fd_sc_hd__nor4_2 _12829_ (.A(_07622_),
    .B(_07738_),
    .C(_07739_),
    .D(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__o22ai_4 _12830_ (.A1(_07738_),
    .A2(_07739_),
    .B1(_07740_),
    .B2(_07622_),
    .Y(_07742_));
 sky130_fd_sc_hd__nand2b_1 _12831_ (.A_N(_07741_),
    .B(_07742_),
    .Y(_07743_));
 sky130_fd_sc_hd__nor2_2 _12832_ (.A(\core.pipe0_currentInstruction[18] ),
    .B(net1290),
    .Y(_07744_));
 sky130_fd_sc_hd__nand2_2 _12833_ (.A(_06637_),
    .B(net1229),
    .Y(_07745_));
 sky130_fd_sc_hd__nor2_1 _12834_ (.A(net459),
    .B(_07518_),
    .Y(_07746_));
 sky130_fd_sc_hd__nor2_1 _12835_ (.A(_07519_),
    .B(_07746_),
    .Y(_07747_));
 sky130_fd_sc_hd__a211o_1 _12836_ (.A1(net2015),
    .A2(net1259),
    .B1(net1229),
    .C1(_07747_),
    .X(_07748_));
 sky130_fd_sc_hd__a21oi_4 _12837_ (.A1(_07745_),
    .A2(_07748_),
    .B1(net1294),
    .Y(_07749_));
 sky130_fd_sc_hd__nor2_2 _12838_ (.A(net459),
    .B(net791),
    .Y(_07750_));
 sky130_fd_sc_hd__or4_4 _12839_ (.A(_07622_),
    .B(_07744_),
    .C(_07749_),
    .D(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__o22ai_4 _12840_ (.A1(_07622_),
    .A2(_07744_),
    .B1(_07749_),
    .B2(_07750_),
    .Y(_07752_));
 sky130_fd_sc_hd__nand2_1 _12841_ (.A(_07751_),
    .B(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__nand4b_2 _12842_ (.A_N(_07741_),
    .B(_07742_),
    .C(_07751_),
    .D(_07752_),
    .Y(_07754_));
 sky130_fd_sc_hd__or2_1 _12843_ (.A(_06405_),
    .B(net1227),
    .X(_07755_));
 sky130_fd_sc_hd__a21oi_1 _12844_ (.A1(net457),
    .A2(_07517_),
    .B1(net458),
    .Y(_07756_));
 sky130_fd_sc_hd__or2_1 _12845_ (.A(_07518_),
    .B(_07756_),
    .X(_07757_));
 sky130_fd_sc_hd__inv_2 _12846_ (.A(_07757_),
    .Y(_07758_));
 sky130_fd_sc_hd__a211o_1 _12847_ (.A1(net2015),
    .A2(net1259),
    .B1(net1229),
    .C1(_07758_),
    .X(_07759_));
 sky130_fd_sc_hd__a21o_1 _12848_ (.A1(_07755_),
    .A2(_07759_),
    .B1(net1294),
    .X(_07760_));
 sky130_fd_sc_hd__or2_1 _12849_ (.A(net458),
    .B(net791),
    .X(_07761_));
 sky130_fd_sc_hd__o211a_1 _12850_ (.A1(net1863),
    .A2(net1290),
    .B1(net793),
    .C1(_07620_),
    .X(_07762_));
 sky130_fd_sc_hd__a21oi_1 _12851_ (.A1(_07760_),
    .A2(_07761_),
    .B1(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__nand3_1 _12852_ (.A(_07760_),
    .B(_07761_),
    .C(_07762_),
    .Y(_07764_));
 sky130_fd_sc_hd__nand2b_2 _12853_ (.A_N(_07763_),
    .B(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__o211a_2 _12854_ (.A1(net1871),
    .A2(net1290),
    .B1(net793),
    .C1(_07620_),
    .X(_07766_));
 sky130_fd_sc_hd__xor2_2 _12855_ (.A(net457),
    .B(_07517_),
    .X(_07767_));
 sky130_fd_sc_hd__o22a_2 _12856_ (.A1(_06483_),
    .A2(net1227),
    .B1(_07397_),
    .B2(_07767_),
    .X(_07768_));
 sky130_fd_sc_hd__or2_2 _12857_ (.A(net457),
    .B(net791),
    .X(_07769_));
 sky130_fd_sc_hd__o21a_1 _12858_ (.A1(net1294),
    .A2(_07768_),
    .B1(_07769_),
    .X(_07770_));
 sky130_fd_sc_hd__o211ai_4 _12859_ (.A1(net1294),
    .A2(_07768_),
    .B1(_07769_),
    .C1(_07766_),
    .Y(_07771_));
 sky130_fd_sc_hd__xnor2_2 _12860_ (.A(_07766_),
    .B(_07770_),
    .Y(_07772_));
 sky130_fd_sc_hd__or3_1 _12861_ (.A(_07754_),
    .B(_07765_),
    .C(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__a211o_4 _12862_ (.A1(_07704_),
    .A2(_07710_),
    .B1(_07734_),
    .C1(_07773_),
    .X(_07774_));
 sky130_fd_sc_hd__o21a_1 _12863_ (.A1(_07763_),
    .A2(_07771_),
    .B1(_07764_),
    .X(_07775_));
 sky130_fd_sc_hd__nand2b_1 _12864_ (.A_N(_07751_),
    .B(_07742_),
    .Y(_07776_));
 sky130_fd_sc_hd__o21ai_1 _12865_ (.A1(_07754_),
    .A2(_07775_),
    .B1(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__nor2_2 _12866_ (.A(_07741_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__o21a_2 _12867_ (.A1(_07714_),
    .A2(_07725_),
    .B1(net785),
    .X(_07779_));
 sky130_fd_sc_hd__o21a_1 _12868_ (.A1(_07718_),
    .A2(_07731_),
    .B1(net785),
    .X(_07780_));
 sky130_fd_sc_hd__nor2_1 _12869_ (.A(_07779_),
    .B(_07780_),
    .Y(_07781_));
 sky130_fd_sc_hd__o21a_1 _12870_ (.A1(_07734_),
    .A2(_07778_),
    .B1(_07781_),
    .X(_07782_));
 sky130_fd_sc_hd__nand2_1 _12871_ (.A(_07774_),
    .B(_07782_),
    .Y(_07783_));
 sky130_fd_sc_hd__nor2_1 _12872_ (.A(net466),
    .B(_07522_),
    .Y(_07784_));
 sky130_fd_sc_hd__or2_1 _12873_ (.A(_07523_),
    .B(_07784_),
    .X(_07785_));
 sky130_fd_sc_hd__o2bb2a_1 _12874_ (.A1_N(_07396_),
    .A2_N(_07785_),
    .B1(_06787_),
    .B2(net1226),
    .X(_07786_));
 sky130_fd_sc_hd__o22a_1 _12875_ (.A1(net466),
    .A2(net790),
    .B1(_07786_),
    .B2(net1291),
    .X(_07787_));
 sky130_fd_sc_hd__and2_1 _12876_ (.A(net786),
    .B(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__nor2_1 _12877_ (.A(net786),
    .B(_07787_),
    .Y(_07789_));
 sky130_fd_sc_hd__nor2_1 _12878_ (.A(_07788_),
    .B(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__nor2_1 _12879_ (.A(net469),
    .B(_07524_),
    .Y(_07791_));
 sky130_fd_sc_hd__or2_2 _12880_ (.A(_07525_),
    .B(_07791_),
    .X(_07792_));
 sky130_fd_sc_hd__o22a_1 _12881_ (.A1(_06943_),
    .A2(net1227),
    .B1(_07397_),
    .B2(_07792_),
    .X(_07793_));
 sky130_fd_sc_hd__a2bb2o_2 _12882_ (.A1_N(net1293),
    .A2_N(_07793_),
    .B1(net789),
    .B2(net469),
    .X(_07794_));
 sky130_fd_sc_hd__xnor2_2 _12883_ (.A(net786),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__xnor2_1 _12884_ (.A(net467),
    .B(_07523_),
    .Y(_07796_));
 sky130_fd_sc_hd__o2bb2a_1 _12885_ (.A1_N(_07396_),
    .A2_N(_07796_),
    .B1(_06865_),
    .B2(net1226),
    .X(_07797_));
 sky130_fd_sc_hd__o22a_2 _12886_ (.A1(net467),
    .A2(net790),
    .B1(_07797_),
    .B2(net1291),
    .X(_07798_));
 sky130_fd_sc_hd__xnor2_2 _12887_ (.A(_07507_),
    .B(_07798_),
    .Y(_07799_));
 sky130_fd_sc_hd__a21oi_1 _12888_ (.A1(net467),
    .A2(_07523_),
    .B1(net468),
    .Y(_07800_));
 sky130_fd_sc_hd__or2_1 _12889_ (.A(_07524_),
    .B(_07800_),
    .X(_07801_));
 sky130_fd_sc_hd__o2bb2a_1 _12890_ (.A1_N(_07396_),
    .A2_N(_07801_),
    .B1(_07020_),
    .B2(net1227),
    .X(_07802_));
 sky130_fd_sc_hd__o22a_1 _12891_ (.A1(net468),
    .A2(net791),
    .B1(_07802_),
    .B2(net1292),
    .X(_07803_));
 sky130_fd_sc_hd__nand2_1 _12892_ (.A(net786),
    .B(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__or2_1 _12893_ (.A(net786),
    .B(_07803_),
    .X(_07805_));
 sky130_fd_sc_hd__and2_1 _12894_ (.A(_07804_),
    .B(_07805_),
    .X(_07806_));
 sky130_fd_sc_hd__nand2_1 _12895_ (.A(_07790_),
    .B(_07799_),
    .Y(_07807_));
 sky130_fd_sc_hd__or3b_1 _12896_ (.A(_07807_),
    .B(_07795_),
    .C_N(_07806_),
    .X(_07808_));
 sky130_fd_sc_hd__a21o_1 _12897_ (.A1(_07774_),
    .A2(_07782_),
    .B1(_07808_),
    .X(_07809_));
 sky130_fd_sc_hd__o21a_1 _12898_ (.A1(_07787_),
    .A2(_07798_),
    .B1(net786),
    .X(_07810_));
 sky130_fd_sc_hd__o21a_1 _12899_ (.A1(_07794_),
    .A2(_07803_),
    .B1(net786),
    .X(_07811_));
 sky130_fd_sc_hd__nor2_1 _12900_ (.A(_07810_),
    .B(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__xnor2_1 _12901_ (.A(net470),
    .B(_07525_),
    .Y(_07813_));
 sky130_fd_sc_hd__inv_2 _12902_ (.A(_07813_),
    .Y(_07814_));
 sky130_fd_sc_hd__o22a_1 _12903_ (.A1(_07107_),
    .A2(net1226),
    .B1(_07397_),
    .B2(_07814_),
    .X(_07815_));
 sky130_fd_sc_hd__o22a_1 _12904_ (.A1(net470),
    .A2(net790),
    .B1(_07815_),
    .B2(net1291),
    .X(_07816_));
 sky130_fd_sc_hd__nand2_2 _12905_ (.A(net785),
    .B(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__or2_1 _12906_ (.A(net785),
    .B(_07816_),
    .X(_07818_));
 sky130_fd_sc_hd__and2_1 _12907_ (.A(_07817_),
    .B(_07818_),
    .X(_07819_));
 sky130_fd_sc_hd__inv_2 _12908_ (.A(_07819_),
    .Y(_07820_));
 sky130_fd_sc_hd__a21o_1 _12909_ (.A1(_07809_),
    .A2(_07812_),
    .B1(_07820_),
    .X(_07821_));
 sky130_fd_sc_hd__a211o_1 _12910_ (.A1(_07809_),
    .A2(_07812_),
    .B1(_07820_),
    .C1(_07541_),
    .X(_07822_));
 sky130_fd_sc_hd__or2_1 _12911_ (.A(net786),
    .B(_07533_),
    .X(_07823_));
 sky130_fd_sc_hd__nand2_1 _12912_ (.A(_07534_),
    .B(_07823_),
    .Y(_07824_));
 sky130_fd_sc_hd__a31o_1 _12913_ (.A1(_07539_),
    .A2(_07817_),
    .A3(_07822_),
    .B1(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__xnor2_2 _12914_ (.A(_04403_),
    .B(_07527_),
    .Y(_07826_));
 sky130_fd_sc_hd__o22a_1 _12915_ (.A1(_07273_),
    .A2(net1226),
    .B1(_07397_),
    .B2(_07826_),
    .X(_07827_));
 sky130_fd_sc_hd__o22a_1 _12916_ (.A1(_04403_),
    .A2(net790),
    .B1(_07827_),
    .B2(net1291),
    .X(_07828_));
 sky130_fd_sc_hd__xnor2_1 _12917_ (.A(_07507_),
    .B(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__a21oi_1 _12918_ (.A1(_07534_),
    .A2(_07825_),
    .B1(_07829_),
    .Y(_07830_));
 sky130_fd_sc_hd__a31o_1 _12919_ (.A1(_07534_),
    .A2(_07825_),
    .A3(_07829_),
    .B1(_07402_),
    .X(_07831_));
 sky130_fd_sc_hd__o21a_1 _12920_ (.A1(_07830_),
    .A2(_07831_),
    .B1(net792),
    .X(_07832_));
 sky130_fd_sc_hd__and3b_4 _12921_ (.A_N(\jtag.managementState[1] ),
    .B(_04397_),
    .C(\jtag.managementState[2] ),
    .X(_07833_));
 sky130_fd_sc_hd__or2_4 _12922_ (.A(\jtag.managementState[2] ),
    .B(\jtag.managementState[1] ),
    .X(_07834_));
 sky130_fd_sc_hd__or2_4 _12923_ (.A(_04397_),
    .B(net1639),
    .X(_07835_));
 sky130_fd_sc_hd__nand2b_4 _12924_ (.A_N(net1369),
    .B(_07835_),
    .Y(_07836_));
 sky130_fd_sc_hd__or2_4 _12925_ (.A(\wbSRAMInterface.state[1] ),
    .B(\wbSRAMInterface.state[0] ),
    .X(_07837_));
 sky130_fd_sc_hd__nand2_2 _12926_ (.A(\wbSRAMInterface.state[1] ),
    .B(\wbSRAMInterface.state[0] ),
    .Y(_07838_));
 sky130_fd_sc_hd__nand2_4 _12927_ (.A(_07837_),
    .B(_07838_),
    .Y(_07839_));
 sky130_fd_sc_hd__or4b_4 _12928_ (.A(net203),
    .B(net202),
    .C(net204),
    .D_N(net205),
    .X(_07840_));
 sky130_fd_sc_hd__nor2_8 _12929_ (.A(_07839_),
    .B(_07840_),
    .Y(_07841_));
 sky130_fd_sc_hd__and2b_2 _12930_ (.A_N(net1307),
    .B(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__a22o_4 _12931_ (.A1(\jtag.managementAddress[3] ),
    .A2(net1306),
    .B1(net1256),
    .B2(\wbSRAMInterface.currentAddress[3] ),
    .X(_07843_));
 sky130_fd_sc_hd__a22o_2 _12932_ (.A1(\jtag.managementAddress[6] ),
    .A2(net1306),
    .B1(net1255),
    .B2(\wbSRAMInterface.currentAddress[6] ),
    .X(_07844_));
 sky130_fd_sc_hd__a22oi_4 _12933_ (.A1(\jtag.managementAddress[14] ),
    .A2(net1307),
    .B1(net1256),
    .B2(\wbSRAMInterface.currentAddress[14] ),
    .Y(_07845_));
 sky130_fd_sc_hd__inv_2 _12934_ (.A(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__a22o_2 _12935_ (.A1(\jtag.managementAddress[15] ),
    .A2(net1307),
    .B1(net1256),
    .B2(\wbSRAMInterface.currentAddress[15] ),
    .X(_07847_));
 sky130_fd_sc_hd__a22o_4 _12936_ (.A1(\jtag.managementAddress[13] ),
    .A2(net1307),
    .B1(_07842_),
    .B2(\wbSRAMInterface.currentAddress[13] ),
    .X(_07848_));
 sky130_fd_sc_hd__a22o_2 _12937_ (.A1(\jtag.managementAddress[8] ),
    .A2(net1306),
    .B1(net1255),
    .B2(\wbSRAMInterface.currentAddress[8] ),
    .X(_07849_));
 sky130_fd_sc_hd__a22o_1 _12938_ (.A1(\jtag.managementAddress[11] ),
    .A2(net1306),
    .B1(net1255),
    .B2(\wbSRAMInterface.currentAddress[11] ),
    .X(_07850_));
 sky130_fd_sc_hd__a22o_2 _12939_ (.A1(\jtag.managementAddress[10] ),
    .A2(net1306),
    .B1(net1255),
    .B2(\wbSRAMInterface.currentAddress[10] ),
    .X(_07851_));
 sky130_fd_sc_hd__a22o_1 _12940_ (.A1(\jtag.managementAddress[9] ),
    .A2(net1306),
    .B1(net1255),
    .B2(\wbSRAMInterface.currentAddress[9] ),
    .X(_07852_));
 sky130_fd_sc_hd__a22o_1 _12941_ (.A1(\jtag.managementAddress[7] ),
    .A2(net1306),
    .B1(net1255),
    .B2(\wbSRAMInterface.currentAddress[7] ),
    .X(_07853_));
 sky130_fd_sc_hd__a22o_2 _12942_ (.A1(\jtag.managementAddress[12] ),
    .A2(net1307),
    .B1(_07842_),
    .B2(\wbSRAMInterface.currentAddress[12] ),
    .X(_07854_));
 sky130_fd_sc_hd__or2_1 _12943_ (.A(_07847_),
    .B(_07853_),
    .X(_07855_));
 sky130_fd_sc_hd__or4_1 _12944_ (.A(_07849_),
    .B(_07850_),
    .C(_07851_),
    .D(_07854_),
    .X(_07856_));
 sky130_fd_sc_hd__or3_1 _12945_ (.A(_07848_),
    .B(_07852_),
    .C(_07856_),
    .X(_07857_));
 sky130_fd_sc_hd__or4_2 _12946_ (.A(_07844_),
    .B(_07846_),
    .C(_07855_),
    .D(_07857_),
    .X(_07858_));
 sky130_fd_sc_hd__a22o_2 _12947_ (.A1(\jtag.managementAddress[16] ),
    .A2(net1307),
    .B1(net1256),
    .B2(\wbSRAMInterface.currentAddress[16] ),
    .X(_07859_));
 sky130_fd_sc_hd__or3_4 _12948_ (.A(\wbSRAMInterface.currentAddress[17] ),
    .B(\wbSRAMInterface.currentAddress[18] ),
    .C(\wbSRAMInterface.currentAddress[19] ),
    .X(_07860_));
 sky130_fd_sc_hd__or3_4 _12949_ (.A(\jtag.managementAddress[19] ),
    .B(\jtag.managementAddress[18] ),
    .C(\jtag.managementAddress[17] ),
    .X(_07861_));
 sky130_fd_sc_hd__a22o_4 _12950_ (.A1(net1256),
    .A2(_07860_),
    .B1(_07861_),
    .B2(net1307),
    .X(_07862_));
 sky130_fd_sc_hd__nor3b_4 _12951_ (.A(net1789),
    .B(_07862_),
    .C_N(_07859_),
    .Y(_07863_));
 sky130_fd_sc_hd__or3b_4 _12952_ (.A(net1789),
    .B(_07862_),
    .C_N(_07859_),
    .X(_07864_));
 sky130_fd_sc_hd__and2b_4 _12953_ (.A_N(\wbSRAMInterface.state[1] ),
    .B(\wbSRAMInterface.state[0] ),
    .X(_07865_));
 sky130_fd_sc_hd__nand2b_4 _12954_ (.A_N(\wbSRAMInterface.state[1] ),
    .B(\wbSRAMInterface.state[0] ),
    .Y(_07866_));
 sky130_fd_sc_hd__a31o_2 _12955_ (.A1(_07835_),
    .A2(_07841_),
    .A3(_07865_),
    .B1(net1369),
    .X(_07867_));
 sky130_fd_sc_hd__nand2_1 _12956_ (.A(_07863_),
    .B(_07867_),
    .Y(_07868_));
 sky130_fd_sc_hd__a22o_1 _12957_ (.A1(\jtag.managementAddress[5] ),
    .A2(net1306),
    .B1(net1256),
    .B2(\wbSRAMInterface.currentAddress[5] ),
    .X(_07869_));
 sky130_fd_sc_hd__a22o_2 _12958_ (.A1(\jtag.managementAddress[4] ),
    .A2(net1306),
    .B1(net1256),
    .B2(\wbSRAMInterface.currentAddress[4] ),
    .X(_07870_));
 sky130_fd_sc_hd__or2_1 _12959_ (.A(_07869_),
    .B(_07870_),
    .X(_07871_));
 sky130_fd_sc_hd__o21a_1 _12960_ (.A1(\wbSRAMInterface.currentAddress[0] ),
    .A2(\wbSRAMInterface.currentAddress[1] ),
    .B1(_07841_),
    .X(_07872_));
 sky130_fd_sc_hd__or2_1 _12961_ (.A(\jtag.managementAddress[1] ),
    .B(\jtag.managementAddress[0] ),
    .X(_07873_));
 sky130_fd_sc_hd__mux2_4 _12962_ (.A0(_07872_),
    .A1(_07873_),
    .S(_07836_),
    .X(_07874_));
 sky130_fd_sc_hd__or4_4 _12963_ (.A(_07858_),
    .B(_07868_),
    .C(_07871_),
    .D(_07874_),
    .X(_07875_));
 sky130_fd_sc_hd__a22o_4 _12964_ (.A1(\jtag.managementAddress[2] ),
    .A2(net1306),
    .B1(net1256),
    .B2(\wbSRAMInterface.currentAddress[2] ),
    .X(_07876_));
 sky130_fd_sc_hd__or3b_1 _12965_ (.A(_07875_),
    .B(_07876_),
    .C_N(_07843_),
    .X(_07877_));
 sky130_fd_sc_hd__nor3b_2 _12966_ (.A(net1791),
    .B(\core.management_pipeStartup ),
    .C_N(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__or4_1 _12967_ (.A(\core.csr.currentInstruction[15] ),
    .B(net1885),
    .C(\core.csr.currentInstruction[11] ),
    .D(\core.csr.currentInstruction[10] ),
    .X(_07879_));
 sky130_fd_sc_hd__or4_1 _12968_ (.A(\core.csr.currentInstruction[9] ),
    .B(\core.csr.currentInstruction[8] ),
    .C(\core.csr.currentInstruction[7] ),
    .D(_07879_),
    .X(_07880_));
 sky130_fd_sc_hd__or3_1 _12969_ (.A(\core.csr.currentInstruction[31] ),
    .B(\core.csr.currentInstruction[14] ),
    .C(\core.csr.currentInstruction[12] ),
    .X(_07881_));
 sky130_fd_sc_hd__or4b_1 _12970_ (.A(\core.csr.currentInstruction[23] ),
    .B(\core.csr.currentInstruction[22] ),
    .C(\core.csr.currentInstruction[20] ),
    .D_N(\core.csr.currentInstruction[21] ),
    .X(_07882_));
 sky130_fd_sc_hd__or3b_1 _12971_ (.A(\core.csr.currentInstruction[24] ),
    .B(_07882_),
    .C_N(\core.csr.currentInstruction[29] ),
    .X(_07883_));
 sky130_fd_sc_hd__or4_2 _12972_ (.A(\core.csr.currentInstruction[30] ),
    .B(_04492_),
    .C(_07881_),
    .D(_07883_),
    .X(_07884_));
 sky130_fd_sc_hd__or4_1 _12973_ (.A(\core.csr.currentInstruction[19] ),
    .B(\core.csr.currentInstruction[18] ),
    .C(\core.csr.currentInstruction[17] ),
    .D(\core.csr.currentInstruction[16] ),
    .X(_07885_));
 sky130_fd_sc_hd__or3b_4 _12974_ (.A(\core.csr.currentInstruction[25] ),
    .B(_07885_),
    .C_N(\core.csr.currentInstruction[28] ),
    .X(_07886_));
 sky130_fd_sc_hd__or4_1 _12975_ (.A(_04519_),
    .B(_07880_),
    .C(_07884_),
    .D(_07886_),
    .X(_07887_));
 sky130_fd_sc_hd__nor2_1 _12976_ (.A(_04504_),
    .B(_04521_),
    .Y(_07888_));
 sky130_fd_sc_hd__a41o_1 _12977_ (.A1(\core.csr.currentInstruction[3] ),
    .A2(\core.csr.currentInstruction[2] ),
    .A3(_04495_),
    .A4(_07888_),
    .B1(_07878_),
    .X(_07889_));
 sky130_fd_sc_hd__or3b_1 _12978_ (.A(_07492_),
    .B(_07889_),
    .C_N(_07887_),
    .X(_07890_));
 sky130_fd_sc_hd__inv_2 _12979_ (.A(_07890_),
    .Y(_07891_));
 sky130_fd_sc_hd__nand2_1 _12980_ (.A(net787),
    .B(_07891_),
    .Y(_07892_));
 sky130_fd_sc_hd__clkinv_2 _12981_ (.A(_07892_),
    .Y(_07893_));
 sky130_fd_sc_hd__and4_2 _12982_ (.A(\core.fetchProgramCounter[2] ),
    .B(net798),
    .C(_07433_),
    .D(_07891_),
    .X(_07894_));
 sky130_fd_sc_hd__and2_1 _12983_ (.A(\core.fetchProgramCounter[3] ),
    .B(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__and4_2 _12984_ (.A(\core.fetchProgramCounter[5] ),
    .B(\core.fetchProgramCounter[4] ),
    .C(\core.fetchProgramCounter[3] ),
    .D(_07894_),
    .X(_07896_));
 sky130_fd_sc_hd__nand2_1 _12985_ (.A(\core.fetchProgramCounter[6] ),
    .B(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__and4_4 _12986_ (.A(\core.fetchProgramCounter[8] ),
    .B(\core.fetchProgramCounter[7] ),
    .C(\core.fetchProgramCounter[6] ),
    .D(_07896_),
    .X(_07898_));
 sky130_fd_sc_hd__and3_1 _12987_ (.A(\core.fetchProgramCounter[10] ),
    .B(\core.fetchProgramCounter[9] ),
    .C(_07898_),
    .X(_07899_));
 sky130_fd_sc_hd__and3_1 _12988_ (.A(\core.fetchProgramCounter[13] ),
    .B(\core.fetchProgramCounter[12] ),
    .C(\core.fetchProgramCounter[11] ),
    .X(_07900_));
 sky130_fd_sc_hd__and4_1 _12989_ (.A(\core.fetchProgramCounter[17] ),
    .B(\core.fetchProgramCounter[16] ),
    .C(\core.fetchProgramCounter[15] ),
    .D(\core.fetchProgramCounter[14] ),
    .X(_07901_));
 sky130_fd_sc_hd__and3_1 _12990_ (.A(\core.fetchProgramCounter[10] ),
    .B(_07900_),
    .C(_07901_),
    .X(_07902_));
 sky130_fd_sc_hd__and4_2 _12991_ (.A(\core.fetchProgramCounter[18] ),
    .B(\core.fetchProgramCounter[9] ),
    .C(_07898_),
    .D(_07902_),
    .X(_07903_));
 sky130_fd_sc_hd__and2_2 _12992_ (.A(\core.fetchProgramCounter[19] ),
    .B(_07903_),
    .X(_07904_));
 sky130_fd_sc_hd__and4_4 _12993_ (.A(\core.fetchProgramCounter[21] ),
    .B(\core.fetchProgramCounter[20] ),
    .C(\core.fetchProgramCounter[19] ),
    .D(_07903_),
    .X(_07905_));
 sky130_fd_sc_hd__nand2_1 _12994_ (.A(\core.fetchProgramCounter[22] ),
    .B(_07905_),
    .Y(_07906_));
 sky130_fd_sc_hd__and4_2 _12995_ (.A(\core.fetchProgramCounter[24] ),
    .B(\core.fetchProgramCounter[23] ),
    .C(\core.fetchProgramCounter[22] ),
    .D(_07905_),
    .X(_07907_));
 sky130_fd_sc_hd__nand3_1 _12996_ (.A(\core.fetchProgramCounter[26] ),
    .B(\core.fetchProgramCounter[25] ),
    .C(_07907_),
    .Y(_07908_));
 sky130_fd_sc_hd__and4_2 _12997_ (.A(\core.fetchProgramCounter[27] ),
    .B(\core.fetchProgramCounter[26] ),
    .C(\core.fetchProgramCounter[25] ),
    .D(_07907_),
    .X(_07909_));
 sky130_fd_sc_hd__nand2_1 _12998_ (.A(\core.fetchProgramCounter[28] ),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__and3_1 _12999_ (.A(\core.fetchProgramCounter[29] ),
    .B(\core.fetchProgramCounter[28] ),
    .C(_07909_),
    .X(_07911_));
 sky130_fd_sc_hd__nand2_1 _13000_ (.A(\core.fetchProgramCounter[30] ),
    .B(_07911_),
    .Y(_07912_));
 sky130_fd_sc_hd__xnor2_1 _13001_ (.A(\core.fetchProgramCounter[31] ),
    .B(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__nor2_1 _13002_ (.A(net792),
    .B(_07913_),
    .Y(_07914_));
 sky130_fd_sc_hd__a21oi_1 _13003_ (.A1(\core.csr.trapReturnVector[31] ),
    .A2(net1177),
    .B1(net771),
    .Y(_07915_));
 sky130_fd_sc_hd__o31a_2 _13004_ (.A1(net1177),
    .A2(_07832_),
    .A3(_07914_),
    .B1(_07915_),
    .X(_07916_));
 sky130_fd_sc_hd__nand2_1 _13005_ (.A(\core.csr.traps.mtvec.csrReadData[30] ),
    .B(\core.csr.traps.mcause.csrReadData[28] ),
    .Y(_07917_));
 sky130_fd_sc_hd__or2_1 _13006_ (.A(\core.csr.traps.mtvec.csrReadData[30] ),
    .B(\core.csr.traps.mcause.csrReadData[28] ),
    .X(_07918_));
 sky130_fd_sc_hd__nor2_1 _13007_ (.A(\core.csr.traps.mtvec.csrReadData[29] ),
    .B(\core.csr.traps.mcause.csrReadData[27] ),
    .Y(_07919_));
 sky130_fd_sc_hd__nand2_1 _13008_ (.A(\core.csr.traps.mtvec.csrReadData[29] ),
    .B(\core.csr.traps.mcause.csrReadData[27] ),
    .Y(_07920_));
 sky130_fd_sc_hd__nor2_1 _13009_ (.A(\core.csr.traps.mtvec.csrReadData[28] ),
    .B(\core.csr.traps.mcause.csrReadData[26] ),
    .Y(_07921_));
 sky130_fd_sc_hd__nand2_1 _13010_ (.A(\core.csr.traps.mtvec.csrReadData[28] ),
    .B(\core.csr.traps.mcause.csrReadData[26] ),
    .Y(_07922_));
 sky130_fd_sc_hd__nand2_1 _13011_ (.A(\core.csr.traps.mtvec.csrReadData[27] ),
    .B(\core.csr.traps.mcause.csrReadData[25] ),
    .Y(_07923_));
 sky130_fd_sc_hd__or2_1 _13012_ (.A(\core.csr.traps.mtvec.csrReadData[27] ),
    .B(\core.csr.traps.mcause.csrReadData[25] ),
    .X(_07924_));
 sky130_fd_sc_hd__and2_2 _13013_ (.A(\core.csr.traps.mtvec.csrReadData[26] ),
    .B(\core.csr.traps.mcause.csrReadData[24] ),
    .X(_07925_));
 sky130_fd_sc_hd__nor2_1 _13014_ (.A(\core.csr.traps.mtvec.csrReadData[26] ),
    .B(\core.csr.traps.mcause.csrReadData[24] ),
    .Y(_07926_));
 sky130_fd_sc_hd__or2_4 _13015_ (.A(\core.csr.traps.mtvec.csrReadData[25] ),
    .B(\core.csr.traps.mcause.csrReadData[23] ),
    .X(_07927_));
 sky130_fd_sc_hd__nand2_2 _13016_ (.A(\core.csr.traps.mtvec.csrReadData[25] ),
    .B(\core.csr.traps.mcause.csrReadData[23] ),
    .Y(_07928_));
 sky130_fd_sc_hd__nor2_2 _13017_ (.A(\core.csr.traps.mtvec.csrReadData[24] ),
    .B(\core.csr.traps.mcause.csrReadData[22] ),
    .Y(_07929_));
 sky130_fd_sc_hd__nand2_2 _13018_ (.A(\core.csr.traps.mtvec.csrReadData[24] ),
    .B(\core.csr.traps.mcause.csrReadData[22] ),
    .Y(_07930_));
 sky130_fd_sc_hd__or2_2 _13019_ (.A(\core.csr.traps.mtvec.csrReadData[23] ),
    .B(\core.csr.traps.mcause.csrReadData[21] ),
    .X(_07931_));
 sky130_fd_sc_hd__nand2_1 _13020_ (.A(\core.csr.traps.mtvec.csrReadData[23] ),
    .B(\core.csr.traps.mcause.csrReadData[21] ),
    .Y(_07932_));
 sky130_fd_sc_hd__nor2_2 _13021_ (.A(\core.csr.traps.mtvec.csrReadData[22] ),
    .B(\core.csr.traps.mcause.csrReadData[20] ),
    .Y(_07933_));
 sky130_fd_sc_hd__nand2_2 _13022_ (.A(\core.csr.traps.mtvec.csrReadData[22] ),
    .B(\core.csr.traps.mcause.csrReadData[20] ),
    .Y(_07934_));
 sky130_fd_sc_hd__or2_2 _13023_ (.A(\core.csr.traps.mtvec.csrReadData[21] ),
    .B(\core.csr.traps.mcause.csrReadData[19] ),
    .X(_07935_));
 sky130_fd_sc_hd__nand2_1 _13024_ (.A(\core.csr.traps.mtvec.csrReadData[21] ),
    .B(\core.csr.traps.mcause.csrReadData[19] ),
    .Y(_07936_));
 sky130_fd_sc_hd__nor2_2 _13025_ (.A(\core.csr.traps.mtvec.csrReadData[20] ),
    .B(\core.csr.traps.mcause.csrReadData[18] ),
    .Y(_07937_));
 sky130_fd_sc_hd__nand2_2 _13026_ (.A(\core.csr.traps.mtvec.csrReadData[20] ),
    .B(\core.csr.traps.mcause.csrReadData[18] ),
    .Y(_07938_));
 sky130_fd_sc_hd__or2_2 _13027_ (.A(\core.csr.traps.mtvec.csrReadData[19] ),
    .B(\core.csr.traps.mcause.csrReadData[17] ),
    .X(_07939_));
 sky130_fd_sc_hd__nand2_1 _13028_ (.A(\core.csr.traps.mtvec.csrReadData[19] ),
    .B(\core.csr.traps.mcause.csrReadData[17] ),
    .Y(_07940_));
 sky130_fd_sc_hd__nor2_2 _13029_ (.A(\core.csr.traps.mtvec.csrReadData[18] ),
    .B(\core.csr.traps.mcause.csrReadData[16] ),
    .Y(_07941_));
 sky130_fd_sc_hd__nand2_2 _13030_ (.A(\core.csr.traps.mtvec.csrReadData[18] ),
    .B(\core.csr.traps.mcause.csrReadData[16] ),
    .Y(_07942_));
 sky130_fd_sc_hd__nor2_1 _13031_ (.A(\core.csr.traps.mtvec.csrReadData[16] ),
    .B(\core.csr.traps.mcause.csrReadData[14] ),
    .Y(_07943_));
 sky130_fd_sc_hd__nand2_1 _13032_ (.A(\core.csr.traps.mtvec.csrReadData[16] ),
    .B(\core.csr.traps.mcause.csrReadData[14] ),
    .Y(_07944_));
 sky130_fd_sc_hd__or2_4 _13033_ (.A(\core.csr.traps.mtvec.csrReadData[15] ),
    .B(\core.csr.traps.mcause.csrReadData[13] ),
    .X(_07945_));
 sky130_fd_sc_hd__nand2_1 _13034_ (.A(\core.csr.traps.mtvec.csrReadData[15] ),
    .B(\core.csr.traps.mcause.csrReadData[13] ),
    .Y(_07946_));
 sky130_fd_sc_hd__nor2_2 _13035_ (.A(\core.csr.traps.mtvec.csrReadData[14] ),
    .B(\core.csr.traps.mcause.csrReadData[12] ),
    .Y(_07947_));
 sky130_fd_sc_hd__nand2_2 _13036_ (.A(\core.csr.traps.mtvec.csrReadData[14] ),
    .B(\core.csr.traps.mcause.csrReadData[12] ),
    .Y(_07948_));
 sky130_fd_sc_hd__or2_2 _13037_ (.A(\core.csr.traps.mtvec.csrReadData[13] ),
    .B(\core.csr.traps.mcause.csrReadData[11] ),
    .X(_07949_));
 sky130_fd_sc_hd__nand2_1 _13038_ (.A(\core.csr.traps.mtvec.csrReadData[13] ),
    .B(\core.csr.traps.mcause.csrReadData[11] ),
    .Y(_07950_));
 sky130_fd_sc_hd__nor2_2 _13039_ (.A(\core.csr.traps.mtvec.csrReadData[12] ),
    .B(\core.csr.traps.mcause.csrReadData[10] ),
    .Y(_07951_));
 sky130_fd_sc_hd__nand2_2 _13040_ (.A(\core.csr.traps.mtvec.csrReadData[12] ),
    .B(\core.csr.traps.mcause.csrReadData[10] ),
    .Y(_07952_));
 sky130_fd_sc_hd__or2_2 _13041_ (.A(\core.csr.traps.mtvec.csrReadData[11] ),
    .B(\core.csr.traps.mcause.csrReadData[9] ),
    .X(_07953_));
 sky130_fd_sc_hd__nand2_1 _13042_ (.A(\core.csr.traps.mtvec.csrReadData[11] ),
    .B(\core.csr.traps.mcause.csrReadData[9] ),
    .Y(_07954_));
 sky130_fd_sc_hd__nor2_2 _13043_ (.A(\core.csr.traps.mtvec.csrReadData[10] ),
    .B(\core.csr.traps.mcause.csrReadData[8] ),
    .Y(_07955_));
 sky130_fd_sc_hd__nand2_2 _13044_ (.A(\core.csr.traps.mtvec.csrReadData[10] ),
    .B(\core.csr.traps.mcause.csrReadData[8] ),
    .Y(_07956_));
 sky130_fd_sc_hd__nor2_1 _13045_ (.A(\core.csr.traps.mtvec.csrReadData[9] ),
    .B(\core.csr.traps.mcause.csrReadData[7] ),
    .Y(_07957_));
 sky130_fd_sc_hd__and2_1 _13046_ (.A(\core.csr.traps.mtvec.csrReadData[9] ),
    .B(\core.csr.traps.mcause.csrReadData[7] ),
    .X(_07958_));
 sky130_fd_sc_hd__or2_2 _13047_ (.A(\core.csr.traps.mtvec.csrReadData[8] ),
    .B(\core.csr.traps.mcause.csrReadData[6] ),
    .X(_07959_));
 sky130_fd_sc_hd__nand2_1 _13048_ (.A(\core.csr.traps.mtvec.csrReadData[8] ),
    .B(\core.csr.traps.mcause.csrReadData[6] ),
    .Y(_07960_));
 sky130_fd_sc_hd__nand2_1 _13049_ (.A(\core.csr.traps.mtvec.csrReadData[7] ),
    .B(\core.csr.traps.mcause.csrReadData[5] ),
    .Y(_07961_));
 sky130_fd_sc_hd__or2_1 _13050_ (.A(\core.csr.traps.mtvec.csrReadData[7] ),
    .B(\core.csr.traps.mcause.csrReadData[5] ),
    .X(_07962_));
 sky130_fd_sc_hd__and2_1 _13051_ (.A(\core.csr.traps.mtvec.csrReadData[6] ),
    .B(\core.csr.traps.mcause.csrReadData[4] ),
    .X(_07963_));
 sky130_fd_sc_hd__nand2_1 _13052_ (.A(\core.csr.traps.mtvec.csrReadData[6] ),
    .B(\core.csr.traps.mcause.csrReadData[4] ),
    .Y(_07964_));
 sky130_fd_sc_hd__or2_1 _13053_ (.A(\core.csr.traps.mtvec.csrReadData[6] ),
    .B(\core.csr.traps.mcause.csrReadData[4] ),
    .X(_07965_));
 sky130_fd_sc_hd__or2_2 _13054_ (.A(\core.csr.traps.mtvec.csrReadData[5] ),
    .B(\core.csr.traps.mcause.csrReadData[3] ),
    .X(_07966_));
 sky130_fd_sc_hd__nand2_1 _13055_ (.A(\core.csr.traps.mtvec.csrReadData[5] ),
    .B(\core.csr.traps.mcause.csrReadData[3] ),
    .Y(_07967_));
 sky130_fd_sc_hd__nor2_1 _13056_ (.A(\core.csr.traps.mtvec.csrReadData[4] ),
    .B(\core.csr.traps.mcause.csrReadData[2] ),
    .Y(_07968_));
 sky130_fd_sc_hd__nand2_1 _13057_ (.A(\core.csr.traps.mtvec.csrReadData[4] ),
    .B(\core.csr.traps.mcause.csrReadData[2] ),
    .Y(_07969_));
 sky130_fd_sc_hd__nand2_1 _13058_ (.A(\core.csr.traps.mtvec.csrReadData[3] ),
    .B(\core.csr.traps.mcause.csrReadData[1] ),
    .Y(_07970_));
 sky130_fd_sc_hd__or2_1 _13059_ (.A(\core.csr.traps.mtvec.csrReadData[3] ),
    .B(\core.csr.traps.mcause.csrReadData[1] ),
    .X(_07971_));
 sky130_fd_sc_hd__and4_1 _13060_ (.A(\core.csr.traps.mtvec.csrReadData[2] ),
    .B(\core.csr.traps.mcause.csrReadData[0] ),
    .C(_07970_),
    .D(_07971_),
    .X(_07972_));
 sky130_fd_sc_hd__a21oi_2 _13061_ (.A1(\core.csr.traps.mtvec.csrReadData[3] ),
    .A2(\core.csr.traps.mcause.csrReadData[1] ),
    .B1(_07972_),
    .Y(_07973_));
 sky130_fd_sc_hd__o21ai_2 _13062_ (.A1(_07968_),
    .A2(_07973_),
    .B1(_07969_),
    .Y(_07974_));
 sky130_fd_sc_hd__a21o_1 _13063_ (.A1(\core.csr.traps.mtvec.csrReadData[5] ),
    .A2(\core.csr.traps.mcause.csrReadData[3] ),
    .B1(_07974_),
    .X(_07975_));
 sky130_fd_sc_hd__and4_2 _13064_ (.A(_07964_),
    .B(_07965_),
    .C(_07966_),
    .D(_07975_),
    .X(_07976_));
 sky130_fd_sc_hd__o211a_1 _13065_ (.A1(_07963_),
    .A2(_07976_),
    .B1(_07961_),
    .C1(_07962_),
    .X(_07977_));
 sky130_fd_sc_hd__a21o_2 _13066_ (.A1(\core.csr.traps.mtvec.csrReadData[7] ),
    .A2(\core.csr.traps.mcause.csrReadData[5] ),
    .B1(_07977_),
    .X(_07978_));
 sky130_fd_sc_hd__a21boi_4 _13067_ (.A1(_07959_),
    .A2(_07978_),
    .B1_N(_07960_),
    .Y(_07979_));
 sky130_fd_sc_hd__o21ba_2 _13068_ (.A1(_07957_),
    .A2(_07979_),
    .B1_N(_07958_),
    .X(_07980_));
 sky130_fd_sc_hd__o21ai_4 _13069_ (.A1(_07955_),
    .A2(_07980_),
    .B1(_07956_),
    .Y(_07981_));
 sky130_fd_sc_hd__a21boi_4 _13070_ (.A1(_07953_),
    .A2(_07981_),
    .B1_N(_07954_),
    .Y(_07982_));
 sky130_fd_sc_hd__o21ai_4 _13071_ (.A1(_07951_),
    .A2(_07982_),
    .B1(_07952_),
    .Y(_07983_));
 sky130_fd_sc_hd__a21boi_4 _13072_ (.A1(_07949_),
    .A2(_07983_),
    .B1_N(_07950_),
    .Y(_07984_));
 sky130_fd_sc_hd__o21ai_4 _13073_ (.A1(_07947_),
    .A2(_07984_),
    .B1(_07948_),
    .Y(_07985_));
 sky130_fd_sc_hd__a21boi_4 _13074_ (.A1(_07945_),
    .A2(_07985_),
    .B1_N(_07946_),
    .Y(_07986_));
 sky130_fd_sc_hd__o21ai_2 _13075_ (.A1(_07943_),
    .A2(_07986_),
    .B1(_07944_),
    .Y(_07987_));
 sky130_fd_sc_hd__a21o_1 _13076_ (.A1(\core.csr.traps.mtvec.csrReadData[17] ),
    .A2(\core.csr.traps.mcause.csrReadData[15] ),
    .B1(_07987_),
    .X(_07988_));
 sky130_fd_sc_hd__o21ai_4 _13077_ (.A1(\core.csr.traps.mtvec.csrReadData[17] ),
    .A2(\core.csr.traps.mcause.csrReadData[15] ),
    .B1(_07988_),
    .Y(_07989_));
 sky130_fd_sc_hd__o21ai_4 _13078_ (.A1(_07941_),
    .A2(_07989_),
    .B1(_07942_),
    .Y(_07990_));
 sky130_fd_sc_hd__a21boi_4 _13079_ (.A1(_07939_),
    .A2(_07990_),
    .B1_N(_07940_),
    .Y(_07991_));
 sky130_fd_sc_hd__o21ai_4 _13080_ (.A1(_07937_),
    .A2(_07991_),
    .B1(_07938_),
    .Y(_07992_));
 sky130_fd_sc_hd__a21boi_4 _13081_ (.A1(_07935_),
    .A2(_07992_),
    .B1_N(_07936_),
    .Y(_07993_));
 sky130_fd_sc_hd__o21ai_4 _13082_ (.A1(_07933_),
    .A2(_07993_),
    .B1(_07934_),
    .Y(_07994_));
 sky130_fd_sc_hd__a21boi_4 _13083_ (.A1(_07931_),
    .A2(_07994_),
    .B1_N(_07932_),
    .Y(_07995_));
 sky130_fd_sc_hd__o21ai_4 _13084_ (.A1(_07929_),
    .A2(_07995_),
    .B1(_07930_),
    .Y(_07996_));
 sky130_fd_sc_hd__a21boi_2 _13085_ (.A1(_07927_),
    .A2(_07996_),
    .B1_N(_07928_),
    .Y(_07997_));
 sky130_fd_sc_hd__nor3_2 _13086_ (.A(_07925_),
    .B(_07926_),
    .C(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__o211a_1 _13087_ (.A1(_07925_),
    .A2(_07998_),
    .B1(_07923_),
    .C1(_07924_),
    .X(_07999_));
 sky130_fd_sc_hd__a21oi_2 _13088_ (.A1(\core.csr.traps.mtvec.csrReadData[27] ),
    .A2(\core.csr.traps.mcause.csrReadData[25] ),
    .B1(_07999_),
    .Y(_08000_));
 sky130_fd_sc_hd__o21a_1 _13089_ (.A1(_07921_),
    .A2(_08000_),
    .B1(_07922_),
    .X(_08001_));
 sky130_fd_sc_hd__o21ai_2 _13090_ (.A1(_07919_),
    .A2(_08001_),
    .B1(_07920_),
    .Y(_08002_));
 sky130_fd_sc_hd__and3_1 _13091_ (.A(_07917_),
    .B(_07918_),
    .C(_08002_),
    .X(_08003_));
 sky130_fd_sc_hd__a21o_1 _13092_ (.A1(\core.csr.traps.mtvec.csrReadData[30] ),
    .A2(\core.csr.traps.mcause.csrReadData[28] ),
    .B1(_08003_),
    .X(_08004_));
 sky130_fd_sc_hd__or3b_4 _13093_ (.A(\core.csr.traps.mtvec.csrReadData[1] ),
    .B(_07468_),
    .C_N(\core.csr.traps.mtvec.csrReadData[0] ),
    .X(_08005_));
 sky130_fd_sc_hd__a21oi_1 _13094_ (.A1(\core.csr.traps.mcause.csrReadData[29] ),
    .A2(_08004_),
    .B1(net1220),
    .Y(_08006_));
 sky130_fd_sc_hd__o21a_1 _13095_ (.A1(\core.csr.traps.mcause.csrReadData[29] ),
    .A2(_08004_),
    .B1(_08006_),
    .X(_08007_));
 sky130_fd_sc_hd__xnor2_2 _13096_ (.A(\core.csr.traps.mtvec.csrReadData[31] ),
    .B(_08007_),
    .Y(_08008_));
 sky130_fd_sc_hd__and2_1 _13097_ (.A(net771),
    .B(_08008_),
    .X(_08009_));
 sky130_fd_sc_hd__o21ai_4 _13098_ (.A1(_07916_),
    .A2(_08009_),
    .B1(net1767),
    .Y(_08010_));
 sky130_fd_sc_hd__o21a_2 _13099_ (.A1(net1767),
    .A2(\core.fetchProgramCounter[31] ),
    .B1(net1889),
    .X(_08011_));
 sky130_fd_sc_hd__and2_1 _13100_ (.A(_08010_),
    .B(_08011_),
    .X(_08012_));
 sky130_fd_sc_hd__a21oi_1 _13101_ (.A1(_07917_),
    .A2(_07918_),
    .B1(_08002_),
    .Y(_08013_));
 sky130_fd_sc_hd__nand2_1 _13102_ (.A(\core.csr.traps.mtvec.csrReadData[30] ),
    .B(net1219),
    .Y(_08014_));
 sky130_fd_sc_hd__o311a_1 _13103_ (.A1(_08003_),
    .A2(net1219),
    .A3(_08013_),
    .B1(_08014_),
    .C1(net769),
    .X(_08015_));
 sky130_fd_sc_hd__or2_1 _13104_ (.A(\core.fetchProgramCounter[30] ),
    .B(_07911_),
    .X(_08016_));
 sky130_fd_sc_hd__a21o_1 _13105_ (.A1(_07912_),
    .A2(_08016_),
    .B1(net792),
    .X(_08017_));
 sky130_fd_sc_hd__nand4_1 _13106_ (.A(_07539_),
    .B(_07817_),
    .C(_07822_),
    .D(_07824_),
    .Y(_08018_));
 sky130_fd_sc_hd__nor2_2 _13107_ (.A(_07402_),
    .B(_07422_),
    .Y(_08019_));
 sky130_fd_sc_hd__a31o_1 _13108_ (.A1(_07825_),
    .A2(_08018_),
    .A3(_08019_),
    .B1(net788),
    .X(_08020_));
 sky130_fd_sc_hd__a21o_1 _13109_ (.A1(\core.csr.trapReturnVector[30] ),
    .A2(net1177),
    .B1(net771),
    .X(_08021_));
 sky130_fd_sc_hd__a21oi_1 _13110_ (.A1(_08017_),
    .A2(_08020_),
    .B1(_08021_),
    .Y(_08022_));
 sky130_fd_sc_hd__o21ai_1 _13111_ (.A1(_08015_),
    .A2(_08022_),
    .B1(net1767),
    .Y(_08023_));
 sky130_fd_sc_hd__o211a_2 _13112_ (.A1(net1767),
    .A2(\core.fetchProgramCounter[30] ),
    .B1(net1888),
    .C1(_08023_),
    .X(_08024_));
 sky130_fd_sc_hd__a21oi_4 _13113_ (.A1(_08010_),
    .A2(_08011_),
    .B1(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__or2_1 _13114_ (.A(\core.fetchProgramCounter[28] ),
    .B(_07909_),
    .X(_08026_));
 sky130_fd_sc_hd__a21o_1 _13115_ (.A1(_07910_),
    .A2(_08026_),
    .B1(net792),
    .X(_08027_));
 sky130_fd_sc_hd__nand3_1 _13116_ (.A(_07809_),
    .B(_07812_),
    .C(_07820_),
    .Y(_08028_));
 sky130_fd_sc_hd__a31o_1 _13117_ (.A1(_07821_),
    .A2(_08019_),
    .A3(_08028_),
    .B1(net788),
    .X(_08029_));
 sky130_fd_sc_hd__a21o_1 _13118_ (.A1(\core.csr.trapReturnVector[28] ),
    .A2(net1177),
    .B1(net771),
    .X(_08030_));
 sky130_fd_sc_hd__a21o_1 _13119_ (.A1(_08027_),
    .A2(_08029_),
    .B1(_08030_),
    .X(_08031_));
 sky130_fd_sc_hd__nand2b_1 _13120_ (.A_N(_07921_),
    .B(_07922_),
    .Y(_08032_));
 sky130_fd_sc_hd__xnor2_1 _13121_ (.A(_08000_),
    .B(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__nor2_1 _13122_ (.A(net1220),
    .B(_08033_),
    .Y(_08034_));
 sky130_fd_sc_hd__a211o_1 _13123_ (.A1(\core.csr.traps.mtvec.csrReadData[28] ),
    .A2(net1220),
    .B1(_08034_),
    .C1(net766),
    .X(_08035_));
 sky130_fd_sc_hd__and2_1 _13124_ (.A(net1766),
    .B(_08035_),
    .X(_08036_));
 sky130_fd_sc_hd__a22oi_4 _13125_ (.A1(net1760),
    .A2(\core.fetchProgramCounter[28] ),
    .B1(_08031_),
    .B2(_08036_),
    .Y(_08037_));
 sky130_fd_sc_hd__nor2_1 _13126_ (.A(net1969),
    .B(_08037_),
    .Y(_08038_));
 sky130_fd_sc_hd__a21oi_1 _13127_ (.A1(\core.fetchProgramCounter[28] ),
    .A2(_07909_),
    .B1(\core.fetchProgramCounter[29] ),
    .Y(_08039_));
 sky130_fd_sc_hd__o21a_1 _13128_ (.A1(_07911_),
    .A2(_08039_),
    .B1(net797),
    .X(_08040_));
 sky130_fd_sc_hd__a21oi_1 _13129_ (.A1(_07817_),
    .A2(_07821_),
    .B1(_07541_),
    .Y(_08041_));
 sky130_fd_sc_hd__a31o_1 _13130_ (.A1(_07541_),
    .A2(_07817_),
    .A3(_07821_),
    .B1(_07402_),
    .X(_08042_));
 sky130_fd_sc_hd__o31a_1 _13131_ (.A1(net1177),
    .A2(_08041_),
    .A3(_08042_),
    .B1(_07439_),
    .X(_08043_));
 sky130_fd_sc_hd__a21oi_1 _13132_ (.A1(\core.csr.trapReturnVector[29] ),
    .A2(net1178),
    .B1(net772),
    .Y(_08044_));
 sky130_fd_sc_hd__o21ai_1 _13133_ (.A1(_08040_),
    .A2(_08043_),
    .B1(_08044_),
    .Y(_08045_));
 sky130_fd_sc_hd__nand2b_1 _13134_ (.A_N(_07919_),
    .B(_07920_),
    .Y(_08046_));
 sky130_fd_sc_hd__nor2_1 _13135_ (.A(_08001_),
    .B(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__a21o_1 _13136_ (.A1(_08001_),
    .A2(_08046_),
    .B1(net1221),
    .X(_08048_));
 sky130_fd_sc_hd__a2bb2o_1 _13137_ (.A1_N(_08047_),
    .A2_N(_08048_),
    .B1(\core.csr.traps.mtvec.csrReadData[29] ),
    .B2(net1221),
    .X(_08049_));
 sky130_fd_sc_hd__o211a_1 _13138_ (.A1(net766),
    .A2(_08049_),
    .B1(_08045_),
    .C1(net1768),
    .X(_08050_));
 sky130_fd_sc_hd__and2_1 _13139_ (.A(net1760),
    .B(\core.fetchProgramCounter[29] ),
    .X(_08051_));
 sky130_fd_sc_hd__or2_4 _13140_ (.A(\core.pipe0_fetch.instructionCached ),
    .B(_07892_),
    .X(_08052_));
 sky130_fd_sc_hd__o21a_2 _13141_ (.A1(_08050_),
    .A2(_08051_),
    .B1(net1891),
    .X(_08053_));
 sky130_fd_sc_hd__and4bb_4 _13142_ (.A_N(_08053_),
    .B_N(_08052_),
    .C(_08038_),
    .D(_08025_),
    .X(_00577_));
 sky130_fd_sc_hd__nor2_2 _13143_ (.A(_06134_),
    .B(_07473_),
    .Y(_08054_));
 sky130_fd_sc_hd__a311o_2 _13144_ (.A1(_06136_),
    .A2(net933),
    .A3(_06227_),
    .B1(_06134_),
    .C1(_06050_),
    .X(_08055_));
 sky130_fd_sc_hd__nand2_2 _13145_ (.A(_06052_),
    .B(_08055_),
    .Y(_08056_));
 sky130_fd_sc_hd__a31o_4 _13146_ (.A1(_05967_),
    .A2(_06052_),
    .A3(_08055_),
    .B1(_05966_),
    .X(_08057_));
 sky130_fd_sc_hd__a21o_4 _13147_ (.A1(_05882_),
    .A2(_08057_),
    .B1(_05881_),
    .X(_08058_));
 sky130_fd_sc_hd__a21oi_4 _13148_ (.A1(_05798_),
    .A2(_08058_),
    .B1(_05796_),
    .Y(_08059_));
 sky130_fd_sc_hd__a211o_2 _13149_ (.A1(_05798_),
    .A2(_08058_),
    .B1(_05711_),
    .C1(_05796_),
    .X(_08060_));
 sky130_fd_sc_hd__nand2_2 _13150_ (.A(_05712_),
    .B(_08060_),
    .Y(_08061_));
 sky130_fd_sc_hd__a31o_4 _13151_ (.A1(_05632_),
    .A2(_05712_),
    .A3(_08060_),
    .B1(_05630_),
    .X(_08062_));
 sky130_fd_sc_hd__a21o_4 _13152_ (.A1(_06314_),
    .A2(_08062_),
    .B1(_06312_),
    .X(_08063_));
 sky130_fd_sc_hd__a21oi_4 _13153_ (.A1(_05551_),
    .A2(_08063_),
    .B1(_05550_),
    .Y(_08064_));
 sky130_fd_sc_hd__a211o_2 _13154_ (.A1(_05551_),
    .A2(_08063_),
    .B1(_05453_),
    .C1(_05550_),
    .X(_08065_));
 sky130_fd_sc_hd__nand2_2 _13155_ (.A(_05454_),
    .B(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__a32o_4 _13156_ (.A1(_05366_),
    .A2(_05454_),
    .A3(_08065_),
    .B1(_05364_),
    .B2(_05330_),
    .X(_08067_));
 sky130_fd_sc_hd__a21bo_4 _13157_ (.A1(_05024_),
    .A2(_08067_),
    .B1_N(_05025_),
    .X(_08068_));
 sky130_fd_sc_hd__a21bo_4 _13158_ (.A1(_05109_),
    .A2(_08068_),
    .B1_N(_05110_),
    .X(_08069_));
 sky130_fd_sc_hd__a21bo_4 _13159_ (.A1(_05280_),
    .A2(_08069_),
    .B1_N(_05278_),
    .X(_08070_));
 sky130_fd_sc_hd__a21oi_4 _13160_ (.A1(_05192_),
    .A2(_08070_),
    .B1(_05189_),
    .Y(_08071_));
 sky130_fd_sc_hd__a211o_2 _13161_ (.A1(_05192_),
    .A2(_08070_),
    .B1(_06487_),
    .C1(_05189_),
    .X(_08072_));
 sky130_fd_sc_hd__nand2_2 _13162_ (.A(_06486_),
    .B(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__a31o_2 _13163_ (.A1(_06407_),
    .A2(_06486_),
    .A3(_08072_),
    .B1(_06409_),
    .X(_08074_));
 sky130_fd_sc_hd__a311o_1 _13164_ (.A1(_06407_),
    .A2(_06486_),
    .A3(_08072_),
    .B1(_06642_),
    .C1(_06409_),
    .X(_08075_));
 sky130_fd_sc_hd__and2_2 _13165_ (.A(_06640_),
    .B(_08075_),
    .X(_08076_));
 sky130_fd_sc_hd__and3_2 _13166_ (.A(_06564_),
    .B(_06640_),
    .C(_08075_),
    .X(_08077_));
 sky130_fd_sc_hd__or2_4 _13167_ (.A(_06563_),
    .B(_08077_),
    .X(_08078_));
 sky130_fd_sc_hd__o31ai_4 _13168_ (.A1(_06563_),
    .A2(_06655_),
    .A3(_08077_),
    .B1(_06653_),
    .Y(_08079_));
 sky130_fd_sc_hd__a21boi_4 _13169_ (.A1(_04852_),
    .A2(_08079_),
    .B1_N(_04851_),
    .Y(_08080_));
 sky130_fd_sc_hd__a21o_4 _13170_ (.A1(_04773_),
    .A2(_08080_),
    .B1(_04774_),
    .X(_08081_));
 sky130_fd_sc_hd__a21oi_4 _13171_ (.A1(_04694_),
    .A2(_08081_),
    .B1(_04696_),
    .Y(_08082_));
 sky130_fd_sc_hd__o21bai_4 _13172_ (.A1(_06792_),
    .A2(_08082_),
    .B1_N(_06790_),
    .Y(_08083_));
 sky130_fd_sc_hd__a21oi_4 _13173_ (.A1(_06869_),
    .A2(_08083_),
    .B1(_06868_),
    .Y(_08084_));
 sky130_fd_sc_hd__o21a_4 _13174_ (.A1(_07022_),
    .A2(_08084_),
    .B1(_07023_),
    .X(_08085_));
 sky130_fd_sc_hd__o21a_4 _13175_ (.A1(_06947_),
    .A2(_08085_),
    .B1(_06948_),
    .X(_08086_));
 sky130_fd_sc_hd__a21oi_4 _13176_ (.A1(_07111_),
    .A2(_08086_),
    .B1(_07110_),
    .Y(_08087_));
 sky130_fd_sc_hd__a21oi_4 _13177_ (.A1(_07194_),
    .A2(_08087_),
    .B1(_07195_),
    .Y(_08088_));
 sky130_fd_sc_hd__xnor2_4 _13178_ (.A(_07350_),
    .B(_08088_),
    .Y(_08089_));
 sky130_fd_sc_hd__o21bai_4 _13179_ (.A1(_07351_),
    .A2(_08088_),
    .B1_N(_07349_),
    .Y(_08090_));
 sky130_fd_sc_hd__xnor2_4 _13180_ (.A(_07360_),
    .B(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__nor2_1 _13181_ (.A(_08089_),
    .B(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__xnor2_4 _13182_ (.A(_07196_),
    .B(_08087_),
    .Y(_08093_));
 sky130_fd_sc_hd__xnor2_4 _13183_ (.A(_07113_),
    .B(_08086_),
    .Y(_08094_));
 sky130_fd_sc_hd__and2_1 _13184_ (.A(net1241),
    .B(_07481_),
    .X(_08095_));
 sky130_fd_sc_hd__nand2_8 _13185_ (.A(net1241),
    .B(_07481_),
    .Y(_08096_));
 sky130_fd_sc_hd__or2_4 _13186_ (.A(\core.memoryOperationCompleted ),
    .B(_08096_),
    .X(_08097_));
 sky130_fd_sc_hd__nor2_1 _13187_ (.A(_08092_),
    .B(_08096_),
    .Y(_08098_));
 sky130_fd_sc_hd__and4b_4 _13188_ (.A_N(\core.memoryOperationCompleted ),
    .B(_08092_),
    .C(_08093_),
    .D(net807),
    .X(_08099_));
 sky130_fd_sc_hd__nand2_8 _13189_ (.A(net765),
    .B(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__nand2b_4 _13190_ (.A_N(net727),
    .B(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__and2_1 _13191_ (.A(_07505_),
    .B(_08101_),
    .X(net333));
 sky130_fd_sc_hd__nor2_8 _13192_ (.A(net1851),
    .B(_07498_),
    .Y(net444));
 sky130_fd_sc_hd__nor2_2 _13193_ (.A(net1730),
    .B(_07498_),
    .Y(net443));
 sky130_fd_sc_hd__nand2b_1 _13194_ (.A_N(_07929_),
    .B(_07930_),
    .Y(_08102_));
 sky130_fd_sc_hd__nor2_1 _13195_ (.A(_07995_),
    .B(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__a211o_1 _13196_ (.A1(_07995_),
    .A2(_08102_),
    .B1(_08103_),
    .C1(net1219),
    .X(_08104_));
 sky130_fd_sc_hd__nand2_1 _13197_ (.A(\core.csr.traps.mtvec.csrReadData[24] ),
    .B(net1219),
    .Y(_08105_));
 sky130_fd_sc_hd__a21boi_1 _13198_ (.A1(_07774_),
    .A2(_07782_),
    .B1_N(_07790_),
    .Y(_08106_));
 sky130_fd_sc_hd__xnor2_1 _13199_ (.A(_07783_),
    .B(_07790_),
    .Y(_08107_));
 sky130_fd_sc_hd__a21oi_1 _13200_ (.A1(\core.csr.trapReturnVector[24] ),
    .A2(net1177),
    .B1(net770),
    .Y(_08108_));
 sky130_fd_sc_hd__a31oi_1 _13201_ (.A1(\core.fetchProgramCounter[23] ),
    .A2(\core.fetchProgramCounter[22] ),
    .A3(_07905_),
    .B1(\core.fetchProgramCounter[24] ),
    .Y(_08109_));
 sky130_fd_sc_hd__o21a_1 _13202_ (.A1(_07907_),
    .A2(_08109_),
    .B1(net797),
    .X(_08110_));
 sky130_fd_sc_hd__a311o_2 _13203_ (.A1(net792),
    .A2(_07403_),
    .A3(_08107_),
    .B1(_08110_),
    .C1(net1178),
    .X(_08111_));
 sky130_fd_sc_hd__a32o_1 _13204_ (.A1(net770),
    .A2(_08104_),
    .A3(_08105_),
    .B1(_08108_),
    .B2(_08111_),
    .X(_08112_));
 sky130_fd_sc_hd__nand2_1 _13205_ (.A(net1766),
    .B(_08112_),
    .Y(_08113_));
 sky130_fd_sc_hd__o211a_4 _13206_ (.A1(net1766),
    .A2(\core.fetchProgramCounter[24] ),
    .B1(net1894),
    .C1(_08113_),
    .X(_08114_));
 sky130_fd_sc_hd__a21oi_1 _13207_ (.A1(_07774_),
    .A2(_07782_),
    .B1(_07807_),
    .Y(_08115_));
 sky130_fd_sc_hd__o21ai_2 _13208_ (.A1(_07810_),
    .A2(_08115_),
    .B1(_07806_),
    .Y(_08116_));
 sky130_fd_sc_hd__nand3_1 _13209_ (.A(_07795_),
    .B(_07804_),
    .C(_08116_),
    .Y(_08117_));
 sky130_fd_sc_hd__a21o_1 _13210_ (.A1(_07804_),
    .A2(_08116_),
    .B1(_07795_),
    .X(_08118_));
 sky130_fd_sc_hd__a31o_1 _13211_ (.A1(\core.fetchProgramCounter[26] ),
    .A2(\core.fetchProgramCounter[25] ),
    .A3(_07907_),
    .B1(\core.fetchProgramCounter[27] ),
    .X(_08119_));
 sky130_fd_sc_hd__and3b_1 _13212_ (.A_N(_07909_),
    .B(_08119_),
    .C(net788),
    .X(_08120_));
 sky130_fd_sc_hd__a211o_1 _13213_ (.A1(\core.csr.trapReturnVector[27] ),
    .A2(net1178),
    .B1(_08120_),
    .C1(net772),
    .X(_08121_));
 sky130_fd_sc_hd__a31o_1 _13214_ (.A1(net792),
    .A2(_08117_),
    .A3(_08118_),
    .B1(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__a211o_1 _13215_ (.A1(_07923_),
    .A2(_07924_),
    .B1(_07925_),
    .C1(_07998_),
    .X(_08123_));
 sky130_fd_sc_hd__nor2_1 _13216_ (.A(_07999_),
    .B(net1220),
    .Y(_08124_));
 sky130_fd_sc_hd__a221o_2 _13217_ (.A1(\core.csr.traps.mtvec.csrReadData[27] ),
    .A2(net1220),
    .B1(_08123_),
    .B2(_08124_),
    .C1(net766),
    .X(_08125_));
 sky130_fd_sc_hd__nand3_1 _13218_ (.A(net1768),
    .B(_08122_),
    .C(_08125_),
    .Y(_08126_));
 sky130_fd_sc_hd__a21boi_2 _13219_ (.A1(net1760),
    .A2(\core.fetchProgramCounter[27] ),
    .B1_N(_08126_),
    .Y(_08127_));
 sky130_fd_sc_hd__clkinv_2 _13220_ (.A(_08127_),
    .Y(_08128_));
 sky130_fd_sc_hd__or3_1 _13221_ (.A(_07806_),
    .B(_07810_),
    .C(_08115_),
    .X(_08129_));
 sky130_fd_sc_hd__a21o_1 _13222_ (.A1(\core.fetchProgramCounter[25] ),
    .A2(_07907_),
    .B1(\core.fetchProgramCounter[26] ),
    .X(_08130_));
 sky130_fd_sc_hd__a21o_1 _13223_ (.A1(\core.csr.trapReturnVector[26] ),
    .A2(net1178),
    .B1(net771),
    .X(_08131_));
 sky130_fd_sc_hd__a31o_1 _13224_ (.A1(net788),
    .A2(_07908_),
    .A3(_08130_),
    .B1(_08131_),
    .X(_08132_));
 sky130_fd_sc_hd__a31o_1 _13225_ (.A1(net793),
    .A2(_08116_),
    .A3(_08129_),
    .B1(_08132_),
    .X(_08133_));
 sky130_fd_sc_hd__o21ai_1 _13226_ (.A1(_07925_),
    .A2(_07926_),
    .B1(_07997_),
    .Y(_08134_));
 sky130_fd_sc_hd__nor2_1 _13227_ (.A(_07998_),
    .B(net1220),
    .Y(_08135_));
 sky130_fd_sc_hd__a221o_1 _13228_ (.A1(\core.csr.traps.mtvec.csrReadData[26] ),
    .A2(net1219),
    .B1(_08134_),
    .B2(_08135_),
    .C1(net766),
    .X(_08136_));
 sky130_fd_sc_hd__and3_1 _13229_ (.A(net1768),
    .B(_08133_),
    .C(_08136_),
    .X(_08137_));
 sky130_fd_sc_hd__a21o_2 _13230_ (.A1(net1760),
    .A2(\core.fetchProgramCounter[26] ),
    .B1(_08137_),
    .X(_08138_));
 sky130_fd_sc_hd__xor2_1 _13231_ (.A(\core.fetchProgramCounter[25] ),
    .B(_07907_),
    .X(_08139_));
 sky130_fd_sc_hd__a221o_1 _13232_ (.A1(\core.csr.trapReturnVector[25] ),
    .A2(net1178),
    .B1(net788),
    .B2(_08139_),
    .C1(net772),
    .X(_08140_));
 sky130_fd_sc_hd__or3_1 _13233_ (.A(_07788_),
    .B(_07799_),
    .C(_08106_),
    .X(_08141_));
 sky130_fd_sc_hd__o21ai_1 _13234_ (.A1(_07788_),
    .A2(_08106_),
    .B1(_07799_),
    .Y(_08142_));
 sky130_fd_sc_hd__a31o_1 _13235_ (.A1(net792),
    .A2(_08141_),
    .A3(_08142_),
    .B1(_08140_),
    .X(_08143_));
 sky130_fd_sc_hd__a21oi_2 _13236_ (.A1(_07927_),
    .A2(_07928_),
    .B1(_07996_),
    .Y(_08144_));
 sky130_fd_sc_hd__a311oi_4 _13237_ (.A1(_07927_),
    .A2(_07928_),
    .A3(_07996_),
    .B1(net1219),
    .C1(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__a211o_1 _13238_ (.A1(\core.csr.traps.mtvec.csrReadData[25] ),
    .A2(net1221),
    .B1(_08145_),
    .C1(net766),
    .X(_08146_));
 sky130_fd_sc_hd__and3_1 _13239_ (.A(net1768),
    .B(_08143_),
    .C(_08146_),
    .X(_08147_));
 sky130_fd_sc_hd__a21o_2 _13240_ (.A1(net1760),
    .A2(\core.fetchProgramCounter[25] ),
    .B1(_08147_),
    .X(_08148_));
 sky130_fd_sc_hd__o21a_1 _13241_ (.A1(_08138_),
    .A2(_08148_),
    .B1(net1899),
    .X(_08149_));
 sky130_fd_sc_hd__or4_2 _13242_ (.A(_08038_),
    .B(_08052_),
    .C(_08114_),
    .D(_08149_),
    .X(_08150_));
 sky130_fd_sc_hd__a211oi_4 _13243_ (.A1(net1900),
    .A2(_08128_),
    .B1(_08150_),
    .C1(_08053_),
    .Y(_08151_));
 sky130_fd_sc_hd__and2_4 _13244_ (.A(_08025_),
    .B(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__nand2_1 _13245_ (.A(_08025_),
    .B(_08151_),
    .Y(_08153_));
 sky130_fd_sc_hd__a21o_1 _13246_ (.A1(_07704_),
    .A2(_07710_),
    .B1(_07772_),
    .X(_08154_));
 sky130_fd_sc_hd__a211o_1 _13247_ (.A1(_07704_),
    .A2(_07710_),
    .B1(_07765_),
    .C1(_07772_),
    .X(_08155_));
 sky130_fd_sc_hd__or2_2 _13248_ (.A(_07754_),
    .B(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__a21oi_1 _13249_ (.A1(_07778_),
    .A2(_08156_),
    .B1(_07727_),
    .Y(_08157_));
 sky130_fd_sc_hd__a21o_2 _13250_ (.A1(_07778_),
    .A2(_08156_),
    .B1(_07727_),
    .X(_08158_));
 sky130_fd_sc_hd__nor2_2 _13251_ (.A(_07715_),
    .B(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__o21ai_4 _13252_ (.A1(_07779_),
    .A2(_08159_),
    .B1(_07721_),
    .Y(_08160_));
 sky130_fd_sc_hd__and3_1 _13253_ (.A(_07719_),
    .B(_07732_),
    .C(_08160_),
    .X(_08161_));
 sky130_fd_sc_hd__a21oi_1 _13254_ (.A1(_07719_),
    .A2(_08160_),
    .B1(_07732_),
    .Y(_08162_));
 sky130_fd_sc_hd__xnor2_1 _13255_ (.A(\core.fetchProgramCounter[23] ),
    .B(_07906_),
    .Y(_08163_));
 sky130_fd_sc_hd__a221oi_2 _13256_ (.A1(\core.csr.trapReturnVector[23] ),
    .A2(net1177),
    .B1(net788),
    .B2(_08163_),
    .C1(net771),
    .Y(_08164_));
 sky130_fd_sc_hd__o31a_2 _13257_ (.A1(net797),
    .A2(_08161_),
    .A3(_08162_),
    .B1(_08164_),
    .X(_08165_));
 sky130_fd_sc_hd__and3_1 _13258_ (.A(_07931_),
    .B(_07932_),
    .C(_07994_),
    .X(_08166_));
 sky130_fd_sc_hd__a21oi_1 _13259_ (.A1(_07931_),
    .A2(_07932_),
    .B1(_07994_),
    .Y(_08167_));
 sky130_fd_sc_hd__nand2_1 _13260_ (.A(\core.csr.traps.mtvec.csrReadData[23] ),
    .B(net1219),
    .Y(_08168_));
 sky130_fd_sc_hd__o311a_2 _13261_ (.A1(net1219),
    .A2(_08166_),
    .A3(_08167_),
    .B1(_08168_),
    .C1(net769),
    .X(_08169_));
 sky130_fd_sc_hd__o21ai_2 _13262_ (.A1(_08165_),
    .A2(_08169_),
    .B1(net1766),
    .Y(_08170_));
 sky130_fd_sc_hd__o211a_4 _13263_ (.A1(net1766),
    .A2(\core.fetchProgramCounter[23] ),
    .B1(net1894),
    .C1(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__and3_1 _13264_ (.A(_07715_),
    .B(_07726_),
    .C(_08158_),
    .X(_08172_));
 sky130_fd_sc_hd__a21oi_1 _13265_ (.A1(_07726_),
    .A2(_08158_),
    .B1(_07715_),
    .Y(_08173_));
 sky130_fd_sc_hd__a21oi_2 _13266_ (.A1(\core.fetchProgramCounter[20] ),
    .A2(_07904_),
    .B1(\core.fetchProgramCounter[21] ),
    .Y(_08174_));
 sky130_fd_sc_hd__a21oi_1 _13267_ (.A1(\core.csr.trapReturnVector[21] ),
    .A2(net1177),
    .B1(net771),
    .Y(_08175_));
 sky130_fd_sc_hd__o31a_1 _13268_ (.A1(_07439_),
    .A2(_07905_),
    .A3(_08174_),
    .B1(_08175_),
    .X(_08176_));
 sky130_fd_sc_hd__o31a_1 _13269_ (.A1(net797),
    .A2(_08172_),
    .A3(_08173_),
    .B1(_08176_),
    .X(_08177_));
 sky130_fd_sc_hd__and3_1 _13270_ (.A(_07935_),
    .B(_07936_),
    .C(_07992_),
    .X(_08178_));
 sky130_fd_sc_hd__a21oi_1 _13271_ (.A1(_07935_),
    .A2(_07936_),
    .B1(_07992_),
    .Y(_08179_));
 sky130_fd_sc_hd__nand2_1 _13272_ (.A(\core.csr.traps.mtvec.csrReadData[21] ),
    .B(net1220),
    .Y(_08180_));
 sky130_fd_sc_hd__o311a_1 _13273_ (.A1(net1220),
    .A2(_08178_),
    .A3(_08179_),
    .B1(_08180_),
    .C1(net773),
    .X(_08181_));
 sky130_fd_sc_hd__o21ai_2 _13274_ (.A1(_08177_),
    .A2(_08181_),
    .B1(net1770),
    .Y(_08182_));
 sky130_fd_sc_hd__o211a_4 _13275_ (.A1(net1770),
    .A2(\core.fetchProgramCounter[21] ),
    .B1(net1899),
    .C1(_08182_),
    .X(_08183_));
 sky130_fd_sc_hd__and2_2 _13276_ (.A(_07613_),
    .B(_07692_),
    .X(_08184_));
 sky130_fd_sc_hd__a21oi_2 _13277_ (.A1(_07701_),
    .A2(_08184_),
    .B1(_07707_),
    .Y(_08185_));
 sky130_fd_sc_hd__a211oi_1 _13278_ (.A1(_07611_),
    .A2(_07612_),
    .B1(_07683_),
    .C1(_07702_),
    .Y(_08186_));
 sky130_fd_sc_hd__or2_1 _13279_ (.A(_07709_),
    .B(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__nand2_1 _13280_ (.A(_07649_),
    .B(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__nand2_1 _13281_ (.A(_07647_),
    .B(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__a21oi_1 _13282_ (.A1(_07660_),
    .A2(_08189_),
    .B1(_07402_),
    .Y(_08190_));
 sky130_fd_sc_hd__o21a_1 _13283_ (.A1(_07660_),
    .A2(_08189_),
    .B1(_08190_),
    .X(_08191_));
 sky130_fd_sc_hd__and2_2 _13284_ (.A(\core.fetchProgramCounter[11] ),
    .B(_07899_),
    .X(_08192_));
 sky130_fd_sc_hd__a21oi_1 _13285_ (.A1(\core.fetchProgramCounter[12] ),
    .A2(_08192_),
    .B1(\core.fetchProgramCounter[13] ),
    .Y(_08193_));
 sky130_fd_sc_hd__and3_1 _13286_ (.A(\core.fetchProgramCounter[13] ),
    .B(\core.fetchProgramCounter[12] ),
    .C(_08192_),
    .X(_08194_));
 sky130_fd_sc_hd__nor2_1 _13287_ (.A(_08193_),
    .B(_08194_),
    .Y(_08195_));
 sky130_fd_sc_hd__a221o_1 _13288_ (.A1(\core.csr.trapReturnVector[13] ),
    .A2(net1180),
    .B1(net787),
    .B2(_08195_),
    .C1(net777),
    .X(_08196_));
 sky130_fd_sc_hd__a21oi_1 _13289_ (.A1(net2013),
    .A2(_08191_),
    .B1(_08196_),
    .Y(_08197_));
 sky130_fd_sc_hd__and3_1 _13290_ (.A(_07949_),
    .B(_07950_),
    .C(_07983_),
    .X(_08198_));
 sky130_fd_sc_hd__a21oi_1 _13291_ (.A1(_07949_),
    .A2(_07950_),
    .B1(_07983_),
    .Y(_08199_));
 sky130_fd_sc_hd__nand2_1 _13292_ (.A(\core.csr.traps.mtvec.csrReadData[13] ),
    .B(net1223),
    .Y(_08200_));
 sky130_fd_sc_hd__o311a_1 _13293_ (.A1(net1223),
    .A2(_08198_),
    .A3(_08199_),
    .B1(_08200_),
    .C1(net777),
    .X(_08201_));
 sky130_fd_sc_hd__o21ai_1 _13294_ (.A1(_08197_),
    .A2(_08201_),
    .B1(net1771),
    .Y(_08202_));
 sky130_fd_sc_hd__o211a_2 _13295_ (.A1(net1771),
    .A2(\core.fetchProgramCounter[13] ),
    .B1(net1915),
    .C1(_08202_),
    .X(_08203_));
 sky130_fd_sc_hd__nor2_1 _13296_ (.A(\core.fetchProgramCounter[19] ),
    .B(_07903_),
    .Y(_08204_));
 sky130_fd_sc_hd__a21oi_1 _13297_ (.A1(\core.csr.trapReturnVector[19] ),
    .A2(net1179),
    .B1(net774),
    .Y(_08205_));
 sky130_fd_sc_hd__o31a_1 _13298_ (.A1(_07439_),
    .A2(_07904_),
    .A3(_08204_),
    .B1(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__a21o_1 _13299_ (.A1(_07775_),
    .A2(_08155_),
    .B1(_07753_),
    .X(_08207_));
 sky130_fd_sc_hd__and3_1 _13300_ (.A(_07743_),
    .B(_07751_),
    .C(_08207_),
    .X(_08208_));
 sky130_fd_sc_hd__a21oi_2 _13301_ (.A1(_07751_),
    .A2(_08207_),
    .B1(_07743_),
    .Y(_08209_));
 sky130_fd_sc_hd__o31a_1 _13302_ (.A1(net797),
    .A2(_08208_),
    .A3(_08209_),
    .B1(_08206_),
    .X(_08210_));
 sky130_fd_sc_hd__and3_1 _13303_ (.A(_07939_),
    .B(_07940_),
    .C(_07990_),
    .X(_08211_));
 sky130_fd_sc_hd__a21oi_1 _13304_ (.A1(_07939_),
    .A2(_07940_),
    .B1(_07990_),
    .Y(_08212_));
 sky130_fd_sc_hd__nand2_1 _13305_ (.A(\core.csr.traps.mtvec.csrReadData[19] ),
    .B(_08005_),
    .Y(_08213_));
 sky130_fd_sc_hd__o311a_1 _13306_ (.A1(net1222),
    .A2(_08211_),
    .A3(_08212_),
    .B1(_08213_),
    .C1(net774),
    .X(_08214_));
 sky130_fd_sc_hd__o21ai_2 _13307_ (.A1(_08210_),
    .A2(_08214_),
    .B1(net1768),
    .Y(_08215_));
 sky130_fd_sc_hd__o211a_1 _13308_ (.A1(net1768),
    .A2(\core.fetchProgramCounter[19] ),
    .B1(net1909),
    .C1(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__or2_1 _13309_ (.A(_07649_),
    .B(_08187_),
    .X(_08217_));
 sky130_fd_sc_hd__a21o_1 _13310_ (.A1(_08188_),
    .A2(_08217_),
    .B1(_07402_),
    .X(_08218_));
 sky130_fd_sc_hd__or2_1 _13311_ (.A(\core.fetchProgramCounter[12] ),
    .B(_08192_),
    .X(_08219_));
 sky130_fd_sc_hd__a21oi_1 _13312_ (.A1(\core.fetchProgramCounter[12] ),
    .A2(_08192_),
    .B1(_07439_),
    .Y(_08220_));
 sky130_fd_sc_hd__a221o_1 _13313_ (.A1(\core.csr.trapReturnVector[12] ),
    .A2(net1180),
    .B1(_08219_),
    .B2(_08220_),
    .C1(net777),
    .X(_08221_));
 sky130_fd_sc_hd__a21oi_1 _13314_ (.A1(net2013),
    .A2(_08218_),
    .B1(_08221_),
    .Y(_08222_));
 sky130_fd_sc_hd__nand2b_1 _13315_ (.A_N(_07951_),
    .B(_07952_),
    .Y(_08223_));
 sky130_fd_sc_hd__or2_2 _13316_ (.A(_07982_),
    .B(_08223_),
    .X(_08224_));
 sky130_fd_sc_hd__a21oi_2 _13317_ (.A1(_07982_),
    .A2(_08223_),
    .B1(net1223),
    .Y(_08225_));
 sky130_fd_sc_hd__a221oi_4 _13318_ (.A1(\core.csr.traps.mtvec.csrReadData[12] ),
    .A2(net1223),
    .B1(_08224_),
    .B2(_08225_),
    .C1(net767),
    .Y(_08226_));
 sky130_fd_sc_hd__o21ai_1 _13319_ (.A1(_08222_),
    .A2(_08226_),
    .B1(net1771),
    .Y(_08227_));
 sky130_fd_sc_hd__o211a_2 _13320_ (.A1(net1771),
    .A2(\core.fetchProgramCounter[12] ),
    .B1(net1915),
    .C1(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__nand3_1 _13321_ (.A(_07753_),
    .B(_07775_),
    .C(_08155_),
    .Y(_08229_));
 sky130_fd_sc_hd__a31o_1 _13322_ (.A1(\core.fetchProgramCounter[9] ),
    .A2(_07898_),
    .A3(_07902_),
    .B1(\core.fetchProgramCounter[18] ),
    .X(_08230_));
 sky130_fd_sc_hd__and3b_1 _13323_ (.A_N(_07903_),
    .B(_08230_),
    .C(net788),
    .X(_08231_));
 sky130_fd_sc_hd__a211o_1 _13324_ (.A1(\core.csr.trapReturnVector[18] ),
    .A2(net1179),
    .B1(_08231_),
    .C1(net774),
    .X(_08232_));
 sky130_fd_sc_hd__a31o_1 _13325_ (.A1(net793),
    .A2(_08207_),
    .A3(_08229_),
    .B1(_08232_),
    .X(_08233_));
 sky130_fd_sc_hd__nand2b_1 _13326_ (.A_N(_07941_),
    .B(_07942_),
    .Y(_08234_));
 sky130_fd_sc_hd__xnor2_1 _13327_ (.A(_07989_),
    .B(_08234_),
    .Y(_08235_));
 sky130_fd_sc_hd__nor2_1 _13328_ (.A(net1222),
    .B(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__a211o_1 _13329_ (.A1(\core.csr.traps.mtvec.csrReadData[18] ),
    .A2(net1222),
    .B1(_08236_),
    .C1(net768),
    .X(_08237_));
 sky130_fd_sc_hd__a21o_1 _13330_ (.A1(_08233_),
    .A2(_08237_),
    .B1(net1761),
    .X(_08238_));
 sky130_fd_sc_hd__o211a_1 _13331_ (.A1(net1769),
    .A2(\core.fetchProgramCounter[18] ),
    .B1(net1909),
    .C1(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__and3_1 _13332_ (.A(_07765_),
    .B(_07771_),
    .C(_08154_),
    .X(_08240_));
 sky130_fd_sc_hd__a21oi_1 _13333_ (.A1(_07771_),
    .A2(_08154_),
    .B1(_07765_),
    .Y(_08241_));
 sky130_fd_sc_hd__or3_1 _13334_ (.A(net797),
    .B(_08240_),
    .C(_08241_),
    .X(_08242_));
 sky130_fd_sc_hd__and4_2 _13335_ (.A(\core.fetchProgramCounter[14] ),
    .B(\core.fetchProgramCounter[13] ),
    .C(\core.fetchProgramCounter[12] ),
    .D(_08192_),
    .X(_08243_));
 sky130_fd_sc_hd__and3_1 _13336_ (.A(\core.fetchProgramCounter[16] ),
    .B(\core.fetchProgramCounter[15] ),
    .C(_08243_),
    .X(_08244_));
 sky130_fd_sc_hd__xor2_1 _13337_ (.A(\core.fetchProgramCounter[17] ),
    .B(_08244_),
    .X(_08245_));
 sky130_fd_sc_hd__a221oi_2 _13338_ (.A1(\core.csr.trapReturnVector[17] ),
    .A2(net1179),
    .B1(net788),
    .B2(_08245_),
    .C1(net775),
    .Y(_08246_));
 sky130_fd_sc_hd__xor2_1 _13339_ (.A(\core.csr.traps.mtvec.csrReadData[17] ),
    .B(\core.csr.traps.mcause.csrReadData[15] ),
    .X(_08247_));
 sky130_fd_sc_hd__nand2_1 _13340_ (.A(_07987_),
    .B(_08247_),
    .Y(_08248_));
 sky130_fd_sc_hd__o21ba_1 _13341_ (.A1(_07987_),
    .A2(_08247_),
    .B1_N(net1222),
    .X(_08249_));
 sky130_fd_sc_hd__a22o_1 _13342_ (.A1(\core.csr.traps.mtvec.csrReadData[17] ),
    .A2(net1222),
    .B1(_08248_),
    .B2(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__o21ai_1 _13343_ (.A1(net768),
    .A2(_08250_),
    .B1(net1769),
    .Y(_08251_));
 sky130_fd_sc_hd__a21oi_1 _13344_ (.A1(_08242_),
    .A2(_08246_),
    .B1(_08251_),
    .Y(_08252_));
 sky130_fd_sc_hd__a21o_1 _13345_ (.A1(net1761),
    .A2(\core.fetchProgramCounter[17] ),
    .B1(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__nand3_1 _13346_ (.A(_07704_),
    .B(_07710_),
    .C(_07772_),
    .Y(_08254_));
 sky130_fd_sc_hd__nand2_1 _13347_ (.A(_08154_),
    .B(_08254_),
    .Y(_08255_));
 sky130_fd_sc_hd__a21o_1 _13348_ (.A1(_07403_),
    .A2(_08255_),
    .B1(net797),
    .X(_08256_));
 sky130_fd_sc_hd__a21o_1 _13349_ (.A1(\core.fetchProgramCounter[15] ),
    .A2(_08243_),
    .B1(\core.fetchProgramCounter[16] ),
    .X(_08257_));
 sky130_fd_sc_hd__or4b_1 _13350_ (.A(net793),
    .B(net1179),
    .C(_08244_),
    .D_N(_08257_),
    .X(_08258_));
 sky130_fd_sc_hd__a21oi_1 _13351_ (.A1(\core.csr.trapReturnVector[16] ),
    .A2(net1179),
    .B1(net775),
    .Y(_08259_));
 sky130_fd_sc_hd__and3_1 _13352_ (.A(_08256_),
    .B(_08258_),
    .C(_08259_),
    .X(_08260_));
 sky130_fd_sc_hd__nand2b_1 _13353_ (.A_N(_07943_),
    .B(_07944_),
    .Y(_08261_));
 sky130_fd_sc_hd__xnor2_1 _13354_ (.A(_07986_),
    .B(_08261_),
    .Y(_08262_));
 sky130_fd_sc_hd__nand2_1 _13355_ (.A(\core.csr.traps.mtvec.csrReadData[16] ),
    .B(net1222),
    .Y(_08263_));
 sky130_fd_sc_hd__o211a_1 _13356_ (.A1(net1222),
    .A2(_08262_),
    .B1(_08263_),
    .C1(net775),
    .X(_08264_));
 sky130_fd_sc_hd__o21a_1 _13357_ (.A1(_08260_),
    .A2(_08264_),
    .B1(net1769),
    .X(_08265_));
 sky130_fd_sc_hd__a211o_1 _13358_ (.A1(net1761),
    .A2(_04410_),
    .B1(net1970),
    .C1(_08265_),
    .X(_08266_));
 sky130_fd_sc_hd__inv_2 _13359_ (.A(_08266_),
    .Y(_08267_));
 sky130_fd_sc_hd__a21bo_1 _13360_ (.A1(net1909),
    .A2(_08253_),
    .B1_N(_08266_),
    .X(_08268_));
 sky130_fd_sc_hd__or4_1 _13361_ (.A(_08216_),
    .B(_08228_),
    .C(_08239_),
    .D(_08268_),
    .X(_08269_));
 sky130_fd_sc_hd__and3_1 _13362_ (.A(_07727_),
    .B(_07778_),
    .C(_08156_),
    .X(_08270_));
 sky130_fd_sc_hd__nand2_1 _13363_ (.A(\core.csr.trapReturnVector[20] ),
    .B(net1177),
    .Y(_08271_));
 sky130_fd_sc_hd__o211a_1 _13364_ (.A1(_08157_),
    .A2(_08270_),
    .B1(net793),
    .C1(_07403_),
    .X(_08272_));
 sky130_fd_sc_hd__xnor2_1 _13365_ (.A(\core.fetchProgramCounter[20] ),
    .B(_07904_),
    .Y(_08273_));
 sky130_fd_sc_hd__a211o_1 _13366_ (.A1(net797),
    .A2(_08273_),
    .B1(_08272_),
    .C1(net1178),
    .X(_08274_));
 sky130_fd_sc_hd__nand2b_1 _13367_ (.A_N(_07937_),
    .B(_07938_),
    .Y(_08275_));
 sky130_fd_sc_hd__nor2_1 _13368_ (.A(_07991_),
    .B(_08275_),
    .Y(_08276_));
 sky130_fd_sc_hd__a21o_1 _13369_ (.A1(_07991_),
    .A2(_08275_),
    .B1(net1221),
    .X(_08277_));
 sky130_fd_sc_hd__nand2_1 _13370_ (.A(\core.csr.traps.mtvec.csrReadData[20] ),
    .B(net1221),
    .Y(_08278_));
 sky130_fd_sc_hd__o211a_1 _13371_ (.A1(_08276_),
    .A2(_08277_),
    .B1(_08278_),
    .C1(net774),
    .X(_08279_));
 sky130_fd_sc_hd__a31o_1 _13372_ (.A1(net766),
    .A2(_08271_),
    .A3(_08274_),
    .B1(_08279_),
    .X(_08280_));
 sky130_fd_sc_hd__nand2_1 _13373_ (.A(net1768),
    .B(_08280_),
    .Y(_08281_));
 sky130_fd_sc_hd__o211a_2 _13374_ (.A1(net1768),
    .A2(\core.fetchProgramCounter[20] ),
    .B1(net1900),
    .C1(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__a31o_1 _13375_ (.A1(_07647_),
    .A2(_07659_),
    .A3(_08188_),
    .B1(_07658_),
    .X(_08283_));
 sky130_fd_sc_hd__and2_1 _13376_ (.A(_07637_),
    .B(_08283_),
    .X(_08284_));
 sky130_fd_sc_hd__nor2_2 _13377_ (.A(_07637_),
    .B(_08283_),
    .Y(_08285_));
 sky130_fd_sc_hd__nor2_1 _13378_ (.A(\core.fetchProgramCounter[14] ),
    .B(_08194_),
    .Y(_08286_));
 sky130_fd_sc_hd__a21oi_1 _13379_ (.A1(\core.csr.trapReturnVector[14] ),
    .A2(net1180),
    .B1(net777),
    .Y(_08287_));
 sky130_fd_sc_hd__o31a_1 _13380_ (.A1(_07439_),
    .A2(_08243_),
    .A3(_08286_),
    .B1(_08287_),
    .X(_08288_));
 sky130_fd_sc_hd__o31a_1 _13381_ (.A1(net798),
    .A2(_08284_),
    .A3(_08285_),
    .B1(_08288_),
    .X(_08289_));
 sky130_fd_sc_hd__nand2b_1 _13382_ (.A_N(_07947_),
    .B(_07948_),
    .Y(_08290_));
 sky130_fd_sc_hd__or2_2 _13383_ (.A(_07984_),
    .B(_08290_),
    .X(_08291_));
 sky130_fd_sc_hd__a21oi_2 _13384_ (.A1(_07984_),
    .A2(_08290_),
    .B1(net1223),
    .Y(_08292_));
 sky130_fd_sc_hd__a221oi_4 _13385_ (.A1(\core.csr.traps.mtvec.csrReadData[14] ),
    .A2(net1223),
    .B1(_08291_),
    .B2(_08292_),
    .C1(net767),
    .Y(_08293_));
 sky130_fd_sc_hd__o21ai_1 _13386_ (.A1(_08289_),
    .A2(_08293_),
    .B1(net1771),
    .Y(_08294_));
 sky130_fd_sc_hd__o211a_1 _13387_ (.A1(net1771),
    .A2(\core.fetchProgramCounter[14] ),
    .B1(net1910),
    .C1(_08294_),
    .X(_08295_));
 sky130_fd_sc_hd__or4_1 _13388_ (.A(_08203_),
    .B(_08269_),
    .C(_08282_),
    .D(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__or3_2 _13389_ (.A(_07721_),
    .B(_07779_),
    .C(_08159_),
    .X(_08297_));
 sky130_fd_sc_hd__or2_1 _13390_ (.A(\core.fetchProgramCounter[22] ),
    .B(_07905_),
    .X(_08298_));
 sky130_fd_sc_hd__a21o_1 _13391_ (.A1(\core.csr.trapReturnVector[22] ),
    .A2(net1177),
    .B1(net770),
    .X(_08299_));
 sky130_fd_sc_hd__a31o_1 _13392_ (.A1(net788),
    .A2(_07906_),
    .A3(_08298_),
    .B1(_08299_),
    .X(_08300_));
 sky130_fd_sc_hd__a31oi_4 _13393_ (.A1(net792),
    .A2(_08160_),
    .A3(_08297_),
    .B1(_08300_),
    .Y(_08301_));
 sky130_fd_sc_hd__nand2b_1 _13394_ (.A_N(_07933_),
    .B(_07934_),
    .Y(_08302_));
 sky130_fd_sc_hd__nor2_1 _13395_ (.A(_07993_),
    .B(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__a21o_1 _13396_ (.A1(_07993_),
    .A2(_08302_),
    .B1(net1219),
    .X(_08304_));
 sky130_fd_sc_hd__nand2_1 _13397_ (.A(\core.csr.traps.mtvec.csrReadData[22] ),
    .B(net1219),
    .Y(_08305_));
 sky130_fd_sc_hd__o211a_2 _13398_ (.A1(_08303_),
    .A2(_08304_),
    .B1(_08305_),
    .C1(net769),
    .X(_08306_));
 sky130_fd_sc_hd__o21ai_2 _13399_ (.A1(_08301_),
    .A2(_08306_),
    .B1(net1766),
    .Y(_08307_));
 sky130_fd_sc_hd__o211a_4 _13400_ (.A1(net1766),
    .A2(\core.fetchProgramCounter[22] ),
    .B1(net1888),
    .C1(_08307_),
    .X(_08308_));
 sky130_fd_sc_hd__o21ai_1 _13401_ (.A1(_07635_),
    .A2(_08285_),
    .B1(_07627_),
    .Y(_08309_));
 sky130_fd_sc_hd__o31a_1 _13402_ (.A1(_07627_),
    .A2(_07635_),
    .A3(_08285_),
    .B1(net2013),
    .X(_08310_));
 sky130_fd_sc_hd__xor2_1 _13403_ (.A(\core.fetchProgramCounter[15] ),
    .B(_08243_),
    .X(_08311_));
 sky130_fd_sc_hd__a221o_1 _13404_ (.A1(\core.csr.trapReturnVector[15] ),
    .A2(net1179),
    .B1(net788),
    .B2(_08311_),
    .C1(net775),
    .X(_08312_));
 sky130_fd_sc_hd__a21o_1 _13405_ (.A1(_08309_),
    .A2(_08310_),
    .B1(_08312_),
    .X(_08313_));
 sky130_fd_sc_hd__a21oi_1 _13406_ (.A1(_07945_),
    .A2(_07946_),
    .B1(_07985_),
    .Y(_08314_));
 sky130_fd_sc_hd__a311oi_2 _13407_ (.A1(_07945_),
    .A2(_07946_),
    .A3(_07985_),
    .B1(net1222),
    .C1(_08314_),
    .Y(_08315_));
 sky130_fd_sc_hd__a211o_1 _13408_ (.A1(\core.csr.traps.mtvec.csrReadData[15] ),
    .A2(net1222),
    .B1(_08315_),
    .C1(net766),
    .X(_08316_));
 sky130_fd_sc_hd__a21o_1 _13409_ (.A1(_08313_),
    .A2(_08316_),
    .B1(net1761),
    .X(_08317_));
 sky130_fd_sc_hd__o211a_1 _13410_ (.A1(net1769),
    .A2(\core.fetchProgramCounter[15] ),
    .B1(net1910),
    .C1(_08317_),
    .X(_08318_));
 sky130_fd_sc_hd__or2_1 _13411_ (.A(_08308_),
    .B(_08318_),
    .X(_08319_));
 sky130_fd_sc_hd__or4_4 _13412_ (.A(_08171_),
    .B(_08183_),
    .C(_08296_),
    .D(_08319_),
    .X(_08320_));
 sky130_fd_sc_hd__xor2_4 _13413_ (.A(_04697_),
    .B(_08081_),
    .X(_08321_));
 sky130_fd_sc_hd__xnor2_4 _13414_ (.A(_04777_),
    .B(_08080_),
    .Y(_08322_));
 sky130_fd_sc_hd__xnor2_4 _13415_ (.A(_04854_),
    .B(_08079_),
    .Y(_08323_));
 sky130_fd_sc_hd__xnor2_4 _13416_ (.A(_06656_),
    .B(_08078_),
    .Y(_08324_));
 sky130_fd_sc_hd__clkinv_2 _13417_ (.A(_08324_),
    .Y(_08325_));
 sky130_fd_sc_hd__xor2_4 _13418_ (.A(_06565_),
    .B(_08076_),
    .X(_08326_));
 sky130_fd_sc_hd__xor2_4 _13419_ (.A(_06643_),
    .B(_08074_),
    .X(_08327_));
 sky130_fd_sc_hd__xnor2_4 _13420_ (.A(_06410_),
    .B(_08073_),
    .Y(_08328_));
 sky130_fd_sc_hd__xnor2_4 _13421_ (.A(_06488_),
    .B(_08071_),
    .Y(_08329_));
 sky130_fd_sc_hd__xnor2_4 _13422_ (.A(_05191_),
    .B(_08070_),
    .Y(_08330_));
 sky130_fd_sc_hd__xnor2_4 _13423_ (.A(_05279_),
    .B(_08069_),
    .Y(_08331_));
 sky130_fd_sc_hd__xnor2_4 _13424_ (.A(_05111_),
    .B(_08068_),
    .Y(_08332_));
 sky130_fd_sc_hd__xnor2_4 _13425_ (.A(_05026_),
    .B(_08067_),
    .Y(_08333_));
 sky130_fd_sc_hd__or4_1 _13426_ (.A(_08330_),
    .B(_08331_),
    .C(_08332_),
    .D(_08333_),
    .X(_08334_));
 sky130_fd_sc_hd__or4_1 _13427_ (.A(_08327_),
    .B(_08328_),
    .C(_08329_),
    .D(_08334_),
    .X(_08335_));
 sky130_fd_sc_hd__or4_1 _13428_ (.A(_08323_),
    .B(_08325_),
    .C(_08326_),
    .D(_08335_),
    .X(_08336_));
 sky130_fd_sc_hd__or3b_2 _13429_ (.A(_08321_),
    .B(_08336_),
    .C_N(_08322_),
    .X(_08337_));
 sky130_fd_sc_hd__inv_2 _13430_ (.A(_08337_),
    .Y(_08338_));
 sky130_fd_sc_hd__xnor2_4 _13431_ (.A(_06949_),
    .B(_08085_),
    .Y(_08339_));
 sky130_fd_sc_hd__xor2_4 _13432_ (.A(_07024_),
    .B(_08084_),
    .X(_08340_));
 sky130_fd_sc_hd__xnor2_4 _13433_ (.A(_06870_),
    .B(_08083_),
    .Y(_08341_));
 sky130_fd_sc_hd__xnor2_4 _13434_ (.A(_06791_),
    .B(_08082_),
    .Y(_08342_));
 sky130_fd_sc_hd__or4_1 _13435_ (.A(_08097_),
    .B(_08340_),
    .C(_08341_),
    .D(_08342_),
    .X(_08343_));
 sky130_fd_sc_hd__or4b_1 _13436_ (.A(net765),
    .B(_08343_),
    .C(_08339_),
    .D_N(_08093_),
    .X(_08344_));
 sky130_fd_sc_hd__or2_4 _13437_ (.A(_08098_),
    .B(_08344_),
    .X(_08345_));
 sky130_fd_sc_hd__a21oi_4 _13438_ (.A1(_08025_),
    .A2(_08151_),
    .B1(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__or3_1 _13439_ (.A(_08339_),
    .B(_08340_),
    .C(_08341_),
    .X(_08347_));
 sky130_fd_sc_hd__or3b_1 _13440_ (.A(_08347_),
    .B(net765),
    .C_N(_08093_),
    .X(_08348_));
 sky130_fd_sc_hd__a2111o_1 _13441_ (.A1(net807),
    .A2(_08348_),
    .B1(_08342_),
    .C1(_08098_),
    .D1(_08097_),
    .X(_08349_));
 sky130_fd_sc_hd__a2bb2o_4 _13442_ (.A1_N(_08153_),
    .A2_N(_08320_),
    .B1(_08338_),
    .B2(net724),
    .X(_08350_));
 sky130_fd_sc_hd__nand2_8 _13443_ (.A(_04467_),
    .B(_07481_),
    .Y(_08351_));
 sky130_fd_sc_hd__inv_4 _13444_ (.A(_08351_),
    .Y(_08352_));
 sky130_fd_sc_hd__a21oi_4 _13445_ (.A1(net2010),
    .A2(_08352_),
    .B1(\localMemoryInterface.coreReadReady ),
    .Y(_08353_));
 sky130_fd_sc_hd__nand2_8 _13446_ (.A(_08350_),
    .B(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__o21a_1 _13447_ (.A1(_07682_),
    .A2(_08185_),
    .B1(_07680_),
    .X(_08355_));
 sky130_fd_sc_hd__xnor2_1 _13448_ (.A(_07673_),
    .B(_08355_),
    .Y(_08356_));
 sky130_fd_sc_hd__nor2_1 _13449_ (.A(\core.fetchProgramCounter[11] ),
    .B(_07899_),
    .Y(_08357_));
 sky130_fd_sc_hd__nor2_1 _13450_ (.A(_08192_),
    .B(_08357_),
    .Y(_08358_));
 sky130_fd_sc_hd__a221o_1 _13451_ (.A1(\core.csr.trapReturnVector[11] ),
    .A2(net1180),
    .B1(net787),
    .B2(_08358_),
    .C1(net777),
    .X(_08359_));
 sky130_fd_sc_hd__a21oi_1 _13452_ (.A1(net2013),
    .A2(_08356_),
    .B1(_08359_),
    .Y(_08360_));
 sky130_fd_sc_hd__and3_1 _13453_ (.A(_07953_),
    .B(_07954_),
    .C(_07981_),
    .X(_08361_));
 sky130_fd_sc_hd__a21oi_1 _13454_ (.A1(_07953_),
    .A2(_07954_),
    .B1(_07981_),
    .Y(_08362_));
 sky130_fd_sc_hd__nand2_1 _13455_ (.A(\core.csr.traps.mtvec.csrReadData[11] ),
    .B(net1223),
    .Y(_08363_));
 sky130_fd_sc_hd__o311a_2 _13456_ (.A1(net1223),
    .A2(_08361_),
    .A3(_08362_),
    .B1(_08363_),
    .C1(net778),
    .X(_08364_));
 sky130_fd_sc_hd__o21a_1 _13457_ (.A1(_08360_),
    .A2(_08364_),
    .B1(net1771),
    .X(_08365_));
 sky130_fd_sc_hd__a211oi_4 _13458_ (.A1(net1765),
    .A2(_04411_),
    .B1(net1970),
    .C1(_08365_),
    .Y(_08366_));
 sky130_fd_sc_hd__xnor2_4 _13459_ (.A(_05368_),
    .B(_08066_),
    .Y(_08367_));
 sky130_fd_sc_hd__a32o_4 _13460_ (.A1(net806),
    .A2(net724),
    .A3(_08367_),
    .B1(_08366_),
    .B2(_08152_),
    .X(_08368_));
 sky130_fd_sc_hd__nand2b_1 _13461_ (.A_N(_08354_),
    .B(_08368_),
    .Y(net375));
 sky130_fd_sc_hd__or2_1 _13462_ (.A(_08354_),
    .B(_08368_),
    .X(net374));
 sky130_fd_sc_hd__and3_4 _13463_ (.A(net724),
    .B(_08350_),
    .C(_08352_),
    .X(_08369_));
 sky130_fd_sc_hd__or4_1 _13464_ (.A(\wbSRAMInterface.currentAddress[16] ),
    .B(\wbSRAMInterface.currentAddress[14] ),
    .C(\wbSRAMInterface.currentAddress[15] ),
    .D(\wbSRAMInterface.currentAddress[13] ),
    .X(_08370_));
 sky130_fd_sc_hd__o31a_1 _13465_ (.A1(\wbSRAMInterface.currentAddress[12] ),
    .A2(_07860_),
    .A3(_08370_),
    .B1(_07837_),
    .X(_08371_));
 sky130_fd_sc_hd__or2_2 _13466_ (.A(net205),
    .B(_07839_),
    .X(_08372_));
 sky130_fd_sc_hd__or4_4 _13467_ (.A(\wbSRAMInterface.currentAddress[20] ),
    .B(\wbSRAMInterface.currentAddress[21] ),
    .C(\wbSRAMInterface.currentAddress[22] ),
    .D(\wbSRAMInterface.currentAddress[23] ),
    .X(_08373_));
 sky130_fd_sc_hd__nor3_4 _13468_ (.A(_08371_),
    .B(net1305),
    .C(_08373_),
    .Y(_08374_));
 sky130_fd_sc_hd__a21oi_4 _13469_ (.A1(_07865_),
    .A2(net1254),
    .B1(net712),
    .Y(net483));
 sky130_fd_sc_hd__nand2_2 _13470_ (.A(_07866_),
    .B(net1254),
    .Y(_08375_));
 sky130_fd_sc_hd__or2_4 _13471_ (.A(\localMemoryInterface.wbReadReady ),
    .B(_08375_),
    .X(_08376_));
 sky130_fd_sc_hd__inv_2 _13472_ (.A(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__and2b_2 _13473_ (.A_N(net712),
    .B(net1254),
    .X(_08378_));
 sky130_fd_sc_hd__a22o_4 _13474_ (.A1(_08368_),
    .A2(net712),
    .B1(net702),
    .B2(\wbSRAMInterface.currentAddress[11] ),
    .X(_08379_));
 sky130_fd_sc_hd__a21bo_1 _13475_ (.A1(net483),
    .A2(_08376_),
    .B1_N(_08379_),
    .X(net373));
 sky130_fd_sc_hd__a21o_1 _13476_ (.A1(net483),
    .A2(_08376_),
    .B1(_08379_),
    .X(net372));
 sky130_fd_sc_hd__and2_1 _13477_ (.A(\coreWBInterface.stb ),
    .B(_08101_),
    .X(net370));
 sky130_fd_sc_hd__and2_2 _13478_ (.A(_07443_),
    .B(net729),
    .X(net305));
 sky130_fd_sc_hd__and2_4 _13479_ (.A(_07437_),
    .B(net727),
    .X(net316));
 sky130_fd_sc_hd__nor2_2 _13480_ (.A(net728),
    .B(_08100_),
    .Y(_08380_));
 sky130_fd_sc_hd__or2_4 _13481_ (.A(net727),
    .B(_08100_),
    .X(_08381_));
 sky130_fd_sc_hd__xor2_4 _13482_ (.A(_06053_),
    .B(_08054_),
    .X(_08382_));
 sky130_fd_sc_hd__a21oi_1 _13483_ (.A1(_07584_),
    .A2(_07586_),
    .B1(_07585_),
    .Y(_08383_));
 sky130_fd_sc_hd__o21ai_1 _13484_ (.A1(_07587_),
    .A2(_08383_),
    .B1(_07403_),
    .Y(_08384_));
 sky130_fd_sc_hd__o21ai_1 _13485_ (.A1(\core.fetchProgramCounter[2] ),
    .A2(_07891_),
    .B1(net787),
    .Y(_08385_));
 sky130_fd_sc_hd__a21oi_2 _13486_ (.A1(\core.csr.trapReturnVector[2] ),
    .A2(net1180),
    .B1(net781),
    .Y(_08386_));
 sky130_fd_sc_hd__o21ai_1 _13487_ (.A1(_07894_),
    .A2(_08385_),
    .B1(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__a21o_1 _13488_ (.A1(net796),
    .A2(_08384_),
    .B1(_08387_),
    .X(_08388_));
 sky130_fd_sc_hd__o21a_1 _13489_ (.A1(_04395_),
    .A2(net1224),
    .B1(\core.csr.traps.mtvec.csrReadData[2] ),
    .X(_08389_));
 sky130_fd_sc_hd__o31ai_1 _13490_ (.A1(\core.csr.traps.mtvec.csrReadData[2] ),
    .A2(_04395_),
    .A3(net1224),
    .B1(net783),
    .Y(_08390_));
 sky130_fd_sc_hd__o211a_2 _13491_ (.A1(_08389_),
    .A2(_08390_),
    .B1(net1774),
    .C1(_08388_),
    .X(_08391_));
 sky130_fd_sc_hd__a21oi_4 _13492_ (.A1(net1763),
    .A2(\core.fetchProgramCounter[2] ),
    .B1(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__nor2_2 _13493_ (.A(net1970),
    .B(_08392_),
    .Y(_08393_));
 sky130_fd_sc_hd__a32o_4 _13494_ (.A1(net806),
    .A2(net723),
    .A3(_08382_),
    .B1(_08393_),
    .B2(net728),
    .X(net325));
 sky130_fd_sc_hd__xnor2_4 _13495_ (.A(_05968_),
    .B(_08056_),
    .Y(_08394_));
 sky130_fd_sc_hd__inv_2 _13496_ (.A(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__nor2_2 _13497_ (.A(_08096_),
    .B(_08394_),
    .Y(_08396_));
 sky130_fd_sc_hd__nor2_1 _13498_ (.A(\core.fetchProgramCounter[3] ),
    .B(_07894_),
    .Y(_08397_));
 sky130_fd_sc_hd__nor2_1 _13499_ (.A(_07895_),
    .B(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__a221o_1 _13500_ (.A1(\core.csr.trapReturnVector[3] ),
    .A2(net1180),
    .B1(_07438_),
    .B2(_08398_),
    .C1(net782),
    .X(_08399_));
 sky130_fd_sc_hd__or3_1 _13501_ (.A(_07573_),
    .B(_07574_),
    .C(_07588_),
    .X(_08400_));
 sky130_fd_sc_hd__o21ai_1 _13502_ (.A1(_07573_),
    .A2(_07574_),
    .B1(_07588_),
    .Y(_08401_));
 sky130_fd_sc_hd__a31o_1 _13503_ (.A1(net795),
    .A2(_08400_),
    .A3(_08401_),
    .B1(_08399_),
    .X(_08402_));
 sky130_fd_sc_hd__a22o_1 _13504_ (.A1(\core.csr.traps.mtvec.csrReadData[2] ),
    .A2(\core.csr.traps.mcause.csrReadData[0] ),
    .B1(_07970_),
    .B2(_07971_),
    .X(_08403_));
 sky130_fd_sc_hd__nor2_1 _13505_ (.A(_07972_),
    .B(net1225),
    .Y(_08404_));
 sky130_fd_sc_hd__a221o_1 _13506_ (.A1(\core.csr.traps.mtvec.csrReadData[3] ),
    .A2(net1225),
    .B1(_08403_),
    .B2(_08404_),
    .C1(net767),
    .X(_08405_));
 sky130_fd_sc_hd__and3_2 _13507_ (.A(net1774),
    .B(_08402_),
    .C(_08405_),
    .X(_08406_));
 sky130_fd_sc_hd__a21oi_4 _13508_ (.A1(net1763),
    .A2(\core.fetchProgramCounter[3] ),
    .B1(_08406_),
    .Y(_08407_));
 sky130_fd_sc_hd__nor2_1 _13509_ (.A(net1970),
    .B(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__a22o_4 _13510_ (.A1(net720),
    .A2(_08396_),
    .B1(_08408_),
    .B2(net728),
    .X(net326));
 sky130_fd_sc_hd__nor2_1 _13511_ (.A(_07590_),
    .B(_07599_),
    .Y(_08409_));
 sky130_fd_sc_hd__or2_1 _13512_ (.A(_07600_),
    .B(_08409_),
    .X(_08410_));
 sky130_fd_sc_hd__a21oi_2 _13513_ (.A1(_07403_),
    .A2(_08410_),
    .B1(net798),
    .Y(_08411_));
 sky130_fd_sc_hd__a21oi_1 _13514_ (.A1(\core.fetchProgramCounter[4] ),
    .A2(_07895_),
    .B1(_07439_),
    .Y(_08412_));
 sky130_fd_sc_hd__o21a_1 _13515_ (.A1(\core.fetchProgramCounter[4] ),
    .A2(_07895_),
    .B1(_08412_),
    .X(_08413_));
 sky130_fd_sc_hd__a2111o_1 _13516_ (.A1(\core.csr.trapReturnVector[4] ),
    .A2(net1181),
    .B1(_08411_),
    .C1(_08413_),
    .D1(net782),
    .X(_08414_));
 sky130_fd_sc_hd__nand2b_1 _13517_ (.A_N(_07968_),
    .B(_07969_),
    .Y(_08415_));
 sky130_fd_sc_hd__xor2_1 _13518_ (.A(_07973_),
    .B(_08415_),
    .X(_08416_));
 sky130_fd_sc_hd__mux2_1 _13519_ (.A0(_08416_),
    .A1(\core.csr.traps.mtvec.csrReadData[4] ),
    .S(net1225),
    .X(_08417_));
 sky130_fd_sc_hd__o211a_2 _13520_ (.A1(net767),
    .A2(_08417_),
    .B1(_08414_),
    .C1(net1775),
    .X(_08418_));
 sky130_fd_sc_hd__a21oi_4 _13521_ (.A1(net1762),
    .A2(\core.fetchProgramCounter[4] ),
    .B1(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__nor2_2 _13522_ (.A(net1970),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__xor2_4 _13523_ (.A(_05883_),
    .B(_08057_),
    .X(_08421_));
 sky130_fd_sc_hd__inv_2 _13524_ (.A(_08421_),
    .Y(_08422_));
 sky130_fd_sc_hd__a22o_4 _13525_ (.A1(net728),
    .A2(_08420_),
    .B1(_08422_),
    .B2(net720),
    .X(net327));
 sky130_fd_sc_hd__or3_1 _13526_ (.A(_07597_),
    .B(_07600_),
    .C(_07603_),
    .X(_08423_));
 sky130_fd_sc_hd__o21ai_1 _13527_ (.A1(_07597_),
    .A2(_07600_),
    .B1(_07603_),
    .Y(_08424_));
 sky130_fd_sc_hd__a31o_1 _13528_ (.A1(\core.fetchProgramCounter[4] ),
    .A2(\core.fetchProgramCounter[3] ),
    .A3(_07894_),
    .B1(\core.fetchProgramCounter[5] ),
    .X(_08425_));
 sky130_fd_sc_hd__and2b_1 _13529_ (.A_N(_07896_),
    .B(_08425_),
    .X(_08426_));
 sky130_fd_sc_hd__a221o_1 _13530_ (.A1(\core.csr.trapReturnVector[5] ),
    .A2(net1181),
    .B1(net787),
    .B2(_08426_),
    .C1(net782),
    .X(_08427_));
 sky130_fd_sc_hd__a31o_1 _13531_ (.A1(net795),
    .A2(_08423_),
    .A3(_08424_),
    .B1(_08427_),
    .X(_08428_));
 sky130_fd_sc_hd__a21oi_1 _13532_ (.A1(_07966_),
    .A2(_07967_),
    .B1(_07974_),
    .Y(_08429_));
 sky130_fd_sc_hd__a31o_1 _13533_ (.A1(_07966_),
    .A2(_07967_),
    .A3(_07974_),
    .B1(net1224),
    .X(_08430_));
 sky130_fd_sc_hd__a2bb2o_1 _13534_ (.A1_N(_08429_),
    .A2_N(_08430_),
    .B1(\core.csr.traps.mtvec.csrReadData[5] ),
    .B2(net1224),
    .X(_08431_));
 sky130_fd_sc_hd__o211a_2 _13535_ (.A1(net767),
    .A2(_08431_),
    .B1(_08428_),
    .C1(net1774),
    .X(_08432_));
 sky130_fd_sc_hd__a21oi_4 _13536_ (.A1(net1762),
    .A2(\core.fetchProgramCounter[5] ),
    .B1(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__nor2_2 _13537_ (.A(net1970),
    .B(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__xnor2_4 _13538_ (.A(_05798_),
    .B(_08058_),
    .Y(_08435_));
 sky130_fd_sc_hd__nor2_2 _13539_ (.A(_08096_),
    .B(_08435_),
    .Y(_08436_));
 sky130_fd_sc_hd__a22o_4 _13540_ (.A1(net728),
    .A2(_08434_),
    .B1(_08436_),
    .B2(net723),
    .X(net328));
 sky130_fd_sc_hd__xnor2_4 _13541_ (.A(_05713_),
    .B(_08059_),
    .Y(_08437_));
 sky130_fd_sc_hd__and2_1 _13542_ (.A(net806),
    .B(_08437_),
    .X(_08438_));
 sky130_fd_sc_hd__or2_1 _13543_ (.A(_07606_),
    .B(_07609_),
    .X(_08439_));
 sky130_fd_sc_hd__nand2_1 _13544_ (.A(_07606_),
    .B(_07609_),
    .Y(_08440_));
 sky130_fd_sc_hd__or2_1 _13545_ (.A(\core.fetchProgramCounter[6] ),
    .B(_07896_),
    .X(_08441_));
 sky130_fd_sc_hd__a21o_1 _13546_ (.A1(\core.csr.trapReturnVector[6] ),
    .A2(net1181),
    .B1(net780),
    .X(_08442_));
 sky130_fd_sc_hd__a31o_1 _13547_ (.A1(net787),
    .A2(_07897_),
    .A3(_08441_),
    .B1(_08442_),
    .X(_08443_));
 sky130_fd_sc_hd__a31o_1 _13548_ (.A1(net796),
    .A2(_08439_),
    .A3(_08440_),
    .B1(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__a22oi_1 _13549_ (.A1(_07964_),
    .A2(_07965_),
    .B1(_07966_),
    .B2(_07975_),
    .Y(_08445_));
 sky130_fd_sc_hd__o31a_1 _13550_ (.A1(_07976_),
    .A2(net1224),
    .A3(_08445_),
    .B1(net781),
    .X(_08446_));
 sky130_fd_sc_hd__a21bo_1 _13551_ (.A1(\core.csr.traps.mtvec.csrReadData[6] ),
    .A2(net1224),
    .B1_N(_08446_),
    .X(_08447_));
 sky130_fd_sc_hd__and3_2 _13552_ (.A(net1774),
    .B(_08444_),
    .C(_08447_),
    .X(_08448_));
 sky130_fd_sc_hd__a21oi_4 _13553_ (.A1(net1764),
    .A2(\core.fetchProgramCounter[6] ),
    .B1(_08448_),
    .Y(_08449_));
 sky130_fd_sc_hd__nor2_2 _13554_ (.A(net1970),
    .B(_08449_),
    .Y(_08450_));
 sky130_fd_sc_hd__a22o_4 _13555_ (.A1(net720),
    .A2(_08438_),
    .B1(_08450_),
    .B2(net728),
    .X(net329));
 sky130_fd_sc_hd__nand2_1 _13556_ (.A(net1764),
    .B(\core.fetchProgramCounter[7] ),
    .Y(_08451_));
 sky130_fd_sc_hd__a21oi_2 _13557_ (.A1(_07606_),
    .A2(_07609_),
    .B1(_07556_),
    .Y(_08452_));
 sky130_fd_sc_hd__xnor2_2 _13558_ (.A(_07608_),
    .B(_08452_),
    .Y(_08453_));
 sky130_fd_sc_hd__xnor2_1 _13559_ (.A(\core.fetchProgramCounter[7] ),
    .B(_07897_),
    .Y(_08454_));
 sky130_fd_sc_hd__a221o_1 _13560_ (.A1(\core.csr.trapReturnVector[7] ),
    .A2(net1181),
    .B1(net787),
    .B2(_08454_),
    .C1(net782),
    .X(_08455_));
 sky130_fd_sc_hd__a21oi_2 _13561_ (.A1(net796),
    .A2(_08453_),
    .B1(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__a211o_1 _13562_ (.A1(_07961_),
    .A2(_07962_),
    .B1(_07963_),
    .C1(_07976_),
    .X(_08457_));
 sky130_fd_sc_hd__or3b_2 _13563_ (.A(_07977_),
    .B(net1224),
    .C_N(_08457_),
    .X(_08458_));
 sky130_fd_sc_hd__nand2_1 _13564_ (.A(\core.csr.traps.mtvec.csrReadData[7] ),
    .B(net1224),
    .Y(_08459_));
 sky130_fd_sc_hd__a311o_4 _13565_ (.A1(net780),
    .A2(_08458_),
    .A3(_08459_),
    .B1(_08456_),
    .C1(net1764),
    .X(_08460_));
 sky130_fd_sc_hd__a21oi_4 _13566_ (.A1(_08451_),
    .A2(_08460_),
    .B1(net1989),
    .Y(_08461_));
 sky130_fd_sc_hd__xor2_4 _13567_ (.A(_05633_),
    .B(_08061_),
    .X(_08462_));
 sky130_fd_sc_hd__inv_2 _13568_ (.A(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__a22o_4 _13569_ (.A1(_00577_),
    .A2(_08461_),
    .B1(_08463_),
    .B2(net720),
    .X(net330));
 sky130_fd_sc_hd__xnor2_4 _13570_ (.A(_06315_),
    .B(_08062_),
    .Y(_08464_));
 sky130_fd_sc_hd__nor2_1 _13571_ (.A(_07613_),
    .B(_07692_),
    .Y(_08465_));
 sky130_fd_sc_hd__or2_1 _13572_ (.A(_08184_),
    .B(_08465_),
    .X(_08466_));
 sky130_fd_sc_hd__a21oi_2 _13573_ (.A1(_07403_),
    .A2(_08466_),
    .B1(net798),
    .Y(_08467_));
 sky130_fd_sc_hd__a31o_1 _13574_ (.A1(\core.fetchProgramCounter[7] ),
    .A2(\core.fetchProgramCounter[6] ),
    .A3(_07896_),
    .B1(\core.fetchProgramCounter[8] ),
    .X(_08468_));
 sky130_fd_sc_hd__and3b_1 _13575_ (.A_N(_07898_),
    .B(_08468_),
    .C(net787),
    .X(_08469_));
 sky130_fd_sc_hd__a211o_1 _13576_ (.A1(\core.csr.trapReturnVector[8] ),
    .A2(net1180),
    .B1(_08469_),
    .C1(net779),
    .X(_08470_));
 sky130_fd_sc_hd__a21oi_1 _13577_ (.A1(_07959_),
    .A2(_07960_),
    .B1(_07978_),
    .Y(_08471_));
 sky130_fd_sc_hd__a31o_1 _13578_ (.A1(_07959_),
    .A2(_07960_),
    .A3(_07978_),
    .B1(net1224),
    .X(_08472_));
 sky130_fd_sc_hd__a2bb2o_2 _13579_ (.A1_N(_08471_),
    .A2_N(_08472_),
    .B1(\core.csr.traps.mtvec.csrReadData[8] ),
    .B2(net1224),
    .X(_08473_));
 sky130_fd_sc_hd__o21a_1 _13580_ (.A1(_08467_),
    .A2(_08470_),
    .B1(net1774),
    .X(_08474_));
 sky130_fd_sc_hd__o21ai_4 _13581_ (.A1(net767),
    .A2(_08473_),
    .B1(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__nand2_1 _13582_ (.A(net1764),
    .B(\core.fetchProgramCounter[8] ),
    .Y(_08476_));
 sky130_fd_sc_hd__a21oi_4 _13583_ (.A1(_08475_),
    .A2(_08476_),
    .B1(net1980),
    .Y(_08477_));
 sky130_fd_sc_hd__a22o_4 _13584_ (.A1(net720),
    .A2(_08464_),
    .B1(_08477_),
    .B2(net729),
    .X(net331));
 sky130_fd_sc_hd__o21ai_1 _13585_ (.A1(_07690_),
    .A2(_08184_),
    .B1(_07701_),
    .Y(_08478_));
 sky130_fd_sc_hd__or3_1 _13586_ (.A(_07690_),
    .B(_07701_),
    .C(_08184_),
    .X(_08479_));
 sky130_fd_sc_hd__xor2_1 _13587_ (.A(\core.fetchProgramCounter[9] ),
    .B(_07898_),
    .X(_08480_));
 sky130_fd_sc_hd__a221o_1 _13588_ (.A1(\core.csr.trapReturnVector[9] ),
    .A2(net1180),
    .B1(net787),
    .B2(_08480_),
    .C1(net778),
    .X(_08481_));
 sky130_fd_sc_hd__a31o_1 _13589_ (.A1(net795),
    .A2(_08478_),
    .A3(_08479_),
    .B1(_08481_),
    .X(_08482_));
 sky130_fd_sc_hd__nor2_1 _13590_ (.A(_07957_),
    .B(_07958_),
    .Y(_08483_));
 sky130_fd_sc_hd__xnor2_1 _13591_ (.A(_07979_),
    .B(_08483_),
    .Y(_08484_));
 sky130_fd_sc_hd__mux2_2 _13592_ (.A0(_08484_),
    .A1(\core.csr.traps.mtvec.csrReadData[9] ),
    .S(net1223),
    .X(_08485_));
 sky130_fd_sc_hd__o211a_1 _13593_ (.A1(net767),
    .A2(_08485_),
    .B1(_08482_),
    .C1(net1773),
    .X(_08486_));
 sky130_fd_sc_hd__a21oi_2 _13594_ (.A1(net1765),
    .A2(\core.fetchProgramCounter[9] ),
    .B1(_08486_),
    .Y(_08487_));
 sky130_fd_sc_hd__nor2_2 _13595_ (.A(net1979),
    .B(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__xor2_4 _13596_ (.A(_05551_),
    .B(_08063_),
    .X(_08489_));
 sky130_fd_sc_hd__a22o_4 _13597_ (.A1(net728),
    .A2(_08488_),
    .B1(_08489_),
    .B2(net720),
    .X(net332));
 sky130_fd_sc_hd__a21oi_1 _13598_ (.A1(\core.csr.trapReturnVector[10] ),
    .A2(net1181),
    .B1(net778),
    .Y(_08490_));
 sky130_fd_sc_hd__a21oi_1 _13599_ (.A1(\core.fetchProgramCounter[9] ),
    .A2(_07898_),
    .B1(\core.fetchProgramCounter[10] ),
    .Y(_08491_));
 sky130_fd_sc_hd__xor2_1 _13600_ (.A(_07682_),
    .B(_08185_),
    .X(_08492_));
 sky130_fd_sc_hd__a21oi_1 _13601_ (.A1(_07403_),
    .A2(_08492_),
    .B1(net798),
    .Y(_08493_));
 sky130_fd_sc_hd__o31a_1 _13602_ (.A1(net1180),
    .A2(_07899_),
    .A3(_08491_),
    .B1(net798),
    .X(_08494_));
 sky130_fd_sc_hd__or2_2 _13603_ (.A(_08493_),
    .B(_08494_),
    .X(_08495_));
 sky130_fd_sc_hd__nand2b_1 _13604_ (.A_N(_07955_),
    .B(_07956_),
    .Y(_08496_));
 sky130_fd_sc_hd__nor2_1 _13605_ (.A(_07980_),
    .B(_08496_),
    .Y(_08497_));
 sky130_fd_sc_hd__a211o_1 _13606_ (.A1(_07980_),
    .A2(_08496_),
    .B1(_08497_),
    .C1(net1225),
    .X(_08498_));
 sky130_fd_sc_hd__nand2_1 _13607_ (.A(\core.csr.traps.mtvec.csrReadData[10] ),
    .B(net1223),
    .Y(_08499_));
 sky130_fd_sc_hd__a32o_1 _13608_ (.A1(net778),
    .A2(_08498_),
    .A3(_08499_),
    .B1(_08490_),
    .B2(_08495_),
    .X(_08500_));
 sky130_fd_sc_hd__nand2_1 _13609_ (.A(net1773),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__o211a_2 _13610_ (.A1(net1772),
    .A2(\core.fetchProgramCounter[10] ),
    .B1(net1913),
    .C1(_08501_),
    .X(_08502_));
 sky130_fd_sc_hd__xnor2_4 _13611_ (.A(_05455_),
    .B(_08064_),
    .Y(_08503_));
 sky130_fd_sc_hd__and2_1 _13612_ (.A(net806),
    .B(_08503_),
    .X(_08504_));
 sky130_fd_sc_hd__a22o_4 _13613_ (.A1(net728),
    .A2(_08502_),
    .B1(_08504_),
    .B2(net723),
    .X(net306));
 sky130_fd_sc_hd__a22o_4 _13614_ (.A1(net728),
    .A2(_08366_),
    .B1(_08367_),
    .B2(net723),
    .X(net307));
 sky130_fd_sc_hd__a22o_2 _13615_ (.A1(net726),
    .A2(_08228_),
    .B1(_08333_),
    .B2(net719),
    .X(net308));
 sky130_fd_sc_hd__a22o_2 _13616_ (.A1(net726),
    .A2(_08203_),
    .B1(_08332_),
    .B2(net719),
    .X(net309));
 sky130_fd_sc_hd__a22o_2 _13617_ (.A1(net726),
    .A2(_08295_),
    .B1(_08331_),
    .B2(net719),
    .X(net310));
 sky130_fd_sc_hd__a22o_2 _13618_ (.A1(net726),
    .A2(_08318_),
    .B1(_08330_),
    .B2(net719),
    .X(net311));
 sky130_fd_sc_hd__a22o_2 _13619_ (.A1(net726),
    .A2(_08267_),
    .B1(_08329_),
    .B2(net719),
    .X(net312));
 sky130_fd_sc_hd__a22o_2 _13620_ (.A1(net726),
    .A2(_08253_),
    .B1(_08328_),
    .B2(net719),
    .X(net313));
 sky130_fd_sc_hd__a22o_2 _13621_ (.A1(net726),
    .A2(_08239_),
    .B1(_08327_),
    .B2(net719),
    .X(net314));
 sky130_fd_sc_hd__a22o_2 _13622_ (.A1(net727),
    .A2(_08216_),
    .B1(_08326_),
    .B2(net719),
    .X(net315));
 sky130_fd_sc_hd__a22o_2 _13623_ (.A1(net726),
    .A2(_08282_),
    .B1(_08325_),
    .B2(net719),
    .X(net317));
 sky130_fd_sc_hd__a22o_2 _13624_ (.A1(net726),
    .A2(_08183_),
    .B1(_08323_),
    .B2(net720),
    .X(net318));
 sky130_fd_sc_hd__o2bb2ai_4 _13625_ (.A1_N(net727),
    .A2_N(_08308_),
    .B1(_08322_),
    .B2(_08381_),
    .Y(net319));
 sky130_fd_sc_hd__a22o_4 _13626_ (.A1(net726),
    .A2(_08171_),
    .B1(_08321_),
    .B2(net719),
    .X(net320));
 sky130_fd_sc_hd__a22o_4 _13627_ (.A1(net729),
    .A2(_08114_),
    .B1(_08342_),
    .B2(net718),
    .X(net321));
 sky130_fd_sc_hd__a22o_4 _13628_ (.A1(net729),
    .A2(_08148_),
    .B1(_08341_),
    .B2(net718),
    .X(net322));
 sky130_fd_sc_hd__a22o_4 _13629_ (.A1(net729),
    .A2(_08138_),
    .B1(_08340_),
    .B2(net718),
    .X(net323));
 sky130_fd_sc_hd__a22o_4 _13630_ (.A1(net729),
    .A2(_08128_),
    .B1(_08339_),
    .B2(net718),
    .X(net324));
 sky130_fd_sc_hd__nor2_8 _13631_ (.A(_07477_),
    .B(_08096_),
    .Y(_08505_));
 sky130_fd_sc_hd__a31o_4 _13632_ (.A1(net765),
    .A2(_08099_),
    .A3(_08505_),
    .B1(net729),
    .X(net366));
 sky130_fd_sc_hd__o211a_4 _13633_ (.A1(_06697_),
    .A2(_07369_),
    .B1(_07475_),
    .C1(net807),
    .X(_08506_));
 sky130_fd_sc_hd__a31o_2 _13634_ (.A1(net765),
    .A2(_08099_),
    .A3(_08506_),
    .B1(net729),
    .X(net367));
 sky130_fd_sc_hd__or2_1 _13635_ (.A(_04465_),
    .B(net817),
    .X(_08507_));
 sky130_fd_sc_hd__nand2_8 _13636_ (.A(_06137_),
    .B(_06697_),
    .Y(_08508_));
 sky130_fd_sc_hd__and3_4 _13637_ (.A(net831),
    .B(net807),
    .C(_08507_),
    .X(_08509_));
 sky130_fd_sc_hd__a31o_2 _13638_ (.A1(net765),
    .A2(_08099_),
    .A3(_08509_),
    .B1(net729),
    .X(net368));
 sky130_fd_sc_hd__o311a_4 _13639_ (.A1(_06697_),
    .A2(_07369_),
    .A3(_07475_),
    .B1(net807),
    .C1(_08507_),
    .X(_08510_));
 sky130_fd_sc_hd__a31o_2 _13640_ (.A1(net765),
    .A2(_08099_),
    .A3(_08510_),
    .B1(net729),
    .X(net369));
 sky130_fd_sc_hd__nand2_2 _13641_ (.A(net1241),
    .B(_06191_),
    .Y(_08511_));
 sky130_fd_sc_hd__inv_6 _13642_ (.A(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__and3_4 _13643_ (.A(net812),
    .B(net723),
    .C(_08512_),
    .X(net334));
 sky130_fd_sc_hd__nor2_8 _13644_ (.A(_04482_),
    .B(_06096_),
    .Y(_08513_));
 sky130_fd_sc_hd__and3_4 _13645_ (.A(net812),
    .B(net723),
    .C(_08513_),
    .X(net345));
 sky130_fd_sc_hd__nor2_8 _13646_ (.A(_04482_),
    .B(_06011_),
    .Y(_08514_));
 sky130_fd_sc_hd__and3_4 _13647_ (.A(net812),
    .B(net723),
    .C(_08514_),
    .X(net356));
 sky130_fd_sc_hd__and2_4 _13648_ (.A(net1241),
    .B(_05926_),
    .X(_08515_));
 sky130_fd_sc_hd__and3_4 _13649_ (.A(net812),
    .B(net723),
    .C(_08515_),
    .X(net359));
 sky130_fd_sc_hd__nor2_8 _13650_ (.A(_04482_),
    .B(_05842_),
    .Y(_08516_));
 sky130_fd_sc_hd__nand2_1 _13651_ (.A(net828),
    .B(_08516_),
    .Y(_08517_));
 sky130_fd_sc_hd__and3_4 _13652_ (.A(net812),
    .B(net723),
    .C(_08516_),
    .X(net360));
 sky130_fd_sc_hd__nand2_2 _13653_ (.A(net1241),
    .B(_05761_),
    .Y(_08518_));
 sky130_fd_sc_hd__or2_4 _13654_ (.A(_06697_),
    .B(_08518_),
    .X(_08519_));
 sky130_fd_sc_hd__nor2_8 _13655_ (.A(net815),
    .B(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__and2_1 _13656_ (.A(net722),
    .B(_08520_),
    .X(net361));
 sky130_fd_sc_hd__or2_4 _13657_ (.A(_04482_),
    .B(_05676_),
    .X(_08521_));
 sky130_fd_sc_hd__or2_4 _13658_ (.A(_06697_),
    .B(_08521_),
    .X(_08522_));
 sky130_fd_sc_hd__nor2_8 _13659_ (.A(net816),
    .B(_08522_),
    .Y(_08523_));
 sky130_fd_sc_hd__and2_1 _13660_ (.A(net722),
    .B(_08523_),
    .X(net362));
 sky130_fd_sc_hd__nand2_2 _13661_ (.A(_04483_),
    .B(_05595_),
    .Y(_08524_));
 sky130_fd_sc_hd__inv_6 _13662_ (.A(_08524_),
    .Y(_08525_));
 sky130_fd_sc_hd__and3_4 _13663_ (.A(net812),
    .B(net723),
    .C(_08525_),
    .X(net363));
 sky130_fd_sc_hd__and2_4 _13664_ (.A(_06279_),
    .B(_07478_),
    .X(_08526_));
 sky130_fd_sc_hd__inv_2 _13665_ (.A(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__nor2_1 _13666_ (.A(net827),
    .B(_08512_),
    .Y(_08528_));
 sky130_fd_sc_hd__a211o_4 _13667_ (.A1(net827),
    .A2(_08527_),
    .B1(_08528_),
    .C1(net815),
    .X(_08529_));
 sky130_fd_sc_hd__inv_2 _13668_ (.A(_08529_),
    .Y(_08530_));
 sky130_fd_sc_hd__nor2_1 _13669_ (.A(_08381_),
    .B(_08529_),
    .Y(net364));
 sky130_fd_sc_hd__o211ai_4 _13670_ (.A1(net1154),
    .A2(net965),
    .B1(_05508_),
    .C1(_07478_),
    .Y(_08531_));
 sky130_fd_sc_hd__nor2_1 _13671_ (.A(net827),
    .B(_08513_),
    .Y(_08532_));
 sky130_fd_sc_hd__a211o_4 _13672_ (.A1(net827),
    .A2(_08531_),
    .B1(_08532_),
    .C1(net815),
    .X(_08533_));
 sky130_fd_sc_hd__inv_2 _13673_ (.A(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__nor2_1 _13674_ (.A(_08381_),
    .B(_08533_),
    .Y(net365));
 sky130_fd_sc_hd__nand4_4 _13675_ (.A(net1266),
    .B(_05388_),
    .C(_05418_),
    .D(_07478_),
    .Y(_08535_));
 sky130_fd_sc_hd__nor2_1 _13676_ (.A(net827),
    .B(_08514_),
    .Y(_08536_));
 sky130_fd_sc_hd__a211o_4 _13677_ (.A1(net827),
    .A2(_08535_),
    .B1(_08536_),
    .C1(net815),
    .X(_08537_));
 sky130_fd_sc_hd__inv_2 _13678_ (.A(_08537_),
    .Y(_08538_));
 sky130_fd_sc_hd__nor2_1 _13679_ (.A(_08381_),
    .B(_08537_),
    .Y(net335));
 sky130_fd_sc_hd__nand2_4 _13680_ (.A(_05362_),
    .B(_07478_),
    .Y(_08539_));
 sky130_fd_sc_hd__nor2_2 _13681_ (.A(net827),
    .B(_08515_),
    .Y(_08540_));
 sky130_fd_sc_hd__a211oi_4 _13682_ (.A1(net827),
    .A2(_08539_),
    .B1(_08540_),
    .C1(net815),
    .Y(_08541_));
 sky130_fd_sc_hd__and2_1 _13683_ (.A(net722),
    .B(_08541_),
    .X(net336));
 sky130_fd_sc_hd__nand2_4 _13684_ (.A(_04989_),
    .B(_07478_),
    .Y(_08542_));
 sky130_fd_sc_hd__nor2_2 _13685_ (.A(net828),
    .B(_08516_),
    .Y(_08543_));
 sky130_fd_sc_hd__a211oi_4 _13686_ (.A1(net828),
    .A2(_08542_),
    .B1(_08543_),
    .C1(net815),
    .Y(_08544_));
 sky130_fd_sc_hd__and2_1 _13687_ (.A(net718),
    .B(_08544_),
    .X(net337));
 sky130_fd_sc_hd__or2_4 _13688_ (.A(_05076_),
    .B(_07479_),
    .X(_08545_));
 sky130_fd_sc_hd__and3_2 _13689_ (.A(_06695_),
    .B(_06696_),
    .C(_08518_),
    .X(_08546_));
 sky130_fd_sc_hd__a211o_4 _13690_ (.A1(net829),
    .A2(_08545_),
    .B1(_08546_),
    .C1(net816),
    .X(_08547_));
 sky130_fd_sc_hd__inv_2 _13691_ (.A(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__nor2_1 _13692_ (.A(_08381_),
    .B(_08547_),
    .Y(net338));
 sky130_fd_sc_hd__or2_2 _13693_ (.A(_05242_),
    .B(_07479_),
    .X(_08549_));
 sky130_fd_sc_hd__and3_2 _13694_ (.A(_06695_),
    .B(_06696_),
    .C(_08521_),
    .X(_08550_));
 sky130_fd_sc_hd__a211o_4 _13695_ (.A1(net830),
    .A2(_08549_),
    .B1(_08550_),
    .C1(net817),
    .X(_08551_));
 sky130_fd_sc_hd__inv_2 _13696_ (.A(_08551_),
    .Y(_08552_));
 sky130_fd_sc_hd__nor2_1 _13697_ (.A(_08381_),
    .B(_08551_),
    .Y(net339));
 sky130_fd_sc_hd__or2_4 _13698_ (.A(_05155_),
    .B(_07479_),
    .X(_08553_));
 sky130_fd_sc_hd__nor2_1 _13699_ (.A(net829),
    .B(_08525_),
    .Y(_08554_));
 sky130_fd_sc_hd__a211o_4 _13700_ (.A1(net829),
    .A2(_08553_),
    .B1(_08554_),
    .C1(net816),
    .X(_08555_));
 sky130_fd_sc_hd__inv_2 _13701_ (.A(_08555_),
    .Y(_08556_));
 sky130_fd_sc_hd__nor2_1 _13702_ (.A(_08381_),
    .B(_08555_),
    .Y(net340));
 sky130_fd_sc_hd__nor2_1 _13703_ (.A(_06448_),
    .B(net1176),
    .Y(_08557_));
 sky130_fd_sc_hd__a22o_1 _13704_ (.A1(net830),
    .A2(_08512_),
    .B1(_08526_),
    .B2(_07475_),
    .X(_08558_));
 sky130_fd_sc_hd__mux2_8 _13705_ (.A0(_08557_),
    .A1(_08558_),
    .S(_07477_),
    .X(_08559_));
 sky130_fd_sc_hd__and2_1 _13706_ (.A(net721),
    .B(_08559_),
    .X(net341));
 sky130_fd_sc_hd__or2_2 _13707_ (.A(_06368_),
    .B(net1175),
    .X(_08560_));
 sky130_fd_sc_hd__nand2_1 _13708_ (.A(net827),
    .B(_08513_),
    .Y(_08561_));
 sky130_fd_sc_hd__o211a_1 _13709_ (.A1(net815),
    .A2(_08531_),
    .B1(_08561_),
    .C1(_07477_),
    .X(_08562_));
 sky130_fd_sc_hd__a21oi_4 _13710_ (.A1(net813),
    .A2(_08560_),
    .B1(_08562_),
    .Y(_08563_));
 sky130_fd_sc_hd__and2_1 _13711_ (.A(net721),
    .B(_08563_),
    .X(net342));
 sky130_fd_sc_hd__or2_1 _13712_ (.A(_06603_),
    .B(net1176),
    .X(_08564_));
 sky130_fd_sc_hd__o2bb2a_1 _13713_ (.A1_N(net828),
    .A2_N(_08514_),
    .B1(_08535_),
    .B2(net815),
    .X(_08565_));
 sky130_fd_sc_hd__mux2_8 _13714_ (.A0(_08564_),
    .A1(_08565_),
    .S(_07477_),
    .X(_08566_));
 sky130_fd_sc_hd__inv_2 _13715_ (.A(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__nor2_1 _13716_ (.A(_08381_),
    .B(_08566_),
    .Y(net343));
 sky130_fd_sc_hd__or2_2 _13717_ (.A(_06526_),
    .B(net1175),
    .X(_08568_));
 sky130_fd_sc_hd__nand2_1 _13718_ (.A(net827),
    .B(_08515_),
    .Y(_08569_));
 sky130_fd_sc_hd__o211a_1 _13719_ (.A1(net815),
    .A2(_08539_),
    .B1(_08569_),
    .C1(_07477_),
    .X(_08570_));
 sky130_fd_sc_hd__a21oi_4 _13720_ (.A1(net812),
    .A2(_08568_),
    .B1(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__and2_1 _13721_ (.A(net721),
    .B(_08571_),
    .X(net344));
 sky130_fd_sc_hd__or2_2 _13722_ (.A(_04895_),
    .B(net1175),
    .X(_08572_));
 sky130_fd_sc_hd__o211a_1 _13723_ (.A1(net815),
    .A2(_08542_),
    .B1(_08517_),
    .C1(_07477_),
    .X(_08573_));
 sky130_fd_sc_hd__a21oi_4 _13724_ (.A1(net813),
    .A2(_08572_),
    .B1(_08573_),
    .Y(_08574_));
 sky130_fd_sc_hd__and2_1 _13725_ (.A(net721),
    .B(_08574_),
    .X(net346));
 sky130_fd_sc_hd__or2_4 _13726_ (.A(_04818_),
    .B(net1175),
    .X(_08575_));
 sky130_fd_sc_hd__o211a_1 _13727_ (.A1(net816),
    .A2(_08545_),
    .B1(_08519_),
    .C1(_07477_),
    .X(_08576_));
 sky130_fd_sc_hd__a21oi_4 _13728_ (.A1(net814),
    .A2(_08575_),
    .B1(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__and2_1 _13729_ (.A(net721),
    .B(_08577_),
    .X(net347));
 sky130_fd_sc_hd__or2_2 _13730_ (.A(_04738_),
    .B(net1176),
    .X(_08578_));
 sky130_fd_sc_hd__o211a_1 _13731_ (.A1(net817),
    .A2(_08549_),
    .B1(_08522_),
    .C1(_07477_),
    .X(_08579_));
 sky130_fd_sc_hd__a21oi_4 _13732_ (.A1(net813),
    .A2(_08578_),
    .B1(_08579_),
    .Y(_08580_));
 sky130_fd_sc_hd__and2_1 _13733_ (.A(net721),
    .B(_08580_),
    .X(net348));
 sky130_fd_sc_hd__or2_4 _13734_ (.A(_04638_),
    .B(net1175),
    .X(_08581_));
 sky130_fd_sc_hd__nand2_1 _13735_ (.A(net829),
    .B(_08525_),
    .Y(_08582_));
 sky130_fd_sc_hd__o211a_1 _13736_ (.A1(net816),
    .A2(_08553_),
    .B1(_08582_),
    .C1(_07477_),
    .X(_08583_));
 sky130_fd_sc_hd__a21oi_4 _13737_ (.A1(net814),
    .A2(_08581_),
    .B1(_08583_),
    .Y(_08584_));
 sky130_fd_sc_hd__and2_1 _13738_ (.A(net721),
    .B(_08584_),
    .X(net349));
 sky130_fd_sc_hd__o21a_2 _13739_ (.A1(_06755_),
    .A2(net1175),
    .B1(net812),
    .X(_08585_));
 sky130_fd_sc_hd__nand2_8 _13740_ (.A(net830),
    .B(net817),
    .Y(_08586_));
 sky130_fd_sc_hd__nand2_8 _13741_ (.A(_08508_),
    .B(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__or3_1 _13742_ (.A(_06448_),
    .B(net1175),
    .C(_08508_),
    .X(_08588_));
 sky130_fd_sc_hd__o221a_4 _13743_ (.A1(_08527_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08528_),
    .C1(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__nor2_8 _13744_ (.A(_08585_),
    .B(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__and2_2 _13745_ (.A(net718),
    .B(_08590_),
    .X(net350));
 sky130_fd_sc_hd__o21a_2 _13746_ (.A1(_06834_),
    .A2(net1175),
    .B1(net812),
    .X(_08591_));
 sky130_fd_sc_hd__or2_1 _13747_ (.A(_08508_),
    .B(_08560_),
    .X(_08592_));
 sky130_fd_sc_hd__o221a_4 _13748_ (.A1(_08531_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08532_),
    .C1(_08592_),
    .X(_08593_));
 sky130_fd_sc_hd__nor2_8 _13749_ (.A(_08591_),
    .B(_08593_),
    .Y(_08594_));
 sky130_fd_sc_hd__and2_2 _13750_ (.A(net718),
    .B(_08594_),
    .X(net351));
 sky130_fd_sc_hd__o21a_2 _13751_ (.A1(_06988_),
    .A2(net1176),
    .B1(net813),
    .X(_08595_));
 sky130_fd_sc_hd__or2_1 _13752_ (.A(_08508_),
    .B(_08564_),
    .X(_08596_));
 sky130_fd_sc_hd__o221a_4 _13753_ (.A1(_08535_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08536_),
    .C1(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__nor2_8 _13754_ (.A(_08595_),
    .B(_08597_),
    .Y(_08598_));
 sky130_fd_sc_hd__and2_1 _13755_ (.A(net721),
    .B(_08598_),
    .X(net352));
 sky130_fd_sc_hd__o21a_2 _13756_ (.A1(_06912_),
    .A2(net1175),
    .B1(net812),
    .X(_08599_));
 sky130_fd_sc_hd__or2_1 _13757_ (.A(_08508_),
    .B(_08568_),
    .X(_08600_));
 sky130_fd_sc_hd__o221a_4 _13758_ (.A1(_08539_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08540_),
    .C1(_08600_),
    .X(_08601_));
 sky130_fd_sc_hd__nor2_8 _13759_ (.A(_08599_),
    .B(_08601_),
    .Y(_08602_));
 sky130_fd_sc_hd__and2_2 _13760_ (.A(net718),
    .B(_08602_),
    .X(net353));
 sky130_fd_sc_hd__o21a_2 _13761_ (.A1(_07070_),
    .A2(net1175),
    .B1(net813),
    .X(_08603_));
 sky130_fd_sc_hd__or2_1 _13762_ (.A(_08508_),
    .B(_08572_),
    .X(_08604_));
 sky130_fd_sc_hd__o221a_4 _13763_ (.A1(_08542_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08543_),
    .C1(_08604_),
    .X(_08605_));
 sky130_fd_sc_hd__nor2_8 _13764_ (.A(_08603_),
    .B(_08605_),
    .Y(_08606_));
 sky130_fd_sc_hd__and2_2 _13765_ (.A(net718),
    .B(_08606_),
    .X(net354));
 sky130_fd_sc_hd__o21a_2 _13766_ (.A1(_07158_),
    .A2(net1176),
    .B1(net813),
    .X(_08607_));
 sky130_fd_sc_hd__or2_1 _13767_ (.A(_08508_),
    .B(_08575_),
    .X(_08608_));
 sky130_fd_sc_hd__o221a_4 _13768_ (.A1(_08545_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08546_),
    .C1(_08608_),
    .X(_08609_));
 sky130_fd_sc_hd__nor2_8 _13769_ (.A(_08607_),
    .B(_08609_),
    .Y(_08610_));
 sky130_fd_sc_hd__and2_1 _13770_ (.A(net721),
    .B(_08610_),
    .X(net355));
 sky130_fd_sc_hd__o21a_2 _13771_ (.A1(_07315_),
    .A2(net1176),
    .B1(net813),
    .X(_08611_));
 sky130_fd_sc_hd__or2_1 _13772_ (.A(_08508_),
    .B(_08578_),
    .X(_08612_));
 sky130_fd_sc_hd__o221a_4 _13773_ (.A1(_08549_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08550_),
    .C1(_08612_),
    .X(_08613_));
 sky130_fd_sc_hd__nor2_8 _13774_ (.A(_08611_),
    .B(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__and2_1 _13775_ (.A(net722),
    .B(_08614_),
    .X(net357));
 sky130_fd_sc_hd__o21a_2 _13776_ (.A1(_07241_),
    .A2(net1176),
    .B1(net813),
    .X(_08615_));
 sky130_fd_sc_hd__or2_1 _13777_ (.A(_08508_),
    .B(_08581_),
    .X(_08616_));
 sky130_fd_sc_hd__o221a_4 _13778_ (.A1(_08553_),
    .A2(_08586_),
    .B1(_08587_),
    .B2(_08554_),
    .C1(_08616_),
    .X(_08617_));
 sky130_fd_sc_hd__nor2_8 _13779_ (.A(_08615_),
    .B(_08617_),
    .Y(_08618_));
 sky130_fd_sc_hd__and2_1 _13780_ (.A(net721),
    .B(_08618_),
    .X(net358));
 sky130_fd_sc_hd__a32o_4 _13781_ (.A1(net806),
    .A2(net2010),
    .A3(_08382_),
    .B1(_08393_),
    .B2(_08152_),
    .X(net294));
 sky130_fd_sc_hd__a22o_4 _13782_ (.A1(net2010),
    .A2(_08396_),
    .B1(_08408_),
    .B2(net725),
    .X(net295));
 sky130_fd_sc_hd__a32o_4 _13783_ (.A1(net806),
    .A2(net724),
    .A3(_08422_),
    .B1(_08420_),
    .B2(net725),
    .X(net296));
 sky130_fd_sc_hd__a22o_4 _13784_ (.A1(net725),
    .A2(_08434_),
    .B1(_08436_),
    .B2(net2010),
    .X(net297));
 sky130_fd_sc_hd__a22o_4 _13785_ (.A1(net2010),
    .A2(_08438_),
    .B1(_08450_),
    .B2(net725),
    .X(net298));
 sky130_fd_sc_hd__a32o_4 _13786_ (.A1(net806),
    .A2(net724),
    .A3(_08463_),
    .B1(_08461_),
    .B2(_08152_),
    .X(net299));
 sky130_fd_sc_hd__a32o_4 _13787_ (.A1(net806),
    .A2(_08346_),
    .A3(_08464_),
    .B1(_08477_),
    .B2(_08152_),
    .X(net300));
 sky130_fd_sc_hd__a32o_4 _13788_ (.A1(net806),
    .A2(_08346_),
    .A3(_08489_),
    .B1(_08488_),
    .B2(net725),
    .X(net301));
 sky130_fd_sc_hd__a22o_4 _13789_ (.A1(net725),
    .A2(_08502_),
    .B1(_08504_),
    .B2(_08346_),
    .X(net302));
 sky130_fd_sc_hd__and2_4 _13790_ (.A(_07865_),
    .B(net702),
    .X(_08619_));
 sky130_fd_sc_hd__a32o_2 _13791_ (.A1(net814),
    .A2(net707),
    .A3(_08512_),
    .B1(net690),
    .B2(net215),
    .X(net376));
 sky130_fd_sc_hd__a32o_2 _13792_ (.A1(net814),
    .A2(net707),
    .A3(_08513_),
    .B1(net690),
    .B2(net226),
    .X(net387));
 sky130_fd_sc_hd__a32o_1 _13793_ (.A1(net814),
    .A2(net707),
    .A3(_08514_),
    .B1(net690),
    .B2(net237),
    .X(net398));
 sky130_fd_sc_hd__a32o_1 _13794_ (.A1(net814),
    .A2(net707),
    .A3(_08515_),
    .B1(net690),
    .B2(net240),
    .X(net401));
 sky130_fd_sc_hd__a32o_1 _13795_ (.A1(net814),
    .A2(net708),
    .A3(_08516_),
    .B1(net691),
    .B2(net241),
    .X(net402));
 sky130_fd_sc_hd__a22o_1 _13796_ (.A1(net708),
    .A2(_08520_),
    .B1(net691),
    .B2(net242),
    .X(net403));
 sky130_fd_sc_hd__a22o_1 _13797_ (.A1(net707),
    .A2(_08523_),
    .B1(net690),
    .B2(net243),
    .X(net404));
 sky130_fd_sc_hd__a32o_1 _13798_ (.A1(net814),
    .A2(net707),
    .A3(_08525_),
    .B1(net690),
    .B2(net244),
    .X(net405));
 sky130_fd_sc_hd__a22o_1 _13799_ (.A1(net709),
    .A2(_08530_),
    .B1(net693),
    .B2(net245),
    .X(net406));
 sky130_fd_sc_hd__a22o_1 _13800_ (.A1(net709),
    .A2(_08534_),
    .B1(net692),
    .B2(net246),
    .X(net407));
 sky130_fd_sc_hd__a22o_1 _13801_ (.A1(net708),
    .A2(_08538_),
    .B1(net691),
    .B2(net216),
    .X(net377));
 sky130_fd_sc_hd__a22o_1 _13802_ (.A1(net708),
    .A2(_08541_),
    .B1(net691),
    .B2(net217),
    .X(net378));
 sky130_fd_sc_hd__a22o_1 _13803_ (.A1(net711),
    .A2(_08544_),
    .B1(_08619_),
    .B2(net218),
    .X(net379));
 sky130_fd_sc_hd__a22o_1 _13804_ (.A1(net711),
    .A2(_08548_),
    .B1(_08619_),
    .B2(net219),
    .X(net380));
 sky130_fd_sc_hd__a22o_1 _13805_ (.A1(net710),
    .A2(_08552_),
    .B1(net691),
    .B2(net220),
    .X(net381));
 sky130_fd_sc_hd__a22o_1 _13806_ (.A1(net710),
    .A2(_08556_),
    .B1(net692),
    .B2(net221),
    .X(net382));
 sky130_fd_sc_hd__a22o_2 _13807_ (.A1(net711),
    .A2(_08559_),
    .B1(_08619_),
    .B2(net222),
    .X(net383));
 sky130_fd_sc_hd__a22o_1 _13808_ (.A1(net709),
    .A2(_08563_),
    .B1(net692),
    .B2(net223),
    .X(net384));
 sky130_fd_sc_hd__a22o_1 _13809_ (.A1(net709),
    .A2(_08567_),
    .B1(net692),
    .B2(net224),
    .X(net385));
 sky130_fd_sc_hd__a22o_1 _13810_ (.A1(net710),
    .A2(_08571_),
    .B1(net693),
    .B2(net225),
    .X(net386));
 sky130_fd_sc_hd__a22o_1 _13811_ (.A1(net709),
    .A2(_08574_),
    .B1(net692),
    .B2(net227),
    .X(net388));
 sky130_fd_sc_hd__a22o_1 _13812_ (.A1(net709),
    .A2(_08577_),
    .B1(net692),
    .B2(net228),
    .X(net389));
 sky130_fd_sc_hd__a22o_1 _13813_ (.A1(net709),
    .A2(_08580_),
    .B1(net692),
    .B2(net229),
    .X(net390));
 sky130_fd_sc_hd__a22o_1 _13814_ (.A1(net709),
    .A2(_08584_),
    .B1(net692),
    .B2(net230),
    .X(net391));
 sky130_fd_sc_hd__a22o_1 _13815_ (.A1(net709),
    .A2(_08590_),
    .B1(net692),
    .B2(net231),
    .X(net392));
 sky130_fd_sc_hd__a22o_1 _13816_ (.A1(net709),
    .A2(_08594_),
    .B1(net692),
    .B2(net232),
    .X(net393));
 sky130_fd_sc_hd__a22o_1 _13817_ (.A1(net711),
    .A2(_08598_),
    .B1(net693),
    .B2(net233),
    .X(net394));
 sky130_fd_sc_hd__a22o_1 _13818_ (.A1(net711),
    .A2(_08602_),
    .B1(net2016),
    .B2(net234),
    .X(net395));
 sky130_fd_sc_hd__a22o_1 _13819_ (.A1(net711),
    .A2(_08606_),
    .B1(net2016),
    .B2(net235),
    .X(net396));
 sky130_fd_sc_hd__a22o_1 _13820_ (.A1(net711),
    .A2(_08610_),
    .B1(net2016),
    .B2(net236),
    .X(net397));
 sky130_fd_sc_hd__a22o_1 _13821_ (.A1(net711),
    .A2(_08614_),
    .B1(net2016),
    .B2(net238),
    .X(net399));
 sky130_fd_sc_hd__a22o_1 _13822_ (.A1(net711),
    .A2(_08618_),
    .B1(net2016),
    .B2(net239),
    .X(net400));
 sky130_fd_sc_hd__a22o_4 _13823_ (.A1(net707),
    .A2(_08505_),
    .B1(net690),
    .B2(\wbSRAMInterface.currentByteSelect[0] ),
    .X(net484));
 sky130_fd_sc_hd__a22o_4 _13824_ (.A1(net707),
    .A2(_08506_),
    .B1(net690),
    .B2(\wbSRAMInterface.currentByteSelect[1] ),
    .X(net485));
 sky130_fd_sc_hd__a22o_4 _13825_ (.A1(net707),
    .A2(_08509_),
    .B1(net690),
    .B2(\wbSRAMInterface.currentByteSelect[2] ),
    .X(net486));
 sky130_fd_sc_hd__a22o_4 _13826_ (.A1(net707),
    .A2(_08510_),
    .B1(net690),
    .B2(\wbSRAMInterface.currentByteSelect[3] ),
    .X(net487));
 sky130_fd_sc_hd__a22o_4 _13827_ (.A1(\wbSRAMInterface.currentAddress[2] ),
    .A2(net702),
    .B1(net294),
    .B2(net712),
    .X(net285));
 sky130_fd_sc_hd__a22o_4 _13828_ (.A1(\wbSRAMInterface.currentAddress[3] ),
    .A2(net702),
    .B1(net295),
    .B2(net712),
    .X(net286));
 sky130_fd_sc_hd__a22o_4 _13829_ (.A1(\wbSRAMInterface.currentAddress[4] ),
    .A2(net702),
    .B1(net296),
    .B2(net2009),
    .X(net287));
 sky130_fd_sc_hd__a22o_4 _13830_ (.A1(\wbSRAMInterface.currentAddress[5] ),
    .A2(_08378_),
    .B1(net297),
    .B2(net2009),
    .X(net288));
 sky130_fd_sc_hd__a22o_4 _13831_ (.A1(\wbSRAMInterface.currentAddress[6] ),
    .A2(_08378_),
    .B1(net298),
    .B2(net2009),
    .X(net289));
 sky130_fd_sc_hd__a22o_4 _13832_ (.A1(\wbSRAMInterface.currentAddress[7] ),
    .A2(net2008),
    .B1(net299),
    .B2(net713),
    .X(net290));
 sky130_fd_sc_hd__a22o_4 _13833_ (.A1(\wbSRAMInterface.currentAddress[8] ),
    .A2(net2008),
    .B1(net300),
    .B2(net713),
    .X(net291));
 sky130_fd_sc_hd__a22o_4 _13834_ (.A1(\wbSRAMInterface.currentAddress[9] ),
    .A2(net2008),
    .B1(net301),
    .B2(net2009),
    .X(net292));
 sky130_fd_sc_hd__a22o_4 _13835_ (.A1(\wbSRAMInterface.currentAddress[10] ),
    .A2(net2008),
    .B1(net302),
    .B2(net2009),
    .X(net293));
 sky130_fd_sc_hd__and2b_4 _13836_ (.A_N(\jtag.state[2] ),
    .B(\jtag.state[3] ),
    .X(_08620_));
 sky130_fd_sc_hd__and2_2 _13837_ (.A(net1778),
    .B(_08620_),
    .X(_08621_));
 sky130_fd_sc_hd__nand2_1 _13838_ (.A(net446),
    .B(net445),
    .Y(_08622_));
 sky130_fd_sc_hd__or4_4 _13839_ (.A(net449),
    .B(net448),
    .C(net447),
    .D(_08622_),
    .X(_08623_));
 sky130_fd_sc_hd__or4b_1 _13840_ (.A(net449),
    .B(net446),
    .C(net445),
    .D_N(net447),
    .X(_08624_));
 sky130_fd_sc_hd__o21a_2 _13841_ (.A1(net448),
    .A2(_08624_),
    .B1(_08623_),
    .X(_08625_));
 sky130_fd_sc_hd__and3_1 _13842_ (.A(net447),
    .B(net446),
    .C(net445),
    .X(_08626_));
 sky130_fd_sc_hd__and3_1 _13843_ (.A(net449),
    .B(net448),
    .C(_08626_),
    .X(_08627_));
 sky130_fd_sc_hd__or3b_1 _13844_ (.A(_08625_),
    .B(_08627_),
    .C_N(\jtag.dataIDRegister.data[31] ),
    .X(_08628_));
 sky130_fd_sc_hd__or3b_2 _13845_ (.A(net448),
    .B(net447),
    .C_N(net445),
    .X(_08629_));
 sky130_fd_sc_hd__nor3_4 _13846_ (.A(net449),
    .B(net446),
    .C(_08629_),
    .Y(_08630_));
 sky130_fd_sc_hd__a21bo_1 _13847_ (.A1(\jtag.dataBypassRegister.data ),
    .A2(_08627_),
    .B1_N(_08628_),
    .X(_08631_));
 sky130_fd_sc_hd__or2_1 _13848_ (.A(net1778),
    .B(net1780),
    .X(_08632_));
 sky130_fd_sc_hd__nand2b_2 _13849_ (.A_N(\jtag.state[3] ),
    .B(\jtag.state[2] ),
    .Y(_08633_));
 sky130_fd_sc_hd__nor2_2 _13850_ (.A(_08632_),
    .B(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__mux2_1 _13851_ (.A0(_08631_),
    .A1(\jtag.dataBSRRegister.data[31] ),
    .S(_08630_),
    .X(_08635_));
 sky130_fd_sc_hd__a32o_4 _13852_ (.A1(net1779),
    .A2(\jtag.instructionRegister.data[4] ),
    .A3(_08621_),
    .B1(_08634_),
    .B2(_08635_),
    .X(net408));
 sky130_fd_sc_hd__nand2_8 _13853_ (.A(\memoryController.last_instruction_enableWB ),
    .B(_04431_),
    .Y(_08636_));
 sky130_fd_sc_hd__a21oi_4 _13854_ (.A1(_07505_),
    .A2(_08101_),
    .B1(_08636_),
    .Y(_08637_));
 sky130_fd_sc_hd__a21oi_4 _13855_ (.A1(\memoryController.last_instruction_enableLocalMemory ),
    .A2(_08354_),
    .B1(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__a211o_4 _13856_ (.A1(\memoryController.last_instruction_enableLocalMemory ),
    .A2(_08354_),
    .B1(_08637_),
    .C1(_08052_),
    .X(_08639_));
 sky130_fd_sc_hd__a211oi_4 _13857_ (.A1(_08350_),
    .A2(_08353_),
    .B1(_04430_),
    .C1(\memoryController.last_instruction_enableLocalMemory ),
    .Y(_08640_));
 sky130_fd_sc_hd__a211oi_4 _13858_ (.A1(_07505_),
    .A2(_08101_),
    .B1(\memoryController.last_instruction_enableWB ),
    .C1(_04561_),
    .Y(_08641_));
 sky130_fd_sc_hd__or2_4 _13859_ (.A(_08640_),
    .B(_08641_),
    .X(_08642_));
 sky130_fd_sc_hd__or3_2 _13860_ (.A(_08097_),
    .B(_08640_),
    .C(_08641_),
    .X(_08643_));
 sky130_fd_sc_hd__o31a_4 _13861_ (.A1(_08097_),
    .A2(_08640_),
    .A3(_08641_),
    .B1(net1772),
    .X(_08644_));
 sky130_fd_sc_hd__and2_4 _13862_ (.A(_08639_),
    .B(net697),
    .X(_08645_));
 sky130_fd_sc_hd__nand2_1 _13863_ (.A(net1665),
    .B(net684),
    .Y(_08646_));
 sky130_fd_sc_hd__o221a_1 _13864_ (.A1(\core.csr.currentInstruction[0] ),
    .A2(net682),
    .B1(net631),
    .B2(\core.pipe0_currentInstruction[0] ),
    .C1(net1926),
    .X(_00000_));
 sky130_fd_sc_hd__o221a_1 _13865_ (.A1(\core.csr.currentInstruction[1] ),
    .A2(net684),
    .B1(net631),
    .B2(\core.pipe0_currentInstruction[1] ),
    .C1(net1922),
    .X(_00001_));
 sky130_fd_sc_hd__o221a_1 _13866_ (.A1(\core.csr.currentInstruction[2] ),
    .A2(net682),
    .B1(net630),
    .B2(\core.pipe0_currentInstruction[2] ),
    .C1(net1926),
    .X(_00002_));
 sky130_fd_sc_hd__nand2_1 _13867_ (.A(_04455_),
    .B(net677),
    .Y(_08647_));
 sky130_fd_sc_hd__o211a_1 _13868_ (.A1(\core.csr.currentInstruction[3] ),
    .A2(net677),
    .B1(_08647_),
    .C1(net1922),
    .X(_00003_));
 sky130_fd_sc_hd__nand2_1 _13869_ (.A(_04447_),
    .B(net677),
    .Y(_08648_));
 sky130_fd_sc_hd__o211a_1 _13870_ (.A1(\core.csr.currentInstruction[4] ),
    .A2(net677),
    .B1(_08648_),
    .C1(net1908),
    .X(_00004_));
 sky130_fd_sc_hd__o221a_1 _13871_ (.A1(\core.csr.currentInstruction[5] ),
    .A2(net684),
    .B1(net629),
    .B2(\core.pipe0_currentInstruction[5] ),
    .C1(net1928),
    .X(_00005_));
 sky130_fd_sc_hd__o221a_1 _13872_ (.A1(\core.csr.currentInstruction[6] ),
    .A2(net683),
    .B1(net629),
    .B2(\core.pipe0_currentInstruction[6] ),
    .C1(net1928),
    .X(_00006_));
 sky130_fd_sc_hd__o221a_1 _13873_ (.A1(\core.csr.currentInstruction[7] ),
    .A2(net682),
    .B1(net631),
    .B2(\core.pipe0_currentInstruction[7] ),
    .C1(net1926),
    .X(_00007_));
 sky130_fd_sc_hd__o221a_1 _13874_ (.A1(\core.csr.currentInstruction[8] ),
    .A2(net682),
    .B1(net631),
    .B2(\core.pipe0_currentInstruction[8] ),
    .C1(net1926),
    .X(_00008_));
 sky130_fd_sc_hd__o221a_1 _13875_ (.A1(\core.csr.currentInstruction[9] ),
    .A2(net682),
    .B1(net631),
    .B2(\core.pipe0_currentInstruction[9] ),
    .C1(net1926),
    .X(_00009_));
 sky130_fd_sc_hd__o221a_1 _13876_ (.A1(\core.csr.currentInstruction[10] ),
    .A2(net682),
    .B1(net631),
    .B2(\core.pipe0_currentInstruction[10] ),
    .C1(net1922),
    .X(_00010_));
 sky130_fd_sc_hd__o221a_1 _13877_ (.A1(\core.csr.currentInstruction[11] ),
    .A2(net682),
    .B1(net631),
    .B2(\core.pipe0_currentInstruction[11] ),
    .C1(net1922),
    .X(_00011_));
 sky130_fd_sc_hd__o221a_1 _13878_ (.A1(\core.csr.currentInstruction[12] ),
    .A2(net683),
    .B1(net630),
    .B2(net1882),
    .C1(net1927),
    .X(_00012_));
 sky130_fd_sc_hd__o221a_1 _13879_ (.A1(net1885),
    .A2(net683),
    .B1(net630),
    .B2(\core.pipe0_currentInstruction[13] ),
    .C1(net1927),
    .X(_00013_));
 sky130_fd_sc_hd__o221a_1 _13880_ (.A1(\core.csr.currentInstruction[14] ),
    .A2(net683),
    .B1(net630),
    .B2(\core.pipe0_currentInstruction[14] ),
    .C1(net1927),
    .X(_00014_));
 sky130_fd_sc_hd__o221a_1 _13881_ (.A1(\core.csr.currentInstruction[15] ),
    .A2(net682),
    .B1(net631),
    .B2(\core.pipe0_currentInstruction[15] ),
    .C1(net1922),
    .X(_00015_));
 sky130_fd_sc_hd__o221a_1 _13882_ (.A1(\core.csr.currentInstruction[16] ),
    .A2(net678),
    .B1(net632),
    .B2(net1871),
    .C1(net1907),
    .X(_00016_));
 sky130_fd_sc_hd__o221a_1 _13883_ (.A1(\core.csr.currentInstruction[17] ),
    .A2(net678),
    .B1(net632),
    .B2(net1867),
    .C1(net1906),
    .X(_00017_));
 sky130_fd_sc_hd__o221a_1 _13884_ (.A1(\core.csr.currentInstruction[18] ),
    .A2(net678),
    .B1(net632),
    .B2(\core.pipe0_currentInstruction[18] ),
    .C1(net1907),
    .X(_00018_));
 sky130_fd_sc_hd__o221a_1 _13885_ (.A1(\core.csr.currentInstruction[19] ),
    .A2(net678),
    .B1(net632),
    .B2(net1861),
    .C1(net1906),
    .X(_00019_));
 sky130_fd_sc_hd__o221a_1 _13886_ (.A1(\core.csr.currentInstruction[20] ),
    .A2(net678),
    .B1(net632),
    .B2(net1852),
    .C1(net1906),
    .X(_00020_));
 sky130_fd_sc_hd__o221a_1 _13887_ (.A1(\core.csr.currentInstruction[21] ),
    .A2(net678),
    .B1(net632),
    .B2(\core.pipe0_currentInstruction[21] ),
    .C1(net1919),
    .X(_00021_));
 sky130_fd_sc_hd__o221a_1 _13888_ (.A1(\core.csr.currentInstruction[22] ),
    .A2(net683),
    .B1(net629),
    .B2(net1837),
    .C1(net1928),
    .X(_00022_));
 sky130_fd_sc_hd__o221a_1 _13889_ (.A1(\core.csr.currentInstruction[23] ),
    .A2(net678),
    .B1(net632),
    .B2(net1831),
    .C1(net1906),
    .X(_00023_));
 sky130_fd_sc_hd__o221a_1 _13890_ (.A1(\core.csr.currentInstruction[24] ),
    .A2(net688),
    .B1(net629),
    .B2(net1828),
    .C1(net1946),
    .X(_00024_));
 sky130_fd_sc_hd__o221a_1 _13891_ (.A1(\core.csr.currentInstruction[25] ),
    .A2(net686),
    .B1(net629),
    .B2(net1822),
    .C1(net1943),
    .X(_00025_));
 sky130_fd_sc_hd__o221a_1 _13892_ (.A1(\core.csr.currentInstruction[26] ),
    .A2(net688),
    .B1(net629),
    .B2(net1821),
    .C1(net1943),
    .X(_00026_));
 sky130_fd_sc_hd__o221a_1 _13893_ (.A1(\core.csr.currentInstruction[27] ),
    .A2(net683),
    .B1(net629),
    .B2(net1820),
    .C1(net1943),
    .X(_00027_));
 sky130_fd_sc_hd__o221a_1 _13894_ (.A1(\core.csr.currentInstruction[28] ),
    .A2(net686),
    .B1(net629),
    .B2(net1819),
    .C1(net1943),
    .X(_00028_));
 sky130_fd_sc_hd__o221a_1 _13895_ (.A1(\core.csr.currentInstruction[29] ),
    .A2(net686),
    .B1(net629),
    .B2(\core.pipe0_currentInstruction[29] ),
    .C1(net1943),
    .X(_00029_));
 sky130_fd_sc_hd__o221a_1 _13896_ (.A1(\core.csr.currentInstruction[30] ),
    .A2(net683),
    .B1(net629),
    .B2(net1818),
    .C1(net1927),
    .X(_00030_));
 sky130_fd_sc_hd__or3b_1 _13897_ (.A(net1816),
    .B(net1668),
    .C_N(net683),
    .X(_08649_));
 sky130_fd_sc_hd__o211a_1 _13898_ (.A1(\core.csr.currentInstruction[31] ),
    .A2(net683),
    .B1(_08649_),
    .C1(net1928),
    .X(_00031_));
 sky130_fd_sc_hd__or2_4 _13899_ (.A(net1990),
    .B(net686),
    .X(_08650_));
 sky130_fd_sc_hd__o22a_1 _13900_ (.A1(net1990),
    .A2(net630),
    .B1(_08650_),
    .B2(net1884),
    .X(_00032_));
 sky130_fd_sc_hd__and3_1 _13901_ (.A(_07893_),
    .B(_08639_),
    .C(net697),
    .X(_08651_));
 sky130_fd_sc_hd__nand2_4 _13902_ (.A(_07893_),
    .B(net677),
    .Y(_08652_));
 sky130_fd_sc_hd__nor2_4 _13903_ (.A(net1970),
    .B(net674),
    .Y(_08653_));
 sky130_fd_sc_hd__a22o_1 _13904_ (.A1(_07443_),
    .A2(net674),
    .B1(_08653_),
    .B2(\core.csr.instruction_memoryAddress[0] ),
    .X(_00033_));
 sky130_fd_sc_hd__o22a_1 _13905_ (.A1(\core.csr.instruction_memoryAddress[1] ),
    .A2(net673),
    .B1(net624),
    .B2(_07437_),
    .X(_00034_));
 sky130_fd_sc_hd__and2_4 _13906_ (.A(net1906),
    .B(net673),
    .X(_08654_));
 sky130_fd_sc_hd__nand2_1 _13907_ (.A(_08392_),
    .B(net672),
    .Y(_08655_));
 sky130_fd_sc_hd__o211a_1 _13908_ (.A1(\core.csr.instruction_memoryAddress[2] ),
    .A2(net672),
    .B1(_08655_),
    .C1(net1913),
    .X(_00035_));
 sky130_fd_sc_hd__nand2_1 _13909_ (.A(_08407_),
    .B(net671),
    .Y(_08656_));
 sky130_fd_sc_hd__o211a_1 _13910_ (.A1(\core.csr.instruction_memoryAddress[3] ),
    .A2(net671),
    .B1(_08656_),
    .C1(net1914),
    .X(_00036_));
 sky130_fd_sc_hd__nand2_1 _13911_ (.A(_08419_),
    .B(net671),
    .Y(_08657_));
 sky130_fd_sc_hd__o211a_1 _13912_ (.A1(\core.csr.instruction_memoryAddress[4] ),
    .A2(net671),
    .B1(_08657_),
    .C1(net1913),
    .X(_00037_));
 sky130_fd_sc_hd__nand2_1 _13913_ (.A(_08433_),
    .B(net671),
    .Y(_08658_));
 sky130_fd_sc_hd__o211a_1 _13914_ (.A1(\core.csr.instruction_memoryAddress[5] ),
    .A2(net671),
    .B1(_08658_),
    .C1(net1930),
    .X(_00038_));
 sky130_fd_sc_hd__nand2_1 _13915_ (.A(_08449_),
    .B(net671),
    .Y(_08659_));
 sky130_fd_sc_hd__o211a_1 _13916_ (.A1(\core.csr.instruction_memoryAddress[6] ),
    .A2(net671),
    .B1(_08659_),
    .C1(net1930),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_1 _13917_ (.A0(\core.csr.instruction_memoryAddress[7] ),
    .A1(_08461_),
    .S(net671),
    .X(_08660_));
 sky130_fd_sc_hd__and2_1 _13918_ (.A(net1930),
    .B(_08660_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _13919_ (.A0(\core.csr.instruction_memoryAddress[8] ),
    .A1(_08477_),
    .S(net671),
    .X(_08661_));
 sky130_fd_sc_hd__and2_1 _13920_ (.A(net1930),
    .B(_08661_),
    .X(_00041_));
 sky130_fd_sc_hd__nand2_1 _13921_ (.A(_08487_),
    .B(net672),
    .Y(_08662_));
 sky130_fd_sc_hd__o211a_1 _13922_ (.A1(\core.csr.instruction_memoryAddress[9] ),
    .A2(net672),
    .B1(_08662_),
    .C1(net1913),
    .X(_00042_));
 sky130_fd_sc_hd__o22a_1 _13923_ (.A1(\core.csr.instruction_memoryAddress[10] ),
    .A2(net672),
    .B1(net624),
    .B2(_08502_),
    .X(_00043_));
 sky130_fd_sc_hd__o22a_1 _13924_ (.A1(\core.csr.instruction_memoryAddress[11] ),
    .A2(net672),
    .B1(net624),
    .B2(_08366_),
    .X(_00044_));
 sky130_fd_sc_hd__o22a_1 _13925_ (.A1(\core.csr.instruction_memoryAddress[12] ),
    .A2(net672),
    .B1(net624),
    .B2(_08228_),
    .X(_00045_));
 sky130_fd_sc_hd__o22a_1 _13926_ (.A1(\core.csr.instruction_memoryAddress[13] ),
    .A2(net673),
    .B1(_08653_),
    .B2(_08203_),
    .X(_00046_));
 sky130_fd_sc_hd__o22a_1 _13927_ (.A1(\core.csr.instruction_memoryAddress[14] ),
    .A2(net673),
    .B1(net624),
    .B2(_08295_),
    .X(_00047_));
 sky130_fd_sc_hd__o22a_1 _13928_ (.A1(\core.csr.instruction_memoryAddress[15] ),
    .A2(net673),
    .B1(net624),
    .B2(_08318_),
    .X(_00048_));
 sky130_fd_sc_hd__o22a_1 _13929_ (.A1(\core.csr.instruction_memoryAddress[16] ),
    .A2(net673),
    .B1(net624),
    .B2(_08267_),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_1 _13930_ (.A1(\core.csr.instruction_memoryAddress[17] ),
    .A2(net624),
    .B1(_08654_),
    .B2(_08253_),
    .X(_00050_));
 sky130_fd_sc_hd__o22a_1 _13931_ (.A1(\core.csr.instruction_memoryAddress[18] ),
    .A2(net674),
    .B1(net624),
    .B2(_08239_),
    .X(_00051_));
 sky130_fd_sc_hd__o22a_1 _13932_ (.A1(\core.csr.instruction_memoryAddress[19] ),
    .A2(net670),
    .B1(net624),
    .B2(_08216_),
    .X(_00052_));
 sky130_fd_sc_hd__o22a_1 _13933_ (.A1(\core.csr.instruction_memoryAddress[20] ),
    .A2(net670),
    .B1(net623),
    .B2(_08282_),
    .X(_00053_));
 sky130_fd_sc_hd__o22a_1 _13934_ (.A1(\core.csr.instruction_memoryAddress[21] ),
    .A2(net670),
    .B1(net623),
    .B2(_08183_),
    .X(_00054_));
 sky130_fd_sc_hd__o22a_1 _13935_ (.A1(\core.csr.instruction_memoryAddress[22] ),
    .A2(net670),
    .B1(net623),
    .B2(_08308_),
    .X(_00055_));
 sky130_fd_sc_hd__o22a_1 _13936_ (.A1(\core.csr.instruction_memoryAddress[23] ),
    .A2(net670),
    .B1(net623),
    .B2(_08171_),
    .X(_00056_));
 sky130_fd_sc_hd__o22a_1 _13937_ (.A1(\core.csr.instruction_memoryAddress[24] ),
    .A2(net670),
    .B1(net623),
    .B2(_08114_),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_1 _13938_ (.A1(\core.csr.instruction_memoryAddress[25] ),
    .A2(net623),
    .B1(_08654_),
    .B2(_08148_),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_1 _13939_ (.A1(\core.csr.instruction_memoryAddress[26] ),
    .A2(net623),
    .B1(_08654_),
    .B2(_08138_),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_1 _13940_ (.A1(\core.csr.instruction_memoryAddress[27] ),
    .A2(net623),
    .B1(_08654_),
    .B2(_08128_),
    .X(_00060_));
 sky130_fd_sc_hd__nand2_1 _13941_ (.A(_08037_),
    .B(net670),
    .Y(_08663_));
 sky130_fd_sc_hd__o211a_1 _13942_ (.A1(\core.csr.instruction_memoryAddress[28] ),
    .A2(net670),
    .B1(_08663_),
    .C1(net1894),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _13943_ (.A0(\core.csr.instruction_memoryAddress[29] ),
    .A1(_08053_),
    .S(net674),
    .X(_08664_));
 sky130_fd_sc_hd__and2_1 _13944_ (.A(net1891),
    .B(_08664_),
    .X(_00062_));
 sky130_fd_sc_hd__o22a_1 _13945_ (.A1(\core.csr.instruction_memoryAddress[30] ),
    .A2(net670),
    .B1(net623),
    .B2(_08024_),
    .X(_00063_));
 sky130_fd_sc_hd__o22a_1 _13946_ (.A1(\core.csr.instruction_memoryAddress[31] ),
    .A2(net670),
    .B1(net623),
    .B2(_08012_),
    .X(_00064_));
 sky130_fd_sc_hd__o21ba_1 _13947_ (.A1(\core.pipe0_fetch.currentPipeStall ),
    .A2(_08650_),
    .B1_N(_08654_),
    .X(_00065_));
 sky130_fd_sc_hd__o32a_1 _13948_ (.A1(net1672),
    .A2(net1655),
    .A3(_06151_),
    .B1(net1362),
    .B2(\coreWBInterface.readDataBuffered[0] ),
    .X(_08665_));
 sky130_fd_sc_hd__mux2_1 _13949_ (.A0(\core.pipe0_fetch.cachedInstruction[0] ),
    .A1(_08665_),
    .S(net1753),
    .X(_08666_));
 sky130_fd_sc_hd__o221a_1 _13950_ (.A1(\core.pipe0_currentInstruction[0] ),
    .A2(net682),
    .B1(net628),
    .B2(_08666_),
    .C1(net1926),
    .X(_00066_));
 sky130_fd_sc_hd__o32a_1 _13951_ (.A1(_04431_),
    .A2(net1655),
    .A3(_06054_),
    .B1(_08636_),
    .B2(\coreWBInterface.readDataBuffered[1] ),
    .X(_08667_));
 sky130_fd_sc_hd__mux2_1 _13952_ (.A0(\core.pipe0_fetch.cachedInstruction[1] ),
    .A1(_08667_),
    .S(net1753),
    .X(_08668_));
 sky130_fd_sc_hd__o221a_1 _13953_ (.A1(\core.pipe0_currentInstruction[1] ),
    .A2(net682),
    .B1(net628),
    .B2(_08668_),
    .C1(net1920),
    .X(_00067_));
 sky130_fd_sc_hd__o32a_1 _13954_ (.A1(net1672),
    .A2(net1655),
    .A3(_05972_),
    .B1(net1362),
    .B2(\coreWBInterface.readDataBuffered[2] ),
    .X(_08669_));
 sky130_fd_sc_hd__mux2_1 _13955_ (.A0(\core.pipe0_fetch.cachedInstruction[2] ),
    .A1(_08669_),
    .S(net1753),
    .X(_08670_));
 sky130_fd_sc_hd__o221a_1 _13956_ (.A1(\core.pipe0_currentInstruction[2] ),
    .A2(net684),
    .B1(net628),
    .B2(_08670_),
    .C1(net1928),
    .X(_00068_));
 sky130_fd_sc_hd__o32a_1 _13957_ (.A1(net1670),
    .A2(net1656),
    .A3(_05887_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[3] ),
    .X(_08671_));
 sky130_fd_sc_hd__mux2_1 _13958_ (.A0(\core.pipe0_fetch.cachedInstruction[3] ),
    .A1(_08671_),
    .S(net1753),
    .X(_08672_));
 sky130_fd_sc_hd__o221a_1 _13959_ (.A1(\core.pipe0_currentInstruction[3] ),
    .A2(net686),
    .B1(net627),
    .B2(_08672_),
    .C1(net1942),
    .X(_00069_));
 sky130_fd_sc_hd__o32a_1 _13960_ (.A1(net1670),
    .A2(net1655),
    .A3(_05803_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[4] ),
    .X(_08673_));
 sky130_fd_sc_hd__mux2_1 _13961_ (.A0(\core.pipe0_fetch.cachedInstruction[4] ),
    .A1(_08673_),
    .S(net1756),
    .X(_08674_));
 sky130_fd_sc_hd__o221a_1 _13962_ (.A1(\core.pipe0_currentInstruction[4] ),
    .A2(net686),
    .B1(net627),
    .B2(_08674_),
    .C1(net1943),
    .X(_00070_));
 sky130_fd_sc_hd__o32a_1 _13963_ (.A1(net1670),
    .A2(net1656),
    .A3(_05722_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[5] ),
    .X(_08675_));
 sky130_fd_sc_hd__mux2_1 _13964_ (.A0(\core.pipe0_fetch.cachedInstruction[5] ),
    .A1(_08675_),
    .S(net1756),
    .X(_08676_));
 sky130_fd_sc_hd__o221a_1 _13965_ (.A1(\core.pipe0_currentInstruction[5] ),
    .A2(net686),
    .B1(net627),
    .B2(_08676_),
    .C1(net1942),
    .X(_00071_));
 sky130_fd_sc_hd__o32a_1 _13966_ (.A1(net1672),
    .A2(net1656),
    .A3(_05637_),
    .B1(net1362),
    .B2(\coreWBInterface.readDataBuffered[6] ),
    .X(_08677_));
 sky130_fd_sc_hd__mux2_1 _13967_ (.A0(\core.pipe0_fetch.cachedInstruction[6] ),
    .A1(_08677_),
    .S(_04413_),
    .X(_08678_));
 sky130_fd_sc_hd__o221a_1 _13968_ (.A1(\core.pipe0_currentInstruction[6] ),
    .A2(net686),
    .B1(net627),
    .B2(_08678_),
    .C1(net1942),
    .X(_00072_));
 sky130_fd_sc_hd__o32a_1 _13969_ (.A1(net1669),
    .A2(net1656),
    .A3(_04569_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[7] ),
    .X(_08679_));
 sky130_fd_sc_hd__mux2_2 _13970_ (.A0(\core.pipe0_fetch.cachedInstruction[7] ),
    .A1(_08679_),
    .S(net1756),
    .X(_08680_));
 sky130_fd_sc_hd__o221a_1 _13971_ (.A1(\core.pipe0_currentInstruction[7] ),
    .A2(net681),
    .B1(net628),
    .B2(_08680_),
    .C1(net1924),
    .X(_00073_));
 sky130_fd_sc_hd__o32a_1 _13972_ (.A1(net1672),
    .A2(net1654),
    .A3(_06144_),
    .B1(net1362),
    .B2(\coreWBInterface.readDataBuffered[8] ),
    .X(_08681_));
 sky130_fd_sc_hd__mux2_1 _13973_ (.A0(\core.pipe0_fetch.cachedInstruction[8] ),
    .A1(_08681_),
    .S(net1753),
    .X(_08682_));
 sky130_fd_sc_hd__o221a_1 _13974_ (.A1(\core.pipe0_currentInstruction[8] ),
    .A2(net685),
    .B1(net628),
    .B2(_08682_),
    .C1(net1925),
    .X(_00074_));
 sky130_fd_sc_hd__o32a_1 _13975_ (.A1(net1672),
    .A2(net1654),
    .A3(_05458_),
    .B1(net1362),
    .B2(\coreWBInterface.readDataBuffered[9] ),
    .X(_08683_));
 sky130_fd_sc_hd__mux2_1 _13976_ (.A0(\core.pipe0_fetch.cachedInstruction[9] ),
    .A1(_08683_),
    .S(net1753),
    .X(_08684_));
 sky130_fd_sc_hd__o221a_1 _13977_ (.A1(\core.pipe0_currentInstruction[9] ),
    .A2(net681),
    .B1(net628),
    .B2(_08684_),
    .C1(net1923),
    .X(_00075_));
 sky130_fd_sc_hd__o32a_2 _13978_ (.A1(net1672),
    .A2(net1654),
    .A3(_05371_),
    .B1(net1362),
    .B2(\coreWBInterface.readDataBuffered[10] ),
    .X(_08685_));
 sky130_fd_sc_hd__mux2_1 _13979_ (.A0(\core.pipe0_fetch.cachedInstruction[10] ),
    .A1(_08685_),
    .S(net1753),
    .X(_08686_));
 sky130_fd_sc_hd__o221a_1 _13980_ (.A1(\core.pipe0_currentInstruction[10] ),
    .A2(net681),
    .B1(net628),
    .B2(_08686_),
    .C1(net1920),
    .X(_00076_));
 sky130_fd_sc_hd__o32a_1 _13981_ (.A1(net1669),
    .A2(net1653),
    .A3(_05283_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[11] ),
    .X(_08687_));
 sky130_fd_sc_hd__mux2_1 _13982_ (.A0(\core.pipe0_fetch.cachedInstruction[11] ),
    .A1(_08687_),
    .S(net1756),
    .X(_08688_));
 sky130_fd_sc_hd__o221a_1 _13983_ (.A1(\core.pipe0_currentInstruction[11] ),
    .A2(net685),
    .B1(net628),
    .B2(_08688_),
    .C1(net1929),
    .X(_00077_));
 sky130_fd_sc_hd__o32a_1 _13984_ (.A1(net1672),
    .A2(net1653),
    .A3(_04938_),
    .B1(net1362),
    .B2(\coreWBInterface.readDataBuffered[12] ),
    .X(_08689_));
 sky130_fd_sc_hd__mux2_1 _13985_ (.A0(\core.pipe0_fetch.cachedInstruction[12] ),
    .A1(_08689_),
    .S(net1753),
    .X(_08690_));
 sky130_fd_sc_hd__o221a_1 _13986_ (.A1(net1882),
    .A2(net685),
    .B1(net628),
    .B2(_08690_),
    .C1(net1925),
    .X(_00078_));
 sky130_fd_sc_hd__o32a_1 _13987_ (.A1(net1669),
    .A2(net1653),
    .A3(_05028_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[13] ),
    .X(_08691_));
 sky130_fd_sc_hd__mux2_1 _13988_ (.A0(\core.pipe0_fetch.cachedInstruction[13] ),
    .A1(_08691_),
    .S(net1754),
    .X(_08692_));
 sky130_fd_sc_hd__o221a_1 _13989_ (.A1(\core.pipe0_currentInstruction[13] ),
    .A2(net689),
    .B1(net625),
    .B2(_08692_),
    .C1(net1947),
    .X(_00079_));
 sky130_fd_sc_hd__o32a_1 _13990_ (.A1(net1670),
    .A2(net1653),
    .A3(_05194_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[14] ),
    .X(_08693_));
 sky130_fd_sc_hd__mux2_1 _13991_ (.A0(\core.pipe0_fetch.cachedInstruction[14] ),
    .A1(_08693_),
    .S(net1755),
    .X(_08694_));
 sky130_fd_sc_hd__o221a_1 _13992_ (.A1(\core.pipe0_currentInstruction[14] ),
    .A2(net687),
    .B1(net626),
    .B2(_08694_),
    .C1(net1944),
    .X(_00080_));
 sky130_fd_sc_hd__o32a_1 _13993_ (.A1(net1670),
    .A2(net1653),
    .A3(_04576_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[15] ),
    .X(_08695_));
 sky130_fd_sc_hd__mux2_1 _13994_ (.A0(\core.pipe0_fetch.cachedInstruction[15] ),
    .A1(_08695_),
    .S(net1756),
    .X(_08696_));
 sky130_fd_sc_hd__o221a_1 _13995_ (.A1(\core.pipe0_currentInstruction[15] ),
    .A2(net686),
    .B1(net627),
    .B2(_08696_),
    .C1(net1944),
    .X(_00081_));
 sky130_fd_sc_hd__o32a_1 _13996_ (.A1(net1669),
    .A2(net1651),
    .A3(_06154_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[16] ),
    .X(_08697_));
 sky130_fd_sc_hd__mux2_1 _13997_ (.A0(\core.pipe0_fetch.cachedInstruction[16] ),
    .A1(_08697_),
    .S(net1754),
    .X(_08698_));
 sky130_fd_sc_hd__o221a_1 _13998_ (.A1(net1877),
    .A2(net689),
    .B1(net625),
    .B2(_08698_),
    .C1(net1947),
    .X(_00082_));
 sky130_fd_sc_hd__o32a_2 _13999_ (.A1(net1669),
    .A2(net1651),
    .A3(_05463_),
    .B1(net1361),
    .B2(\coreWBInterface.readDataBuffered[17] ),
    .X(_08699_));
 sky130_fd_sc_hd__mux2_1 _14000_ (.A0(\core.pipe0_fetch.cachedInstruction[17] ),
    .A1(_08699_),
    .S(net1754),
    .X(_08700_));
 sky130_fd_sc_hd__o221a_1 _14001_ (.A1(net1866),
    .A2(net687),
    .B1(net625),
    .B2(_08700_),
    .C1(net1947),
    .X(_00083_));
 sky130_fd_sc_hd__o32a_1 _14002_ (.A1(net1672),
    .A2(_04583_),
    .A3(_05375_),
    .B1(net1362),
    .B2(\coreWBInterface.readDataBuffered[18] ),
    .X(_08701_));
 sky130_fd_sc_hd__mux2_1 _14003_ (.A0(\core.pipe0_fetch.cachedInstruction[18] ),
    .A1(_08701_),
    .S(net1753),
    .X(_08702_));
 sky130_fd_sc_hd__o221a_1 _14004_ (.A1(\core.pipe0_currentInstruction[18] ),
    .A2(net681),
    .B1(net628),
    .B2(_08702_),
    .C1(net1920),
    .X(_00084_));
 sky130_fd_sc_hd__o32a_2 _14005_ (.A1(net1669),
    .A2(net1651),
    .A3(_05287_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[19] ),
    .X(_08703_));
 sky130_fd_sc_hd__mux2_1 _14006_ (.A0(\core.pipe0_fetch.cachedInstruction[19] ),
    .A1(_08703_),
    .S(net1754),
    .X(_08704_));
 sky130_fd_sc_hd__o221a_1 _14007_ (.A1(net1860),
    .A2(net689),
    .B1(net625),
    .B2(_08704_),
    .C1(net1947),
    .X(_00085_));
 sky130_fd_sc_hd__o32a_1 _14008_ (.A1(net1671),
    .A2(net1652),
    .A3(_04856_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[20] ),
    .X(_08705_));
 sky130_fd_sc_hd__mux2_1 _14009_ (.A0(\core.pipe0_fetch.cachedInstruction[20] ),
    .A1(_08705_),
    .S(net1754),
    .X(_08706_));
 sky130_fd_sc_hd__o221a_1 _14010_ (.A1(net1851),
    .A2(net687),
    .B1(net626),
    .B2(_08706_),
    .C1(net1949),
    .X(_00086_));
 sky130_fd_sc_hd__o32a_1 _14011_ (.A1(net1669),
    .A2(net1651),
    .A3(_04779_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[21] ),
    .X(_08707_));
 sky130_fd_sc_hd__mux2_1 _14012_ (.A0(\core.pipe0_fetch.cachedInstruction[21] ),
    .A1(_08707_),
    .S(net1754),
    .X(_08708_));
 sky130_fd_sc_hd__o221a_1 _14013_ (.A1(net1849),
    .A2(net689),
    .B1(net625),
    .B2(_08708_),
    .C1(net1947),
    .X(_00087_));
 sky130_fd_sc_hd__o32a_1 _14014_ (.A1(net1670),
    .A2(net1652),
    .A3(_04699_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[22] ),
    .X(_08709_));
 sky130_fd_sc_hd__mux2_1 _14015_ (.A0(\core.pipe0_fetch.cachedInstruction[22] ),
    .A1(_08709_),
    .S(net1755),
    .X(_08710_));
 sky130_fd_sc_hd__o221a_1 _14016_ (.A1(net1837),
    .A2(net687),
    .B1(net626),
    .B2(_08710_),
    .C1(net1949),
    .X(_00088_));
 sky130_fd_sc_hd__o32a_1 _14017_ (.A1(net1670),
    .A2(net1652),
    .A3(_04584_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[23] ),
    .X(_08711_));
 sky130_fd_sc_hd__mux2_1 _14018_ (.A0(\core.pipe0_fetch.cachedInstruction[23] ),
    .A1(_08711_),
    .S(net1755),
    .X(_08712_));
 sky130_fd_sc_hd__o221a_1 _14019_ (.A1(net1831),
    .A2(net687),
    .B1(net626),
    .B2(_08712_),
    .C1(net1949),
    .X(_00089_));
 sky130_fd_sc_hd__o32a_1 _14020_ (.A1(net1669),
    .A2(net1660),
    .A3(_06140_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[24] ),
    .X(_08713_));
 sky130_fd_sc_hd__mux2_1 _14021_ (.A0(\core.pipe0_fetch.cachedInstruction[24] ),
    .A1(_08713_),
    .S(net1754),
    .X(_08714_));
 sky130_fd_sc_hd__o221a_1 _14022_ (.A1(net1828),
    .A2(net687),
    .B1(net625),
    .B2(_08714_),
    .C1(net1948),
    .X(_00090_));
 sky130_fd_sc_hd__o32a_1 _14023_ (.A1(net1671),
    .A2(net1660),
    .A3(_05468_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[25] ),
    .X(_08715_));
 sky130_fd_sc_hd__mux2_1 _14024_ (.A0(\core.pipe0_fetch.cachedInstruction[25] ),
    .A1(_08715_),
    .S(net1756),
    .X(_08716_));
 sky130_fd_sc_hd__o221a_1 _14025_ (.A1(net1822),
    .A2(net689),
    .B1(net627),
    .B2(_08716_),
    .C1(net1939),
    .X(_00091_));
 sky130_fd_sc_hd__o32a_1 _14026_ (.A1(net1669),
    .A2(net1660),
    .A3(_05380_),
    .B1(net1361),
    .B2(\coreWBInterface.readDataBuffered[26] ),
    .X(_08717_));
 sky130_fd_sc_hd__mux2_1 _14027_ (.A0(\core.pipe0_fetch.cachedInstruction[26] ),
    .A1(_08717_),
    .S(net1754),
    .X(_08718_));
 sky130_fd_sc_hd__o221a_1 _14028_ (.A1(\core.pipe0_currentInstruction[26] ),
    .A2(net687),
    .B1(net625),
    .B2(_08718_),
    .C1(net1939),
    .X(_00092_));
 sky130_fd_sc_hd__o32a_1 _14029_ (.A1(net1671),
    .A2(net1660),
    .A3(_05292_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[27] ),
    .X(_08719_));
 sky130_fd_sc_hd__mux2_1 _14030_ (.A0(\core.pipe0_fetch.cachedInstruction[27] ),
    .A1(_08719_),
    .S(net1754),
    .X(_08720_));
 sky130_fd_sc_hd__o221a_1 _14031_ (.A1(\core.pipe0_currentInstruction[27] ),
    .A2(net689),
    .B1(net625),
    .B2(_08720_),
    .C1(net1939),
    .X(_00093_));
 sky130_fd_sc_hd__o32a_1 _14032_ (.A1(net1670),
    .A2(net1661),
    .A3(_04951_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[28] ),
    .X(_08721_));
 sky130_fd_sc_hd__mux2_1 _14033_ (.A0(\core.pipe0_fetch.cachedInstruction[28] ),
    .A1(_08721_),
    .S(net1755),
    .X(_08722_));
 sky130_fd_sc_hd__o221a_1 _14034_ (.A1(\core.pipe0_currentInstruction[28] ),
    .A2(net687),
    .B1(net626),
    .B2(_08722_),
    .C1(net1944),
    .X(_00094_));
 sky130_fd_sc_hd__o32a_1 _14035_ (.A1(net1669),
    .A2(net1661),
    .A3(_05034_),
    .B1(net1359),
    .B2(\coreWBInterface.readDataBuffered[29] ),
    .X(_08723_));
 sky130_fd_sc_hd__mux2_1 _14036_ (.A0(\core.pipe0_fetch.cachedInstruction[29] ),
    .A1(_08723_),
    .S(net1754),
    .X(_08724_));
 sky130_fd_sc_hd__o221a_1 _14037_ (.A1(\core.pipe0_currentInstruction[29] ),
    .A2(net687),
    .B1(net625),
    .B2(_08724_),
    .C1(net1948),
    .X(_00095_));
 sky130_fd_sc_hd__o32a_1 _14038_ (.A1(net1670),
    .A2(net1660),
    .A3(_05200_),
    .B1(net1361),
    .B2(\coreWBInterface.readDataBuffered[30] ),
    .X(_08725_));
 sky130_fd_sc_hd__mux2_1 _14039_ (.A0(\core.pipe0_fetch.cachedInstruction[30] ),
    .A1(_08725_),
    .S(net1755),
    .X(_08726_));
 sky130_fd_sc_hd__o221a_1 _14040_ (.A1(net1818),
    .A2(net688),
    .B1(net625),
    .B2(_08726_),
    .C1(net1949),
    .X(_00096_));
 sky130_fd_sc_hd__o32a_1 _14041_ (.A1(net1670),
    .A2(net1661),
    .A3(_04560_),
    .B1(net1360),
    .B2(\coreWBInterface.readDataBuffered[31] ),
    .X(_08727_));
 sky130_fd_sc_hd__mux2_1 _14042_ (.A0(\core.pipe0_fetch.cachedInstruction[31] ),
    .A1(_08727_),
    .S(net1756),
    .X(_08728_));
 sky130_fd_sc_hd__o221a_1 _14043_ (.A1(net1816),
    .A2(net687),
    .B1(net627),
    .B2(_08728_),
    .C1(net1944),
    .X(_00097_));
 sky130_fd_sc_hd__nor2_1 _14044_ (.A(net699),
    .B(net696),
    .Y(_08729_));
 sky130_fd_sc_hd__or3_1 _14045_ (.A(net701),
    .B(net697),
    .C(_08665_),
    .X(_08730_));
 sky130_fd_sc_hd__o211a_1 _14046_ (.A1(\core.pipe0_fetch.cachedInstruction[0] ),
    .A2(net669),
    .B1(_08730_),
    .C1(net1923),
    .X(_00098_));
 sky130_fd_sc_hd__or3_1 _14047_ (.A(net701),
    .B(net697),
    .C(_08667_),
    .X(_08731_));
 sky130_fd_sc_hd__o211a_1 _14048_ (.A1(\core.pipe0_fetch.cachedInstruction[1] ),
    .A2(net669),
    .B1(_08731_),
    .C1(net1923),
    .X(_00099_));
 sky130_fd_sc_hd__or3_1 _14049_ (.A(net701),
    .B(net696),
    .C(_08669_),
    .X(_08732_));
 sky130_fd_sc_hd__o211a_1 _14050_ (.A1(\core.pipe0_fetch.cachedInstruction[2] ),
    .A2(net669),
    .B1(_08732_),
    .C1(net1927),
    .X(_00100_));
 sky130_fd_sc_hd__or3_1 _14051_ (.A(net701),
    .B(net696),
    .C(_08671_),
    .X(_08733_));
 sky130_fd_sc_hd__o211a_1 _14052_ (.A1(\core.pipe0_fetch.cachedInstruction[3] ),
    .A2(net669),
    .B1(_08733_),
    .C1(net1942),
    .X(_00101_));
 sky130_fd_sc_hd__or3_1 _14053_ (.A(net700),
    .B(net694),
    .C(_08673_),
    .X(_08734_));
 sky130_fd_sc_hd__o211a_1 _14054_ (.A1(\core.pipe0_fetch.cachedInstruction[4] ),
    .A2(net668),
    .B1(_08734_),
    .C1(net1942),
    .X(_00102_));
 sky130_fd_sc_hd__or3_1 _14055_ (.A(net700),
    .B(net694),
    .C(_08675_),
    .X(_08735_));
 sky130_fd_sc_hd__o211a_1 _14056_ (.A1(\core.pipe0_fetch.cachedInstruction[5] ),
    .A2(net668),
    .B1(_08735_),
    .C1(net1943),
    .X(_00103_));
 sky130_fd_sc_hd__or3_1 _14057_ (.A(net700),
    .B(net696),
    .C(_08677_),
    .X(_08736_));
 sky130_fd_sc_hd__o211a_1 _14058_ (.A1(\core.pipe0_fetch.cachedInstruction[6] ),
    .A2(net668),
    .B1(_08736_),
    .C1(net1943),
    .X(_00104_));
 sky130_fd_sc_hd__or3_1 _14059_ (.A(net700),
    .B(net696),
    .C(_08679_),
    .X(_08737_));
 sky130_fd_sc_hd__o211a_1 _14060_ (.A1(\core.pipe0_fetch.cachedInstruction[7] ),
    .A2(net668),
    .B1(_08737_),
    .C1(net1940),
    .X(_00105_));
 sky130_fd_sc_hd__or3_1 _14061_ (.A(net701),
    .B(net696),
    .C(_08681_),
    .X(_08738_));
 sky130_fd_sc_hd__o211a_1 _14062_ (.A1(\core.pipe0_fetch.cachedInstruction[8] ),
    .A2(net669),
    .B1(_08738_),
    .C1(net1925),
    .X(_00106_));
 sky130_fd_sc_hd__or3_1 _14063_ (.A(net701),
    .B(net696),
    .C(_08683_),
    .X(_08739_));
 sky130_fd_sc_hd__o211a_1 _14064_ (.A1(\core.pipe0_fetch.cachedInstruction[9] ),
    .A2(net669),
    .B1(_08739_),
    .C1(net1923),
    .X(_00107_));
 sky130_fd_sc_hd__or3_1 _14065_ (.A(net701),
    .B(net697),
    .C(_08685_),
    .X(_08740_));
 sky130_fd_sc_hd__o211a_1 _14066_ (.A1(\core.pipe0_fetch.cachedInstruction[10] ),
    .A2(net669),
    .B1(_08740_),
    .C1(net1923),
    .X(_00108_));
 sky130_fd_sc_hd__or3_1 _14067_ (.A(net700),
    .B(net696),
    .C(_08687_),
    .X(_08741_));
 sky130_fd_sc_hd__o211a_1 _14068_ (.A1(\core.pipe0_fetch.cachedInstruction[11] ),
    .A2(net668),
    .B1(_08741_),
    .C1(net1940),
    .X(_00109_));
 sky130_fd_sc_hd__or3_1 _14069_ (.A(net701),
    .B(net696),
    .C(_08689_),
    .X(_08742_));
 sky130_fd_sc_hd__o211a_1 _14070_ (.A1(\core.pipe0_fetch.cachedInstruction[12] ),
    .A2(net669),
    .B1(_08742_),
    .C1(net1929),
    .X(_00110_));
 sky130_fd_sc_hd__or3_1 _14071_ (.A(net698),
    .B(net695),
    .C(_08691_),
    .X(_08743_));
 sky130_fd_sc_hd__o211a_1 _14072_ (.A1(\core.pipe0_fetch.cachedInstruction[13] ),
    .A2(net666),
    .B1(_08743_),
    .C1(net1947),
    .X(_00111_));
 sky130_fd_sc_hd__or3_1 _14073_ (.A(net698),
    .B(_08644_),
    .C(_08693_),
    .X(_08744_));
 sky130_fd_sc_hd__o211a_1 _14074_ (.A1(\core.pipe0_fetch.cachedInstruction[14] ),
    .A2(net667),
    .B1(_08744_),
    .C1(net1945),
    .X(_00112_));
 sky130_fd_sc_hd__or3_1 _14075_ (.A(net700),
    .B(net694),
    .C(_08695_),
    .X(_08745_));
 sky130_fd_sc_hd__o211a_1 _14076_ (.A1(\core.pipe0_fetch.cachedInstruction[15] ),
    .A2(net668),
    .B1(_08745_),
    .C1(net1944),
    .X(_00113_));
 sky130_fd_sc_hd__or3_1 _14077_ (.A(net698),
    .B(net695),
    .C(_08697_),
    .X(_08746_));
 sky130_fd_sc_hd__o211a_1 _14078_ (.A1(\core.pipe0_fetch.cachedInstruction[16] ),
    .A2(net666),
    .B1(_08746_),
    .C1(net1947),
    .X(_00114_));
 sky130_fd_sc_hd__or3_1 _14079_ (.A(net698),
    .B(net695),
    .C(_08699_),
    .X(_08747_));
 sky130_fd_sc_hd__o211a_1 _14080_ (.A1(\core.pipe0_fetch.cachedInstruction[17] ),
    .A2(net666),
    .B1(_08747_),
    .C1(net1947),
    .X(_00115_));
 sky130_fd_sc_hd__or3_1 _14081_ (.A(net701),
    .B(net697),
    .C(_08701_),
    .X(_08748_));
 sky130_fd_sc_hd__o211a_1 _14082_ (.A1(\core.pipe0_fetch.cachedInstruction[18] ),
    .A2(net669),
    .B1(_08748_),
    .C1(net1923),
    .X(_00116_));
 sky130_fd_sc_hd__or3_1 _14083_ (.A(net698),
    .B(net695),
    .C(_08703_),
    .X(_08749_));
 sky130_fd_sc_hd__o211a_1 _14084_ (.A1(\core.pipe0_fetch.cachedInstruction[19] ),
    .A2(net666),
    .B1(_08749_),
    .C1(net1947),
    .X(_00117_));
 sky130_fd_sc_hd__or3_1 _14085_ (.A(net698),
    .B(net694),
    .C(_08705_),
    .X(_08750_));
 sky130_fd_sc_hd__o211a_1 _14086_ (.A1(\core.pipe0_fetch.cachedInstruction[20] ),
    .A2(net666),
    .B1(_08750_),
    .C1(net1949),
    .X(_00118_));
 sky130_fd_sc_hd__or3_1 _14087_ (.A(net698),
    .B(net695),
    .C(_08707_),
    .X(_08751_));
 sky130_fd_sc_hd__o211a_1 _14088_ (.A1(\core.pipe0_fetch.cachedInstruction[21] ),
    .A2(net666),
    .B1(_08751_),
    .C1(net1947),
    .X(_00119_));
 sky130_fd_sc_hd__or3_1 _14089_ (.A(net699),
    .B(net694),
    .C(_08709_),
    .X(_08752_));
 sky130_fd_sc_hd__o211a_1 _14090_ (.A1(\core.pipe0_fetch.cachedInstruction[22] ),
    .A2(net667),
    .B1(_08752_),
    .C1(net1949),
    .X(_00120_));
 sky130_fd_sc_hd__or3_1 _14091_ (.A(net699),
    .B(net694),
    .C(_08711_),
    .X(_08753_));
 sky130_fd_sc_hd__o211a_1 _14092_ (.A1(\core.pipe0_fetch.cachedInstruction[23] ),
    .A2(net666),
    .B1(_08753_),
    .C1(net1949),
    .X(_00121_));
 sky130_fd_sc_hd__or3_1 _14093_ (.A(net698),
    .B(net695),
    .C(_08713_),
    .X(_08754_));
 sky130_fd_sc_hd__o211a_1 _14094_ (.A1(\core.pipe0_fetch.cachedInstruction[24] ),
    .A2(net667),
    .B1(_08754_),
    .C1(net1948),
    .X(_00122_));
 sky130_fd_sc_hd__or3_1 _14095_ (.A(net700),
    .B(net695),
    .C(_08715_),
    .X(_08755_));
 sky130_fd_sc_hd__o211a_1 _14096_ (.A1(\core.pipe0_fetch.cachedInstruction[25] ),
    .A2(net668),
    .B1(_08755_),
    .C1(net1939),
    .X(_00123_));
 sky130_fd_sc_hd__or3_1 _14097_ (.A(net698),
    .B(net695),
    .C(_08717_),
    .X(_08756_));
 sky130_fd_sc_hd__o211a_1 _14098_ (.A1(\core.pipe0_fetch.cachedInstruction[26] ),
    .A2(net666),
    .B1(_08756_),
    .C1(net1941),
    .X(_00124_));
 sky130_fd_sc_hd__or3_1 _14099_ (.A(net698),
    .B(net695),
    .C(_08719_),
    .X(_08757_));
 sky130_fd_sc_hd__o211a_1 _14100_ (.A1(\core.pipe0_fetch.cachedInstruction[27] ),
    .A2(net666),
    .B1(_08757_),
    .C1(net1939),
    .X(_00125_));
 sky130_fd_sc_hd__or3_1 _14101_ (.A(net699),
    .B(net694),
    .C(_08721_),
    .X(_08758_));
 sky130_fd_sc_hd__o211a_1 _14102_ (.A1(\core.pipe0_fetch.cachedInstruction[28] ),
    .A2(net667),
    .B1(_08758_),
    .C1(net1944),
    .X(_00126_));
 sky130_fd_sc_hd__or3_1 _14103_ (.A(net699),
    .B(net694),
    .C(_08723_),
    .X(_08759_));
 sky130_fd_sc_hd__o211a_1 _14104_ (.A1(\core.pipe0_fetch.cachedInstruction[29] ),
    .A2(net666),
    .B1(_08759_),
    .C1(net1948),
    .X(_00127_));
 sky130_fd_sc_hd__or3_1 _14105_ (.A(net699),
    .B(net694),
    .C(_08725_),
    .X(_08760_));
 sky130_fd_sc_hd__o211a_1 _14106_ (.A1(\core.pipe0_fetch.cachedInstruction[30] ),
    .A2(net667),
    .B1(_08760_),
    .C1(net1949),
    .X(_00128_));
 sky130_fd_sc_hd__or3_1 _14107_ (.A(net700),
    .B(net694),
    .C(_08727_),
    .X(_08761_));
 sky130_fd_sc_hd__o211a_1 _14108_ (.A1(\core.pipe0_fetch.cachedInstruction[31] ),
    .A2(net668),
    .B1(_08761_),
    .C1(net1945),
    .X(_00129_));
 sky130_fd_sc_hd__a21oi_1 _14109_ (.A1(net1753),
    .A2(net701),
    .B1(_08650_),
    .Y(_00130_));
 sky130_fd_sc_hd__or3_2 _14110_ (.A(net782),
    .B(_07439_),
    .C(_07891_),
    .X(_08762_));
 sky130_fd_sc_hd__nand2_1 _14111_ (.A(net1928),
    .B(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__and3_1 _14112_ (.A(net1884),
    .B(net1668),
    .C(_07878_),
    .X(_08764_));
 sky130_fd_sc_hd__or4b_2 _14113_ (.A(net1775),
    .B(_07843_),
    .C(_07875_),
    .D_N(_08764_),
    .X(_08765_));
 sky130_fd_sc_hd__o21a_1 _14114_ (.A1(net1763),
    .A2(_08763_),
    .B1(_08765_),
    .X(_08766_));
 sky130_fd_sc_hd__a21oi_4 _14115_ (.A1(_08639_),
    .A2(_08643_),
    .B1(net1765),
    .Y(_08767_));
 sky130_fd_sc_hd__nor2_1 _14116_ (.A(net739),
    .B(net663),
    .Y(_08768_));
 sky130_fd_sc_hd__nor3_4 _14117_ (.A(net1370),
    .B(_07840_),
    .C(_07866_),
    .Y(_08769_));
 sky130_fd_sc_hd__a22o_4 _14118_ (.A1(\jtag.managementReadData[0] ),
    .A2(net1369),
    .B1(net1300),
    .B2(net215),
    .X(_08770_));
 sky130_fd_sc_hd__or2_2 _14119_ (.A(_07843_),
    .B(_07876_),
    .X(_08771_));
 sky130_fd_sc_hd__nor2_2 _14120_ (.A(_07875_),
    .B(_08771_),
    .Y(_08772_));
 sky130_fd_sc_hd__or2_4 _14121_ (.A(_07875_),
    .B(_08771_),
    .X(_08773_));
 sky130_fd_sc_hd__a21oi_1 _14122_ (.A1(net450),
    .A2(net951),
    .B1(_08770_),
    .Y(_08774_));
 sky130_fd_sc_hd__nand2_1 _14123_ (.A(net450),
    .B(_08770_),
    .Y(_08775_));
 sky130_fd_sc_hd__a31o_1 _14124_ (.A1(net450),
    .A2(_08770_),
    .A3(net951),
    .B1(net1774),
    .X(_08776_));
 sky130_fd_sc_hd__a2bb2o_1 _14125_ (.A1_N(_08774_),
    .A2_N(_08776_),
    .B1(net1774),
    .B2(_07442_),
    .X(_08777_));
 sky130_fd_sc_hd__or3_1 _14126_ (.A(net741),
    .B(net664),
    .C(_08777_),
    .X(_08778_));
 sky130_fd_sc_hd__o211a_1 _14127_ (.A1(\core.fetchProgramCounter[0] ),
    .A2(net622),
    .B1(_08778_),
    .C1(net1934),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_4 _14128_ (.A1(\jtag.managementReadData[1] ),
    .A2(net1370),
    .B1(net1300),
    .B2(net226),
    .X(_08779_));
 sky130_fd_sc_hd__and2_1 _14129_ (.A(net461),
    .B(_08779_),
    .X(_08780_));
 sky130_fd_sc_hd__xor2_4 _14130_ (.A(net461),
    .B(_08779_),
    .X(_08781_));
 sky130_fd_sc_hd__xnor2_1 _14131_ (.A(_08775_),
    .B(_08781_),
    .Y(_08782_));
 sky130_fd_sc_hd__mux2_1 _14132_ (.A0(_08779_),
    .A1(_08782_),
    .S(net951),
    .X(_08783_));
 sky130_fd_sc_hd__o21ba_1 _14133_ (.A1(net1775),
    .A2(_08783_),
    .B1_N(_07436_),
    .X(_08784_));
 sky130_fd_sc_hd__or3_1 _14134_ (.A(net740),
    .B(net665),
    .C(_08784_),
    .X(_08785_));
 sky130_fd_sc_hd__o211a_1 _14135_ (.A1(\core.fetchProgramCounter[1] ),
    .A2(net621),
    .B1(_08785_),
    .C1(net1934),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_4 _14136_ (.A1(\jtag.managementReadData[2] ),
    .A2(net1370),
    .B1(net1300),
    .B2(net237),
    .X(_08786_));
 sky130_fd_sc_hd__a31oi_4 _14137_ (.A1(net450),
    .A2(_08770_),
    .A3(_08781_),
    .B1(_08780_),
    .Y(_08787_));
 sky130_fd_sc_hd__nor2_1 _14138_ (.A(net472),
    .B(_08786_),
    .Y(_08788_));
 sky130_fd_sc_hd__nand2_1 _14139_ (.A(net472),
    .B(_08786_),
    .Y(_08789_));
 sky130_fd_sc_hd__and2b_1 _14140_ (.A_N(_08788_),
    .B(_08789_),
    .X(_08790_));
 sky130_fd_sc_hd__xnor2_1 _14141_ (.A(_08787_),
    .B(_08790_),
    .Y(_08791_));
 sky130_fd_sc_hd__mux2_1 _14142_ (.A0(_08786_),
    .A1(_08791_),
    .S(net951),
    .X(_08792_));
 sky130_fd_sc_hd__a21o_1 _14143_ (.A1(net1763),
    .A2(_08792_),
    .B1(_08391_),
    .X(_08793_));
 sky130_fd_sc_hd__or3_1 _14144_ (.A(net740),
    .B(net665),
    .C(_08793_),
    .X(_08794_));
 sky130_fd_sc_hd__o211a_1 _14145_ (.A1(\core.fetchProgramCounter[2] ),
    .A2(net621),
    .B1(_08794_),
    .C1(net1934),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_2 _14146_ (.A1(\jtag.managementReadData[3] ),
    .A2(net1370),
    .B1(net1300),
    .B2(net240),
    .X(_08795_));
 sky130_fd_sc_hd__nor2_1 _14147_ (.A(net475),
    .B(_08795_),
    .Y(_08796_));
 sky130_fd_sc_hd__and2_1 _14148_ (.A(net475),
    .B(_08795_),
    .X(_08797_));
 sky130_fd_sc_hd__or2_1 _14149_ (.A(_08796_),
    .B(_08797_),
    .X(_08798_));
 sky130_fd_sc_hd__o21ai_2 _14150_ (.A1(_08787_),
    .A2(_08788_),
    .B1(_08789_),
    .Y(_08799_));
 sky130_fd_sc_hd__xnor2_1 _14151_ (.A(_08798_),
    .B(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__mux2_1 _14152_ (.A0(_08795_),
    .A1(_08800_),
    .S(net951),
    .X(_08801_));
 sky130_fd_sc_hd__a21o_1 _14153_ (.A1(net1762),
    .A2(_08801_),
    .B1(_08406_),
    .X(_08802_));
 sky130_fd_sc_hd__or3_1 _14154_ (.A(net740),
    .B(net665),
    .C(_08802_),
    .X(_08803_));
 sky130_fd_sc_hd__o211a_1 _14155_ (.A1(\core.fetchProgramCounter[3] ),
    .A2(net621),
    .B1(_08803_),
    .C1(net1934),
    .X(_00134_));
 sky130_fd_sc_hd__a22o_4 _14156_ (.A1(\jtag.managementReadData[4] ),
    .A2(net1370),
    .B1(net1301),
    .B2(net241),
    .X(_08804_));
 sky130_fd_sc_hd__nor2_1 _14157_ (.A(net476),
    .B(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__nand2_1 _14158_ (.A(net476),
    .B(_08804_),
    .Y(_08806_));
 sky130_fd_sc_hd__and2b_1 _14159_ (.A_N(_08805_),
    .B(_08806_),
    .X(_08807_));
 sky130_fd_sc_hd__nor2_1 _14160_ (.A(_08797_),
    .B(_08799_),
    .Y(_08808_));
 sky130_fd_sc_hd__or2_2 _14161_ (.A(_08796_),
    .B(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__xnor2_1 _14162_ (.A(_08807_),
    .B(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__mux2_1 _14163_ (.A0(_08804_),
    .A1(_08810_),
    .S(net951),
    .X(_08811_));
 sky130_fd_sc_hd__a21o_1 _14164_ (.A1(net1762),
    .A2(_08811_),
    .B1(_08418_),
    .X(_08812_));
 sky130_fd_sc_hd__or3_1 _14165_ (.A(net740),
    .B(net665),
    .C(_08812_),
    .X(_08813_));
 sky130_fd_sc_hd__o211a_1 _14166_ (.A1(\core.fetchProgramCounter[4] ),
    .A2(net621),
    .B1(_08813_),
    .C1(net1934),
    .X(_00135_));
 sky130_fd_sc_hd__a22o_4 _14167_ (.A1(\jtag.managementReadData[5] ),
    .A2(net1369),
    .B1(net1300),
    .B2(net242),
    .X(_08814_));
 sky130_fd_sc_hd__xnor2_1 _14168_ (.A(net477),
    .B(_08814_),
    .Y(_08815_));
 sky130_fd_sc_hd__o21ai_2 _14169_ (.A1(_08805_),
    .A2(_08809_),
    .B1(_08806_),
    .Y(_08816_));
 sky130_fd_sc_hd__xnor2_1 _14170_ (.A(_08815_),
    .B(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__or2_1 _14171_ (.A(net952),
    .B(_08814_),
    .X(_08818_));
 sky130_fd_sc_hd__o211a_1 _14172_ (.A1(net956),
    .A2(_08817_),
    .B1(_08818_),
    .C1(net1762),
    .X(_08819_));
 sky130_fd_sc_hd__or3_1 _14173_ (.A(_08432_),
    .B(net740),
    .C(net664),
    .X(_08820_));
 sky130_fd_sc_hd__o221a_1 _14174_ (.A1(\core.fetchProgramCounter[5] ),
    .A2(net622),
    .B1(_08819_),
    .B2(_08820_),
    .C1(net1931),
    .X(_00136_));
 sky130_fd_sc_hd__a22o_4 _14175_ (.A1(\jtag.managementReadData[6] ),
    .A2(net1369),
    .B1(net1300),
    .B2(net243),
    .X(_08821_));
 sky130_fd_sc_hd__nor2_2 _14176_ (.A(net478),
    .B(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__nand2_2 _14177_ (.A(net478),
    .B(_08821_),
    .Y(_08823_));
 sky130_fd_sc_hd__nand2b_1 _14178_ (.A_N(_08822_),
    .B(_08823_),
    .Y(_08824_));
 sky130_fd_sc_hd__o21a_1 _14179_ (.A1(net477),
    .A2(_08814_),
    .B1(_08816_),
    .X(_08825_));
 sky130_fd_sc_hd__a21oi_4 _14180_ (.A1(net477),
    .A2(_08814_),
    .B1(_08825_),
    .Y(_08826_));
 sky130_fd_sc_hd__xnor2_1 _14181_ (.A(_08824_),
    .B(_08826_),
    .Y(_08827_));
 sky130_fd_sc_hd__nand2_1 _14182_ (.A(net951),
    .B(_08827_),
    .Y(_08828_));
 sky130_fd_sc_hd__o211a_1 _14183_ (.A1(net951),
    .A2(_08821_),
    .B1(_08828_),
    .C1(net1762),
    .X(_08829_));
 sky130_fd_sc_hd__or3_1 _14184_ (.A(_08448_),
    .B(net741),
    .C(net664),
    .X(_08830_));
 sky130_fd_sc_hd__o221a_1 _14185_ (.A1(\core.fetchProgramCounter[6] ),
    .A2(net621),
    .B1(_08829_),
    .B2(_08830_),
    .C1(net1938),
    .X(_00137_));
 sky130_fd_sc_hd__a22o_4 _14186_ (.A1(\jtag.managementReadData[7] ),
    .A2(net1369),
    .B1(net1300),
    .B2(net244),
    .X(_08831_));
 sky130_fd_sc_hd__or2_2 _14187_ (.A(net479),
    .B(_08831_),
    .X(_08832_));
 sky130_fd_sc_hd__nand2_1 _14188_ (.A(net479),
    .B(_08831_),
    .Y(_08833_));
 sky130_fd_sc_hd__nand2_1 _14189_ (.A(_08832_),
    .B(_08833_),
    .Y(_08834_));
 sky130_fd_sc_hd__o21ai_4 _14190_ (.A1(_08822_),
    .A2(_08826_),
    .B1(_08823_),
    .Y(_08835_));
 sky130_fd_sc_hd__xnor2_1 _14191_ (.A(_08834_),
    .B(_08835_),
    .Y(_08836_));
 sky130_fd_sc_hd__mux2_1 _14192_ (.A0(_08831_),
    .A1(_08836_),
    .S(net951),
    .X(_08837_));
 sky130_fd_sc_hd__a21bo_1 _14193_ (.A1(net1764),
    .A2(_08837_),
    .B1_N(_08460_),
    .X(_08838_));
 sky130_fd_sc_hd__or3_1 _14194_ (.A(net741),
    .B(net664),
    .C(_08838_),
    .X(_08839_));
 sky130_fd_sc_hd__o211a_1 _14195_ (.A1(\core.fetchProgramCounter[7] ),
    .A2(net622),
    .B1(_08839_),
    .C1(net1930),
    .X(_00138_));
 sky130_fd_sc_hd__a22o_4 _14196_ (.A1(\jtag.managementReadData[8] ),
    .A2(net1369),
    .B1(net1300),
    .B2(net245),
    .X(_08840_));
 sky130_fd_sc_hd__nor2_2 _14197_ (.A(net480),
    .B(_08840_),
    .Y(_08841_));
 sky130_fd_sc_hd__nand2_2 _14198_ (.A(net480),
    .B(_08840_),
    .Y(_08842_));
 sky130_fd_sc_hd__and2b_1 _14199_ (.A_N(_08841_),
    .B(_08842_),
    .X(_08843_));
 sky130_fd_sc_hd__a21boi_4 _14200_ (.A1(_08832_),
    .A2(_08835_),
    .B1_N(_08833_),
    .Y(_08844_));
 sky130_fd_sc_hd__xnor2_1 _14201_ (.A(_08843_),
    .B(_08844_),
    .Y(_08845_));
 sky130_fd_sc_hd__mux2_1 _14202_ (.A0(_08840_),
    .A1(_08845_),
    .S(net951),
    .X(_08846_));
 sky130_fd_sc_hd__a21bo_1 _14203_ (.A1(net1764),
    .A2(_08846_),
    .B1_N(_08475_),
    .X(_08847_));
 sky130_fd_sc_hd__or3_1 _14204_ (.A(net741),
    .B(net665),
    .C(_08847_),
    .X(_08848_));
 sky130_fd_sc_hd__o211a_1 _14205_ (.A1(\core.fetchProgramCounter[8] ),
    .A2(net622),
    .B1(_08848_),
    .C1(net1930),
    .X(_00139_));
 sky130_fd_sc_hd__a22o_4 _14206_ (.A1(\jtag.managementReadData[9] ),
    .A2(net1369),
    .B1(net1300),
    .B2(net246),
    .X(_08849_));
 sky130_fd_sc_hd__or2_1 _14207_ (.A(net481),
    .B(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__nand2_1 _14208_ (.A(net481),
    .B(_08849_),
    .Y(_08851_));
 sky130_fd_sc_hd__nand2_1 _14209_ (.A(_08850_),
    .B(_08851_),
    .Y(_08852_));
 sky130_fd_sc_hd__o21ai_4 _14210_ (.A1(_08841_),
    .A2(_08844_),
    .B1(_08842_),
    .Y(_08853_));
 sky130_fd_sc_hd__xnor2_1 _14211_ (.A(_08852_),
    .B(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__mux2_1 _14212_ (.A0(_08849_),
    .A1(_08854_),
    .S(net952),
    .X(_08855_));
 sky130_fd_sc_hd__a21o_1 _14213_ (.A1(net1765),
    .A2(_08855_),
    .B1(_08486_),
    .X(_08856_));
 sky130_fd_sc_hd__or3_1 _14214_ (.A(net740),
    .B(net664),
    .C(_08856_),
    .X(_08857_));
 sky130_fd_sc_hd__o211a_1 _14215_ (.A1(\core.fetchProgramCounter[9] ),
    .A2(net621),
    .B1(_08857_),
    .C1(net1913),
    .X(_00140_));
 sky130_fd_sc_hd__a22o_4 _14216_ (.A1(\jtag.managementReadData[10] ),
    .A2(net1370),
    .B1(net1300),
    .B2(net216),
    .X(_08858_));
 sky130_fd_sc_hd__nand2_1 _14217_ (.A(net451),
    .B(_08858_),
    .Y(_08859_));
 sky130_fd_sc_hd__or2_1 _14218_ (.A(net451),
    .B(_08858_),
    .X(_08860_));
 sky130_fd_sc_hd__nand2_1 _14219_ (.A(_08859_),
    .B(_08860_),
    .Y(_08861_));
 sky130_fd_sc_hd__a21bo_1 _14220_ (.A1(_08850_),
    .A2(_08853_),
    .B1_N(_08851_),
    .X(_08862_));
 sky130_fd_sc_hd__xnor2_1 _14221_ (.A(_08861_),
    .B(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__mux2_1 _14222_ (.A0(_08858_),
    .A1(_08863_),
    .S(net952),
    .X(_08864_));
 sky130_fd_sc_hd__o21a_1 _14223_ (.A1(net1773),
    .A2(_08864_),
    .B1(_08501_),
    .X(_08865_));
 sky130_fd_sc_hd__or3_1 _14224_ (.A(net740),
    .B(net664),
    .C(_08865_),
    .X(_08866_));
 sky130_fd_sc_hd__o211a_1 _14225_ (.A1(\core.fetchProgramCounter[10] ),
    .A2(net621),
    .B1(_08866_),
    .C1(net1913),
    .X(_00141_));
 sky130_fd_sc_hd__a21bo_1 _14226_ (.A1(_08860_),
    .A2(_08862_),
    .B1_N(_08859_),
    .X(_08867_));
 sky130_fd_sc_hd__a22o_4 _14227_ (.A1(\jtag.managementReadData[11] ),
    .A2(net1369),
    .B1(net1301),
    .B2(net217),
    .X(_08868_));
 sky130_fd_sc_hd__nand2_1 _14228_ (.A(net452),
    .B(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__or2_1 _14229_ (.A(net452),
    .B(_08868_),
    .X(_08870_));
 sky130_fd_sc_hd__and2_1 _14230_ (.A(_08869_),
    .B(_08870_),
    .X(_08871_));
 sky130_fd_sc_hd__nand2_1 _14231_ (.A(_08867_),
    .B(_08871_),
    .Y(_08872_));
 sky130_fd_sc_hd__xor2_1 _14232_ (.A(_08867_),
    .B(_08871_),
    .X(_08873_));
 sky130_fd_sc_hd__mux2_1 _14233_ (.A0(_08868_),
    .A1(_08873_),
    .S(net952),
    .X(_08874_));
 sky130_fd_sc_hd__o21ba_1 _14234_ (.A1(net1772),
    .A2(_08874_),
    .B1_N(_08365_),
    .X(_08875_));
 sky130_fd_sc_hd__or3_1 _14235_ (.A(net740),
    .B(net664),
    .C(_08875_),
    .X(_08876_));
 sky130_fd_sc_hd__o211a_1 _14236_ (.A1(\core.fetchProgramCounter[11] ),
    .A2(net621),
    .B1(_08876_),
    .C1(net1915),
    .X(_00142_));
 sky130_fd_sc_hd__a22o_4 _14237_ (.A1(\jtag.managementReadData[12] ),
    .A2(net1369),
    .B1(net1301),
    .B2(net218),
    .X(_08877_));
 sky130_fd_sc_hd__nand2_1 _14238_ (.A(net453),
    .B(_08877_),
    .Y(_08878_));
 sky130_fd_sc_hd__xnor2_1 _14239_ (.A(net453),
    .B(_08877_),
    .Y(_08879_));
 sky130_fd_sc_hd__and3_1 _14240_ (.A(_08869_),
    .B(_08872_),
    .C(_08879_),
    .X(_08880_));
 sky130_fd_sc_hd__a21o_1 _14241_ (.A1(_08869_),
    .A2(_08872_),
    .B1(_08879_),
    .X(_08881_));
 sky130_fd_sc_hd__or3b_1 _14242_ (.A(net956),
    .B(_08880_),
    .C_N(_08881_),
    .X(_08882_));
 sky130_fd_sc_hd__a21bo_1 _14243_ (.A1(net956),
    .A2(_08877_),
    .B1_N(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__o21a_1 _14244_ (.A1(net1772),
    .A2(_08883_),
    .B1(_08227_),
    .X(_08884_));
 sky130_fd_sc_hd__or3_1 _14245_ (.A(net740),
    .B(net664),
    .C(_08884_),
    .X(_08885_));
 sky130_fd_sc_hd__o211a_1 _14246_ (.A1(\core.fetchProgramCounter[12] ),
    .A2(net621),
    .B1(_08885_),
    .C1(net1915),
    .X(_00143_));
 sky130_fd_sc_hd__a22o_4 _14247_ (.A1(\jtag.managementReadData[13] ),
    .A2(net1371),
    .B1(net1301),
    .B2(net219),
    .X(_08886_));
 sky130_fd_sc_hd__nand2_1 _14248_ (.A(net454),
    .B(_08886_),
    .Y(_08887_));
 sky130_fd_sc_hd__xnor2_1 _14249_ (.A(net454),
    .B(_08886_),
    .Y(_08888_));
 sky130_fd_sc_hd__and3_1 _14250_ (.A(_08878_),
    .B(_08881_),
    .C(_08888_),
    .X(_08889_));
 sky130_fd_sc_hd__a21o_1 _14251_ (.A1(_08878_),
    .A2(_08881_),
    .B1(_08888_),
    .X(_08890_));
 sky130_fd_sc_hd__or3b_1 _14252_ (.A(net956),
    .B(_08889_),
    .C_N(_08890_),
    .X(_08891_));
 sky130_fd_sc_hd__a21bo_1 _14253_ (.A1(net956),
    .A2(_08886_),
    .B1_N(_08891_),
    .X(_08892_));
 sky130_fd_sc_hd__o21a_1 _14254_ (.A1(net1771),
    .A2(_08892_),
    .B1(_08202_),
    .X(_08893_));
 sky130_fd_sc_hd__or3_1 _14255_ (.A(net740),
    .B(net664),
    .C(_08893_),
    .X(_08894_));
 sky130_fd_sc_hd__o211a_1 _14256_ (.A1(\core.fetchProgramCounter[13] ),
    .A2(net621),
    .B1(_08894_),
    .C1(net1915),
    .X(_00144_));
 sky130_fd_sc_hd__a22o_4 _14257_ (.A1(\jtag.managementReadData[14] ),
    .A2(net1371),
    .B1(net1301),
    .B2(net220),
    .X(_08895_));
 sky130_fd_sc_hd__nand2_1 _14258_ (.A(net455),
    .B(_08895_),
    .Y(_08896_));
 sky130_fd_sc_hd__xnor2_1 _14259_ (.A(net455),
    .B(_08895_),
    .Y(_08897_));
 sky130_fd_sc_hd__and3_1 _14260_ (.A(_08887_),
    .B(_08890_),
    .C(_08897_),
    .X(_08898_));
 sky130_fd_sc_hd__a21o_1 _14261_ (.A1(_08887_),
    .A2(_08890_),
    .B1(_08897_),
    .X(_08899_));
 sky130_fd_sc_hd__or3b_1 _14262_ (.A(net956),
    .B(_08898_),
    .C_N(_08899_),
    .X(_08900_));
 sky130_fd_sc_hd__a21bo_1 _14263_ (.A1(net956),
    .A2(_08895_),
    .B1_N(_08900_),
    .X(_08901_));
 sky130_fd_sc_hd__o21a_1 _14264_ (.A1(net1771),
    .A2(_08901_),
    .B1(_08294_),
    .X(_08902_));
 sky130_fd_sc_hd__or3_1 _14265_ (.A(net739),
    .B(net663),
    .C(_08902_),
    .X(_08903_));
 sky130_fd_sc_hd__o211a_1 _14266_ (.A1(\core.fetchProgramCounter[14] ),
    .A2(net620),
    .B1(_08903_),
    .C1(net1910),
    .X(_00145_));
 sky130_fd_sc_hd__a22o_4 _14267_ (.A1(\jtag.managementReadData[15] ),
    .A2(net1371),
    .B1(net1301),
    .B2(net221),
    .X(_08904_));
 sky130_fd_sc_hd__and2_1 _14268_ (.A(net456),
    .B(_08904_),
    .X(_08905_));
 sky130_fd_sc_hd__nor2_1 _14269_ (.A(net456),
    .B(_08904_),
    .Y(_08906_));
 sky130_fd_sc_hd__or2_1 _14270_ (.A(_08905_),
    .B(_08906_),
    .X(_08907_));
 sky130_fd_sc_hd__and3_1 _14271_ (.A(_08896_),
    .B(_08899_),
    .C(_08907_),
    .X(_08908_));
 sky130_fd_sc_hd__a21oi_2 _14272_ (.A1(_08896_),
    .A2(_08899_),
    .B1(_08907_),
    .Y(_08909_));
 sky130_fd_sc_hd__nor2_1 _14273_ (.A(_08908_),
    .B(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__mux2_1 _14274_ (.A0(_08904_),
    .A1(_08910_),
    .S(net953),
    .X(_08911_));
 sky130_fd_sc_hd__o21a_1 _14275_ (.A1(net1771),
    .A2(_08911_),
    .B1(_08317_),
    .X(_08912_));
 sky130_fd_sc_hd__or3_1 _14276_ (.A(net739),
    .B(net663),
    .C(_08912_),
    .X(_08913_));
 sky130_fd_sc_hd__o211a_1 _14277_ (.A1(\core.fetchProgramCounter[15] ),
    .A2(net620),
    .B1(_08913_),
    .C1(net1910),
    .X(_00146_));
 sky130_fd_sc_hd__nor2_2 _14278_ (.A(_08905_),
    .B(_08909_),
    .Y(_08914_));
 sky130_fd_sc_hd__a22o_4 _14279_ (.A1(\jtag.managementReadData[16] ),
    .A2(net1368),
    .B1(net1299),
    .B2(net222),
    .X(_08915_));
 sky130_fd_sc_hd__nor2_1 _14280_ (.A(net457),
    .B(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__nand2_1 _14281_ (.A(net457),
    .B(_08915_),
    .Y(_08917_));
 sky130_fd_sc_hd__and2b_1 _14282_ (.A_N(_08916_),
    .B(_08917_),
    .X(_08918_));
 sky130_fd_sc_hd__xnor2_1 _14283_ (.A(_08914_),
    .B(_08918_),
    .Y(_08919_));
 sky130_fd_sc_hd__mux2_1 _14284_ (.A0(_08915_),
    .A1(_08919_),
    .S(net953),
    .X(_08920_));
 sky130_fd_sc_hd__o21ba_1 _14285_ (.A1(net1769),
    .A2(_08920_),
    .B1_N(_08265_),
    .X(_08921_));
 sky130_fd_sc_hd__or3_1 _14286_ (.A(net739),
    .B(net663),
    .C(_08921_),
    .X(_08922_));
 sky130_fd_sc_hd__o211a_1 _14287_ (.A1(\core.fetchProgramCounter[16] ),
    .A2(net620),
    .B1(_08922_),
    .C1(net1909),
    .X(_00147_));
 sky130_fd_sc_hd__a22o_4 _14288_ (.A1(\jtag.managementReadData[17] ),
    .A2(net1368),
    .B1(net1299),
    .B2(net223),
    .X(_08923_));
 sky130_fd_sc_hd__nor2_1 _14289_ (.A(net458),
    .B(_08923_),
    .Y(_08924_));
 sky130_fd_sc_hd__and2_1 _14290_ (.A(net458),
    .B(_08923_),
    .X(_08925_));
 sky130_fd_sc_hd__or2_1 _14291_ (.A(_08924_),
    .B(_08925_),
    .X(_08926_));
 sky130_fd_sc_hd__o21ai_2 _14292_ (.A1(_08914_),
    .A2(_08916_),
    .B1(_08917_),
    .Y(_08927_));
 sky130_fd_sc_hd__xnor2_1 _14293_ (.A(_08926_),
    .B(_08927_),
    .Y(_08928_));
 sky130_fd_sc_hd__or2_1 _14294_ (.A(net953),
    .B(_08923_),
    .X(_08929_));
 sky130_fd_sc_hd__o211a_1 _14295_ (.A1(net955),
    .A2(_08928_),
    .B1(_08929_),
    .C1(net1761),
    .X(_08930_));
 sky130_fd_sc_hd__or3_1 _14296_ (.A(_08252_),
    .B(net739),
    .C(net663),
    .X(_08931_));
 sky130_fd_sc_hd__o221a_1 _14297_ (.A1(\core.fetchProgramCounter[17] ),
    .A2(net620),
    .B1(_08930_),
    .B2(_08931_),
    .C1(net1909),
    .X(_00148_));
 sky130_fd_sc_hd__a22o_4 _14298_ (.A1(\jtag.managementReadData[18] ),
    .A2(net1368),
    .B1(net1299),
    .B2(net224),
    .X(_08932_));
 sky130_fd_sc_hd__nand2_1 _14299_ (.A(net459),
    .B(_08932_),
    .Y(_08933_));
 sky130_fd_sc_hd__or2_1 _14300_ (.A(net459),
    .B(_08932_),
    .X(_08934_));
 sky130_fd_sc_hd__nand2_1 _14301_ (.A(_08933_),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__nor2_1 _14302_ (.A(_08925_),
    .B(_08927_),
    .Y(_08936_));
 sky130_fd_sc_hd__nor2_1 _14303_ (.A(_08924_),
    .B(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__xnor2_1 _14304_ (.A(_08935_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__mux2_1 _14305_ (.A0(_08932_),
    .A1(_08938_),
    .S(net953),
    .X(_08939_));
 sky130_fd_sc_hd__o21a_1 _14306_ (.A1(net1769),
    .A2(_08939_),
    .B1(_08238_),
    .X(_08940_));
 sky130_fd_sc_hd__or3_1 _14307_ (.A(net739),
    .B(net663),
    .C(_08940_),
    .X(_08941_));
 sky130_fd_sc_hd__o211a_1 _14308_ (.A1(\core.fetchProgramCounter[18] ),
    .A2(net620),
    .B1(_08941_),
    .C1(net1909),
    .X(_00149_));
 sky130_fd_sc_hd__a21boi_1 _14309_ (.A1(_08934_),
    .A2(_08937_),
    .B1_N(_08933_),
    .Y(_08942_));
 sky130_fd_sc_hd__a22o_4 _14310_ (.A1(\jtag.managementReadData[19] ),
    .A2(net1368),
    .B1(net1299),
    .B2(net225),
    .X(_08943_));
 sky130_fd_sc_hd__nand2_1 _14311_ (.A(net460),
    .B(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__xnor2_1 _14312_ (.A(net460),
    .B(_08943_),
    .Y(_08945_));
 sky130_fd_sc_hd__and2_1 _14313_ (.A(_08942_),
    .B(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__or2_1 _14314_ (.A(_08942_),
    .B(_08945_),
    .X(_08947_));
 sky130_fd_sc_hd__or3b_1 _14315_ (.A(net955),
    .B(_08946_),
    .C_N(_08947_),
    .X(_08948_));
 sky130_fd_sc_hd__a21bo_1 _14316_ (.A1(net955),
    .A2(_08943_),
    .B1_N(_08948_),
    .X(_08949_));
 sky130_fd_sc_hd__o21a_1 _14317_ (.A1(net1768),
    .A2(_08949_),
    .B1(_08215_),
    .X(_08950_));
 sky130_fd_sc_hd__or3_1 _14318_ (.A(net739),
    .B(net663),
    .C(_08950_),
    .X(_08951_));
 sky130_fd_sc_hd__o211a_1 _14319_ (.A1(\core.fetchProgramCounter[19] ),
    .A2(net620),
    .B1(_08951_),
    .C1(net1909),
    .X(_00150_));
 sky130_fd_sc_hd__a22o_4 _14320_ (.A1(\jtag.managementReadData[20] ),
    .A2(net1368),
    .B1(net1299),
    .B2(net227),
    .X(_08952_));
 sky130_fd_sc_hd__nand2_1 _14321_ (.A(net462),
    .B(_08952_),
    .Y(_08953_));
 sky130_fd_sc_hd__xnor2_1 _14322_ (.A(net462),
    .B(_08952_),
    .Y(_08954_));
 sky130_fd_sc_hd__and3_1 _14323_ (.A(_08944_),
    .B(_08947_),
    .C(_08954_),
    .X(_08955_));
 sky130_fd_sc_hd__a21o_1 _14324_ (.A1(_08944_),
    .A2(_08947_),
    .B1(_08954_),
    .X(_08956_));
 sky130_fd_sc_hd__or3b_1 _14325_ (.A(net955),
    .B(_08955_),
    .C_N(_08956_),
    .X(_08957_));
 sky130_fd_sc_hd__a21bo_1 _14326_ (.A1(net955),
    .A2(_08952_),
    .B1_N(_08957_),
    .X(_08958_));
 sky130_fd_sc_hd__o21a_1 _14327_ (.A1(net1768),
    .A2(_08958_),
    .B1(_08281_),
    .X(_08959_));
 sky130_fd_sc_hd__or3_1 _14328_ (.A(net739),
    .B(net662),
    .C(_08959_),
    .X(_08960_));
 sky130_fd_sc_hd__o211a_1 _14329_ (.A1(\core.fetchProgramCounter[20] ),
    .A2(net619),
    .B1(_08960_),
    .C1(net1900),
    .X(_00151_));
 sky130_fd_sc_hd__a22o_4 _14330_ (.A1(\jtag.managementReadData[21] ),
    .A2(net1368),
    .B1(net1299),
    .B2(net228),
    .X(_08961_));
 sky130_fd_sc_hd__nand2_1 _14331_ (.A(net463),
    .B(_08961_),
    .Y(_08962_));
 sky130_fd_sc_hd__xnor2_1 _14332_ (.A(net463),
    .B(_08961_),
    .Y(_08963_));
 sky130_fd_sc_hd__and3_1 _14333_ (.A(_08953_),
    .B(_08956_),
    .C(_08963_),
    .X(_08964_));
 sky130_fd_sc_hd__a21o_1 _14334_ (.A1(_08953_),
    .A2(_08956_),
    .B1(_08963_),
    .X(_08965_));
 sky130_fd_sc_hd__or3b_1 _14335_ (.A(net954),
    .B(_08964_),
    .C_N(_08965_),
    .X(_08966_));
 sky130_fd_sc_hd__a21bo_1 _14336_ (.A1(net954),
    .A2(_08961_),
    .B1_N(_08966_),
    .X(_08967_));
 sky130_fd_sc_hd__o21a_1 _14337_ (.A1(net1767),
    .A2(_08967_),
    .B1(_08182_),
    .X(_08968_));
 sky130_fd_sc_hd__or3_1 _14338_ (.A(net738),
    .B(net662),
    .C(_08968_),
    .X(_08969_));
 sky130_fd_sc_hd__o211a_1 _14339_ (.A1(\core.fetchProgramCounter[21] ),
    .A2(net619),
    .B1(_08969_),
    .C1(net1899),
    .X(_00152_));
 sky130_fd_sc_hd__a22o_4 _14340_ (.A1(\jtag.managementReadData[22] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net229),
    .X(_08970_));
 sky130_fd_sc_hd__nand2_1 _14341_ (.A(net464),
    .B(_08970_),
    .Y(_08971_));
 sky130_fd_sc_hd__xnor2_1 _14342_ (.A(net464),
    .B(_08970_),
    .Y(_08972_));
 sky130_fd_sc_hd__and3_1 _14343_ (.A(_08962_),
    .B(_08965_),
    .C(_08972_),
    .X(_08973_));
 sky130_fd_sc_hd__a21o_1 _14344_ (.A1(_08962_),
    .A2(_08965_),
    .B1(_08972_),
    .X(_08974_));
 sky130_fd_sc_hd__or3b_1 _14345_ (.A(net954),
    .B(_08973_),
    .C_N(_08974_),
    .X(_08975_));
 sky130_fd_sc_hd__a21bo_1 _14346_ (.A1(net954),
    .A2(_08970_),
    .B1_N(_08975_),
    .X(_08976_));
 sky130_fd_sc_hd__o21a_1 _14347_ (.A1(net1766),
    .A2(_08976_),
    .B1(_08307_),
    .X(_08977_));
 sky130_fd_sc_hd__or3_1 _14348_ (.A(net738),
    .B(net662),
    .C(_08977_),
    .X(_08978_));
 sky130_fd_sc_hd__o211a_1 _14349_ (.A1(\core.fetchProgramCounter[22] ),
    .A2(net619),
    .B1(_08978_),
    .C1(net1888),
    .X(_00153_));
 sky130_fd_sc_hd__a22o_2 _14350_ (.A1(\jtag.managementReadData[23] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net230),
    .X(_08979_));
 sky130_fd_sc_hd__and2_1 _14351_ (.A(net465),
    .B(_08979_),
    .X(_08980_));
 sky130_fd_sc_hd__nor2_1 _14352_ (.A(net465),
    .B(_08979_),
    .Y(_08981_));
 sky130_fd_sc_hd__or2_1 _14353_ (.A(_08980_),
    .B(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__and3_1 _14354_ (.A(_08971_),
    .B(_08974_),
    .C(_08982_),
    .X(_08983_));
 sky130_fd_sc_hd__a21oi_1 _14355_ (.A1(_08971_),
    .A2(_08974_),
    .B1(_08982_),
    .Y(_08984_));
 sky130_fd_sc_hd__nor2_1 _14356_ (.A(_08983_),
    .B(_08984_),
    .Y(_08985_));
 sky130_fd_sc_hd__mux2_1 _14357_ (.A0(_08979_),
    .A1(_08985_),
    .S(net953),
    .X(_08986_));
 sky130_fd_sc_hd__o21a_1 _14358_ (.A1(net1766),
    .A2(_08986_),
    .B1(_08170_),
    .X(_08987_));
 sky130_fd_sc_hd__or3_1 _14359_ (.A(net738),
    .B(net662),
    .C(_08987_),
    .X(_08988_));
 sky130_fd_sc_hd__o211a_1 _14360_ (.A1(\core.fetchProgramCounter[23] ),
    .A2(net619),
    .B1(_08988_),
    .C1(net1894),
    .X(_00154_));
 sky130_fd_sc_hd__nor2_1 _14361_ (.A(_08980_),
    .B(_08984_),
    .Y(_08989_));
 sky130_fd_sc_hd__a22o_2 _14362_ (.A1(\jtag.managementReadData[24] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net231),
    .X(_08990_));
 sky130_fd_sc_hd__nor2_1 _14363_ (.A(net466),
    .B(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__nand2_1 _14364_ (.A(net466),
    .B(_08990_),
    .Y(_08992_));
 sky130_fd_sc_hd__nand2b_1 _14365_ (.A_N(_08991_),
    .B(_08992_),
    .Y(_08993_));
 sky130_fd_sc_hd__xnor2_1 _14366_ (.A(_08989_),
    .B(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__nor2_1 _14367_ (.A(net954),
    .B(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__a211o_1 _14368_ (.A1(net954),
    .A2(_08990_),
    .B1(_08995_),
    .C1(net1766),
    .X(_08996_));
 sky130_fd_sc_hd__a211o_1 _14369_ (.A1(_08113_),
    .A2(_08996_),
    .B1(net662),
    .C1(net738),
    .X(_08997_));
 sky130_fd_sc_hd__o211a_1 _14370_ (.A1(\core.fetchProgramCounter[24] ),
    .A2(net619),
    .B1(_08997_),
    .C1(net1894),
    .X(_00155_));
 sky130_fd_sc_hd__a22o_2 _14371_ (.A1(\jtag.managementReadData[25] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net232),
    .X(_08998_));
 sky130_fd_sc_hd__nor2_1 _14372_ (.A(net467),
    .B(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__nand2_1 _14373_ (.A(net467),
    .B(_08998_),
    .Y(_09000_));
 sky130_fd_sc_hd__and2b_1 _14374_ (.A_N(_08999_),
    .B(_09000_),
    .X(_09001_));
 sky130_fd_sc_hd__o21a_1 _14375_ (.A1(_08989_),
    .A2(_08991_),
    .B1(_08992_),
    .X(_09002_));
 sky130_fd_sc_hd__xnor2_1 _14376_ (.A(_09001_),
    .B(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__mux2_1 _14377_ (.A0(_08998_),
    .A1(_09003_),
    .S(net953),
    .X(_09004_));
 sky130_fd_sc_hd__a21o_1 _14378_ (.A1(net1760),
    .A2(_09004_),
    .B1(_08147_),
    .X(_09005_));
 sky130_fd_sc_hd__or3_1 _14379_ (.A(net738),
    .B(net662),
    .C(_09005_),
    .X(_09006_));
 sky130_fd_sc_hd__o211a_1 _14380_ (.A1(\core.fetchProgramCounter[25] ),
    .A2(net619),
    .B1(_09006_),
    .C1(net1899),
    .X(_00156_));
 sky130_fd_sc_hd__a22o_2 _14381_ (.A1(\jtag.managementReadData[26] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net233),
    .X(_09007_));
 sky130_fd_sc_hd__nor2_1 _14382_ (.A(net468),
    .B(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__nand2_1 _14383_ (.A(net468),
    .B(_09007_),
    .Y(_09009_));
 sky130_fd_sc_hd__nand2b_1 _14384_ (.A_N(_09008_),
    .B(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__o21a_1 _14385_ (.A1(_08999_),
    .A2(_09002_),
    .B1(_09000_),
    .X(_09011_));
 sky130_fd_sc_hd__xor2_1 _14386_ (.A(_09010_),
    .B(_09011_),
    .X(_09012_));
 sky130_fd_sc_hd__mux2_1 _14387_ (.A0(_09007_),
    .A1(_09012_),
    .S(net953),
    .X(_09013_));
 sky130_fd_sc_hd__a21o_1 _14388_ (.A1(net1760),
    .A2(_09013_),
    .B1(_08137_),
    .X(_09014_));
 sky130_fd_sc_hd__or3_1 _14389_ (.A(net738),
    .B(net663),
    .C(_09014_),
    .X(_09015_));
 sky130_fd_sc_hd__o211a_1 _14390_ (.A1(\core.fetchProgramCounter[26] ),
    .A2(net620),
    .B1(_09015_),
    .C1(net1900),
    .X(_00157_));
 sky130_fd_sc_hd__a22o_4 _14391_ (.A1(\jtag.managementReadData[27] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net234),
    .X(_09016_));
 sky130_fd_sc_hd__xnor2_1 _14392_ (.A(net469),
    .B(_09016_),
    .Y(_09017_));
 sky130_fd_sc_hd__o21ai_2 _14393_ (.A1(_09008_),
    .A2(_09011_),
    .B1(_09009_),
    .Y(_09018_));
 sky130_fd_sc_hd__xnor2_1 _14394_ (.A(_09017_),
    .B(_09018_),
    .Y(_09019_));
 sky130_fd_sc_hd__mux2_1 _14395_ (.A0(_09016_),
    .A1(_09019_),
    .S(net953),
    .X(_09020_));
 sky130_fd_sc_hd__a21bo_1 _14396_ (.A1(net1760),
    .A2(_09020_),
    .B1_N(_08126_),
    .X(_09021_));
 sky130_fd_sc_hd__or3_1 _14397_ (.A(net739),
    .B(net663),
    .C(_09021_),
    .X(_09022_));
 sky130_fd_sc_hd__o211a_1 _14398_ (.A1(\core.fetchProgramCounter[27] ),
    .A2(net620),
    .B1(_09022_),
    .C1(net1899),
    .X(_00158_));
 sky130_fd_sc_hd__a22o_2 _14399_ (.A1(\jtag.managementReadData[28] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net235),
    .X(_09023_));
 sky130_fd_sc_hd__nor2_1 _14400_ (.A(net470),
    .B(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__nand2_1 _14401_ (.A(net470),
    .B(_09023_),
    .Y(_09025_));
 sky130_fd_sc_hd__nand2b_1 _14402_ (.A_N(_09024_),
    .B(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__a21o_1 _14403_ (.A1(net469),
    .A2(_09016_),
    .B1(_09018_),
    .X(_09027_));
 sky130_fd_sc_hd__o21ai_4 _14404_ (.A1(net469),
    .A2(_09016_),
    .B1(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__xor2_1 _14405_ (.A(_09026_),
    .B(_09028_),
    .X(_09029_));
 sky130_fd_sc_hd__or2_1 _14406_ (.A(net953),
    .B(_09023_),
    .X(_09030_));
 sky130_fd_sc_hd__o211a_1 _14407_ (.A1(net954),
    .A2(_09029_),
    .B1(_09030_),
    .C1(net1760),
    .X(_09031_));
 sky130_fd_sc_hd__a31o_1 _14408_ (.A1(net1767),
    .A2(_08031_),
    .A3(_08035_),
    .B1(_09031_),
    .X(_09032_));
 sky130_fd_sc_hd__or3_1 _14409_ (.A(net738),
    .B(net662),
    .C(_09032_),
    .X(_09033_));
 sky130_fd_sc_hd__o211a_1 _14410_ (.A1(\core.fetchProgramCounter[28] ),
    .A2(net619),
    .B1(_09033_),
    .C1(net1899),
    .X(_00159_));
 sky130_fd_sc_hd__a22o_4 _14411_ (.A1(\jtag.managementReadData[29] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net236),
    .X(_09034_));
 sky130_fd_sc_hd__nor2_1 _14412_ (.A(net471),
    .B(_09034_),
    .Y(_09035_));
 sky130_fd_sc_hd__and2_1 _14413_ (.A(net471),
    .B(_09034_),
    .X(_09036_));
 sky130_fd_sc_hd__or2_1 _14414_ (.A(_09035_),
    .B(_09036_),
    .X(_09037_));
 sky130_fd_sc_hd__o21ai_2 _14415_ (.A1(_09024_),
    .A2(_09028_),
    .B1(_09025_),
    .Y(_09038_));
 sky130_fd_sc_hd__xnor2_1 _14416_ (.A(_09037_),
    .B(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__mux2_1 _14417_ (.A0(_09034_),
    .A1(_09039_),
    .S(net953),
    .X(_09040_));
 sky130_fd_sc_hd__a21o_1 _14418_ (.A1(net1760),
    .A2(_09040_),
    .B1(_08050_),
    .X(_09041_));
 sky130_fd_sc_hd__or3_1 _14419_ (.A(net738),
    .B(net662),
    .C(_09041_),
    .X(_09042_));
 sky130_fd_sc_hd__o211a_1 _14420_ (.A1(\core.fetchProgramCounter[29] ),
    .A2(net619),
    .B1(_09042_),
    .C1(net1891),
    .X(_00160_));
 sky130_fd_sc_hd__a22o_2 _14421_ (.A1(\jtag.managementReadData[30] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net238),
    .X(_09043_));
 sky130_fd_sc_hd__and2_1 _14422_ (.A(net473),
    .B(_09043_),
    .X(_09044_));
 sky130_fd_sc_hd__nor2_1 _14423_ (.A(net473),
    .B(_09043_),
    .Y(_09045_));
 sky130_fd_sc_hd__nor2_1 _14424_ (.A(_09036_),
    .B(_09038_),
    .Y(_09046_));
 sky130_fd_sc_hd__o22a_1 _14425_ (.A1(_09044_),
    .A2(_09045_),
    .B1(_09046_),
    .B2(_09035_),
    .X(_09047_));
 sky130_fd_sc_hd__nor4_1 _14426_ (.A(_09035_),
    .B(_09044_),
    .C(_09045_),
    .D(_09046_),
    .Y(_09048_));
 sky130_fd_sc_hd__nor3_1 _14427_ (.A(net954),
    .B(_09047_),
    .C(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__a211o_1 _14428_ (.A1(net954),
    .A2(_09043_),
    .B1(_09049_),
    .C1(net1767),
    .X(_09050_));
 sky130_fd_sc_hd__a211o_1 _14429_ (.A1(_08023_),
    .A2(_09050_),
    .B1(net662),
    .C1(net738),
    .X(_09051_));
 sky130_fd_sc_hd__o211a_1 _14430_ (.A1(\core.fetchProgramCounter[30] ),
    .A2(net619),
    .B1(_09051_),
    .C1(net1889),
    .X(_00161_));
 sky130_fd_sc_hd__a22o_4 _14431_ (.A1(\jtag.managementReadData[31] ),
    .A2(net1367),
    .B1(net1298),
    .B2(net239),
    .X(_09052_));
 sky130_fd_sc_hd__nor2_1 _14432_ (.A(_09044_),
    .B(_09048_),
    .Y(_09053_));
 sky130_fd_sc_hd__nor2_1 _14433_ (.A(_04403_),
    .B(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__a211o_1 _14434_ (.A1(_04403_),
    .A2(_09053_),
    .B1(_09054_),
    .C1(net954),
    .X(_09055_));
 sky130_fd_sc_hd__xnor2_1 _14435_ (.A(_09052_),
    .B(_09055_),
    .Y(_09056_));
 sky130_fd_sc_hd__o21a_1 _14436_ (.A1(net1767),
    .A2(_09056_),
    .B1(_08010_),
    .X(_09057_));
 sky130_fd_sc_hd__or3_1 _14437_ (.A(net738),
    .B(net662),
    .C(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__o211a_1 _14438_ (.A1(\core.fetchProgramCounter[31] ),
    .A2(net619),
    .B1(_09058_),
    .C1(net1889),
    .X(_00162_));
 sky130_fd_sc_hd__or3b_2 _14439_ (.A(net1778),
    .B(net1779),
    .C_N(_08620_),
    .X(_09059_));
 sky130_fd_sc_hd__inv_2 _14440_ (.A(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__nand2_4 _14441_ (.A(net1781),
    .B(_08630_),
    .Y(_09061_));
 sky130_fd_sc_hd__nor2_1 _14442_ (.A(_09059_),
    .B(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__or3_1 _14443_ (.A(\jtag.dataBSRRegister.data[26] ),
    .B(_09059_),
    .C(_09061_),
    .X(_09063_));
 sky130_fd_sc_hd__or3_2 _14444_ (.A(\jtag.managementState[0] ),
    .B(net1639),
    .C(_09063_),
    .X(_09064_));
 sky130_fd_sc_hd__mux2_1 _14445_ (.A0(\jtag.dataBSRRegister.data[0] ),
    .A1(\jtag.managementAddress[0] ),
    .S(net1217),
    .X(_09065_));
 sky130_fd_sc_hd__and2_1 _14446_ (.A(net1932),
    .B(_09065_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _14447_ (.A0(\jtag.dataBSRRegister.data[1] ),
    .A1(\jtag.managementAddress[1] ),
    .S(net1217),
    .X(_09066_));
 sky130_fd_sc_hd__and2_1 _14448_ (.A(net1933),
    .B(_09066_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _14449_ (.A0(\jtag.dataBSRRegister.data[2] ),
    .A1(\jtag.managementAddress[2] ),
    .S(net1217),
    .X(_09067_));
 sky130_fd_sc_hd__and2_1 _14450_ (.A(net1936),
    .B(_09067_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _14451_ (.A0(\jtag.dataBSRRegister.data[3] ),
    .A1(\jtag.managementAddress[3] ),
    .S(net1216),
    .X(_09068_));
 sky130_fd_sc_hd__and2_1 _14452_ (.A(net1935),
    .B(_09068_),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _14453_ (.A0(\jtag.dataBSRRegister.data[4] ),
    .A1(\jtag.managementAddress[4] ),
    .S(net1216),
    .X(_09069_));
 sky130_fd_sc_hd__and2_1 _14454_ (.A(net1935),
    .B(_09069_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _14455_ (.A0(\jtag.dataBSRRegister.data[5] ),
    .A1(\jtag.managementAddress[5] ),
    .S(net1216),
    .X(_09070_));
 sky130_fd_sc_hd__and2_1 _14456_ (.A(net1953),
    .B(_09070_),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _14457_ (.A0(\jtag.dataBSRRegister.data[6] ),
    .A1(\jtag.managementAddress[6] ),
    .S(net1216),
    .X(_09071_));
 sky130_fd_sc_hd__and2_1 _14458_ (.A(net1943),
    .B(_09071_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _14459_ (.A0(\jtag.dataBSRRegister.data[7] ),
    .A1(\jtag.managementAddress[7] ),
    .S(net1216),
    .X(_09072_));
 sky130_fd_sc_hd__and2_1 _14460_ (.A(net1953),
    .B(_09072_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _14461_ (.A0(\jtag.dataBSRRegister.data[8] ),
    .A1(\jtag.managementAddress[8] ),
    .S(net1216),
    .X(_09073_));
 sky130_fd_sc_hd__and2_1 _14462_ (.A(net1953),
    .B(_09073_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _14463_ (.A0(\jtag.dataBSRRegister.data[9] ),
    .A1(\jtag.managementAddress[9] ),
    .S(net1216),
    .X(_09074_));
 sky130_fd_sc_hd__and2_1 _14464_ (.A(net1935),
    .B(_09074_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _14465_ (.A0(\jtag.dataBSRRegister.data[10] ),
    .A1(\jtag.managementAddress[10] ),
    .S(net1216),
    .X(_09075_));
 sky130_fd_sc_hd__and2_1 _14466_ (.A(net1936),
    .B(_09075_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _14467_ (.A0(\jtag.dataBSRRegister.data[11] ),
    .A1(\jtag.managementAddress[11] ),
    .S(net1216),
    .X(_09076_));
 sky130_fd_sc_hd__and2_1 _14468_ (.A(net1936),
    .B(_09076_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _14469_ (.A0(\jtag.dataBSRRegister.data[12] ),
    .A1(\jtag.managementAddress[12] ),
    .S(net1216),
    .X(_09077_));
 sky130_fd_sc_hd__and2_1 _14470_ (.A(net1936),
    .B(_09077_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _14471_ (.A0(\jtag.dataBSRRegister.data[13] ),
    .A1(\jtag.managementAddress[13] ),
    .S(net1217),
    .X(_09078_));
 sky130_fd_sc_hd__and2_1 _14472_ (.A(net1933),
    .B(_09078_),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _14473_ (.A0(\jtag.dataBSRRegister.data[14] ),
    .A1(\jtag.managementAddress[14] ),
    .S(net1217),
    .X(_09079_));
 sky130_fd_sc_hd__and2_1 _14474_ (.A(net1932),
    .B(_09079_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _14475_ (.A0(\jtag.dataBSRRegister.data[15] ),
    .A1(\jtag.managementAddress[15] ),
    .S(net1217),
    .X(_09080_));
 sky130_fd_sc_hd__and2_1 _14476_ (.A(net1917),
    .B(_09080_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _14477_ (.A0(\jtag.dataBSRRegister.data[16] ),
    .A1(\jtag.managementAddress[16] ),
    .S(net1217),
    .X(_09081_));
 sky130_fd_sc_hd__and2_1 _14478_ (.A(net1917),
    .B(_09081_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _14479_ (.A0(\jtag.dataBSRRegister.data[17] ),
    .A1(\jtag.managementAddress[17] ),
    .S(net1218),
    .X(_09082_));
 sky130_fd_sc_hd__and2_1 _14480_ (.A(net1901),
    .B(_09082_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _14481_ (.A0(\jtag.dataBSRRegister.data[18] ),
    .A1(\jtag.managementAddress[18] ),
    .S(net1218),
    .X(_09083_));
 sky130_fd_sc_hd__and2_1 _14482_ (.A(net1904),
    .B(_09083_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _14483_ (.A0(\jtag.dataBSRRegister.data[19] ),
    .A1(\jtag.managementAddress[19] ),
    .S(net1218),
    .X(_09084_));
 sky130_fd_sc_hd__and2_1 _14484_ (.A(net1901),
    .B(_09084_),
    .X(_00182_));
 sky130_fd_sc_hd__o211a_1 _14485_ (.A1(_04512_),
    .A2(_04516_),
    .B1(_04526_),
    .C1(net1923),
    .X(_09085_));
 sky130_fd_sc_hd__or3_2 _14486_ (.A(\core.csr.currentInstruction[10] ),
    .B(_04424_),
    .C(_04513_),
    .X(_09086_));
 sky130_fd_sc_hd__nor2_1 _14487_ (.A(_04512_),
    .B(_09086_),
    .Y(_09087_));
 sky130_fd_sc_hd__and3_4 _14488_ (.A(net676),
    .B(net1072),
    .C(_09087_),
    .X(_09088_));
 sky130_fd_sc_hd__mux2_1 _14489_ (.A0(\core.registers[20][0] ),
    .A1(net1037),
    .S(net617),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _14490_ (.A0(\core.registers[20][1] ),
    .A1(net1039),
    .S(net617),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _14491_ (.A0(\core.registers[20][2] ),
    .A1(net1044),
    .S(net618),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _14492_ (.A0(\core.registers[20][3] ),
    .A1(net1048),
    .S(net617),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _14493_ (.A0(\core.registers[20][4] ),
    .A1(net1053),
    .S(net617),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _14494_ (.A0(\core.registers[20][5] ),
    .A1(net1057),
    .S(net618),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _14495_ (.A0(\core.registers[20][6] ),
    .A1(net1061),
    .S(net618),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _14496_ (.A0(\core.registers[20][7] ),
    .A1(net1133),
    .S(net618),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _14497_ (.A0(\core.registers[20][8] ),
    .A1(net959),
    .S(net618),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _14498_ (.A0(\core.registers[20][9] ),
    .A1(net962),
    .S(net616),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _14499_ (.A0(\core.registers[20][10] ),
    .A1(net969),
    .S(net617),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _14500_ (.A0(\core.registers[20][11] ),
    .A1(net972),
    .S(net616),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _14501_ (.A0(\core.registers[20][12] ),
    .A1(net989),
    .S(net616),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _14502_ (.A0(\core.registers[20][13] ),
    .A1(net985),
    .S(net617),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _14503_ (.A0(\core.registers[20][14] ),
    .A1(net974),
    .S(net617),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _14504_ (.A0(\core.registers[20][15] ),
    .A1(net981),
    .S(net617),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _14505_ (.A0(\core.registers[20][16] ),
    .A1(net1124),
    .S(net615),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _14506_ (.A0(\core.registers[20][17] ),
    .A1(net1129),
    .S(net615),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _14507_ (.A0(\core.registers[20][18] ),
    .A1(net1116),
    .S(net615),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _14508_ (.A0(\core.registers[20][19] ),
    .A1(net1120),
    .S(net615),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _14509_ (.A0(\core.registers[20][20] ),
    .A1(net1138),
    .S(net615),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _14510_ (.A0(\core.registers[20][21] ),
    .A1(net1142),
    .S(net615),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _14511_ (.A0(\core.registers[20][22] ),
    .A1(net1147),
    .S(net616),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _14512_ (.A0(\core.registers[20][23] ),
    .A1(net1151),
    .S(net615),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _14513_ (.A0(\core.registers[20][24] ),
    .A1(net1115),
    .S(net615),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _14514_ (.A0(\core.registers[20][25] ),
    .A1(net1108),
    .S(net615),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _14515_ (.A0(\core.registers[20][26] ),
    .A1(net1102),
    .S(net616),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _14516_ (.A0(\core.registers[20][27] ),
    .A1(net1106),
    .S(net616),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _14517_ (.A0(\core.registers[20][28] ),
    .A1(net1098),
    .S(net615),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _14518_ (.A0(\core.registers[20][29] ),
    .A1(net1092),
    .S(net617),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _14519_ (.A0(\core.registers[20][30] ),
    .A1(net1084),
    .S(net618),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _14520_ (.A0(\core.registers[20][31] ),
    .A1(net1089),
    .S(net617),
    .X(_00214_));
 sky130_fd_sc_hd__a21oi_1 _14521_ (.A1(net806),
    .A2(net697),
    .B1(\core.memoryOperationCompleted ),
    .Y(_09089_));
 sky130_fd_sc_hd__nor2_1 _14522_ (.A(_08650_),
    .B(_09089_),
    .Y(_00215_));
 sky130_fd_sc_hd__o21ba_1 _14523_ (.A1(_08096_),
    .A2(_08642_),
    .B1_N(_08639_),
    .X(_09090_));
 sky130_fd_sc_hd__o21a_1 _14524_ (.A1(net1765),
    .A2(_09090_),
    .B1(net1814),
    .X(_09091_));
 sky130_fd_sc_hd__and3_1 _14525_ (.A(\core.memoryOperationCompleted ),
    .B(net807),
    .C(net678),
    .X(_09092_));
 sky130_fd_sc_hd__o21a_1 _14526_ (.A1(_09091_),
    .A2(_09092_),
    .B1(net1908),
    .X(_00216_));
 sky130_fd_sc_hd__a311oi_1 _14527_ (.A1(\core.management_pipeStartup ),
    .A2(net683),
    .A3(_08762_),
    .B1(net1989),
    .C1(_07878_),
    .Y(_00217_));
 sky130_fd_sc_hd__or2_4 _14528_ (.A(_04425_),
    .B(_04511_),
    .X(_09093_));
 sky130_fd_sc_hd__or3_2 _14529_ (.A(\core.csr.currentInstruction[10] ),
    .B(\core.csr.currentInstruction[9] ),
    .C(_04513_),
    .X(_09094_));
 sky130_fd_sc_hd__nor2_1 _14530_ (.A(_09093_),
    .B(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__and3_4 _14531_ (.A(net679),
    .B(net1075),
    .C(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__mux2_1 _14532_ (.A0(\core.registers[19][0] ),
    .A1(net1037),
    .S(net613),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _14533_ (.A0(\core.registers[19][1] ),
    .A1(net1040),
    .S(net613),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _14534_ (.A0(\core.registers[19][2] ),
    .A1(net1044),
    .S(net613),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _14535_ (.A0(\core.registers[19][3] ),
    .A1(net1048),
    .S(net613),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _14536_ (.A0(\core.registers[19][4] ),
    .A1(net1054),
    .S(net613),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _14537_ (.A0(\core.registers[19][5] ),
    .A1(net1057),
    .S(net614),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _14538_ (.A0(\core.registers[19][6] ),
    .A1(net1061),
    .S(net614),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _14539_ (.A0(\core.registers[19][7] ),
    .A1(net1133),
    .S(net614),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _14540_ (.A0(\core.registers[19][8] ),
    .A1(net960),
    .S(net614),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _14541_ (.A0(\core.registers[19][9] ),
    .A1(net963),
    .S(net612),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _14542_ (.A0(\core.registers[19][10] ),
    .A1(net968),
    .S(net613),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _14543_ (.A0(\core.registers[19][11] ),
    .A1(net972),
    .S(net612),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _14544_ (.A0(\core.registers[19][12] ),
    .A1(net989),
    .S(net612),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _14545_ (.A0(\core.registers[19][13] ),
    .A1(net986),
    .S(net614),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _14546_ (.A0(\core.registers[19][14] ),
    .A1(net974),
    .S(net613),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _14547_ (.A0(\core.registers[19][15] ),
    .A1(net981),
    .S(net613),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _14548_ (.A0(\core.registers[19][16] ),
    .A1(net1124),
    .S(net611),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _14549_ (.A0(\core.registers[19][17] ),
    .A1(net1130),
    .S(net611),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _14550_ (.A0(\core.registers[19][18] ),
    .A1(net1117),
    .S(net612),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _14551_ (.A0(\core.registers[19][19] ),
    .A1(net1123),
    .S(net611),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _14552_ (.A0(\core.registers[19][20] ),
    .A1(net1138),
    .S(net611),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _14553_ (.A0(\core.registers[19][21] ),
    .A1(net1142),
    .S(net611),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _14554_ (.A0(\core.registers[19][22] ),
    .A1(net1147),
    .S(net612),
    .X(_00240_));
 sky130_fd_sc_hd__mux2_1 _14555_ (.A0(\core.registers[19][23] ),
    .A1(net1151),
    .S(net611),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _14556_ (.A0(\core.registers[19][24] ),
    .A1(net1114),
    .S(net611),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _14557_ (.A0(\core.registers[19][25] ),
    .A1(net1109),
    .S(net611),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _14558_ (.A0(\core.registers[19][26] ),
    .A1(net1102),
    .S(net612),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _14559_ (.A0(\core.registers[19][27] ),
    .A1(net1106),
    .S(net611),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _14560_ (.A0(\core.registers[19][28] ),
    .A1(net1096),
    .S(net611),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _14561_ (.A0(\core.registers[19][29] ),
    .A1(net1092),
    .S(net613),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _14562_ (.A0(\core.registers[19][30] ),
    .A1(net1084),
    .S(net614),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _14563_ (.A0(\core.registers[19][31] ),
    .A1(net1089),
    .S(net613),
    .X(_00249_));
 sky130_fd_sc_hd__or2_4 _14564_ (.A(\core.csr.currentInstruction[7] ),
    .B(_04511_),
    .X(_09097_));
 sky130_fd_sc_hd__or3_2 _14565_ (.A(_04424_),
    .B(_04513_),
    .C(_04514_),
    .X(_09098_));
 sky130_fd_sc_hd__nor2_1 _14566_ (.A(_09097_),
    .B(_09098_),
    .Y(_09099_));
 sky130_fd_sc_hd__and3_4 _14567_ (.A(net679),
    .B(net1074),
    .C(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__mux2_1 _14568_ (.A0(\core.registers[30][0] ),
    .A1(net1035),
    .S(net610),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _14569_ (.A0(\core.registers[30][1] ),
    .A1(net1041),
    .S(net610),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _14570_ (.A0(\core.registers[30][2] ),
    .A1(net1043),
    .S(net609),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _14571_ (.A0(\core.registers[30][3] ),
    .A1(net1050),
    .S(net609),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _14572_ (.A0(\core.registers[30][4] ),
    .A1(net1055),
    .S(net610),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _14573_ (.A0(\core.registers[30][5] ),
    .A1(net1059),
    .S(net609),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _14574_ (.A0(\core.registers[30][6] ),
    .A1(net1064),
    .S(net609),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _14575_ (.A0(\core.registers[30][7] ),
    .A1(net1134),
    .S(net609),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _14576_ (.A0(\core.registers[30][8] ),
    .A1(net957),
    .S(net609),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _14577_ (.A0(\core.registers[30][9] ),
    .A1(net962),
    .S(net608),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _14578_ (.A0(\core.registers[30][10] ),
    .A1(net966),
    .S(net610),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _14579_ (.A0(\core.registers[30][11] ),
    .A1(net970),
    .S(net608),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _14580_ (.A0(\core.registers[30][12] ),
    .A1(net988),
    .S(net610),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _14581_ (.A0(\core.registers[30][13] ),
    .A1(net984),
    .S(net609),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _14582_ (.A0(\core.registers[30][14] ),
    .A1(net974),
    .S(net610),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _14583_ (.A0(\core.registers[30][15] ),
    .A1(net979),
    .S(net609),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _14584_ (.A0(\core.registers[30][16] ),
    .A1(net1127),
    .S(net607),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _14585_ (.A0(\core.registers[30][17] ),
    .A1(net1131),
    .S(net607),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _14586_ (.A0(\core.registers[30][18] ),
    .A1(net1117),
    .S(net608),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _14587_ (.A0(\core.registers[30][19] ),
    .A1(net1121),
    .S(net607),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _14588_ (.A0(\core.registers[30][20] ),
    .A1(net1137),
    .S(net607),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _14589_ (.A0(\core.registers[30][21] ),
    .A1(net1141),
    .S(net607),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _14590_ (.A0(\core.registers[30][22] ),
    .A1(net1146),
    .S(net608),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _14591_ (.A0(\core.registers[30][23] ),
    .A1(net1149),
    .S(net607),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _14592_ (.A0(\core.registers[30][24] ),
    .A1(net1113),
    .S(net607),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _14593_ (.A0(\core.registers[30][25] ),
    .A1(net1108),
    .S(net607),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _14594_ (.A0(\core.registers[30][26] ),
    .A1(net1100),
    .S(net608),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _14595_ (.A0(\core.registers[30][27] ),
    .A1(net1104),
    .S(net607),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _14596_ (.A0(\core.registers[30][28] ),
    .A1(net1098),
    .S(net607),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _14597_ (.A0(\core.registers[30][29] ),
    .A1(net1095),
    .S(net609),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _14598_ (.A0(\core.registers[30][30] ),
    .A1(net1086),
    .S(net609),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _14599_ (.A0(\core.registers[30][31] ),
    .A1(net1091),
    .S(net610),
    .X(_00281_));
 sky130_fd_sc_hd__nor2_1 _14600_ (.A(_04516_),
    .B(_09097_),
    .Y(_09101_));
 sky130_fd_sc_hd__and3_4 _14601_ (.A(net679),
    .B(net1075),
    .C(_09101_),
    .X(_09102_));
 sky130_fd_sc_hd__mux2_1 _14602_ (.A0(\core.registers[2][0] ),
    .A1(net1038),
    .S(net605),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _14603_ (.A0(\core.registers[2][1] ),
    .A1(net1042),
    .S(net605),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _14604_ (.A0(\core.registers[2][2] ),
    .A1(net1045),
    .S(net605),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _14605_ (.A0(\core.registers[2][3] ),
    .A1(net1049),
    .S(net605),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _14606_ (.A0(\core.registers[2][4] ),
    .A1(net1053),
    .S(net605),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _14607_ (.A0(\core.registers[2][5] ),
    .A1(net1060),
    .S(net606),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _14608_ (.A0(\core.registers[2][6] ),
    .A1(net1063),
    .S(net606),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _14609_ (.A0(\core.registers[2][7] ),
    .A1(net1135),
    .S(net606),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _14610_ (.A0(\core.registers[2][8] ),
    .A1(net960),
    .S(net606),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _14611_ (.A0(\core.registers[2][9] ),
    .A1(net965),
    .S(net604),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _14612_ (.A0(\core.registers[2][10] ),
    .A1(net969),
    .S(net605),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _14613_ (.A0(\core.registers[2][11] ),
    .A1(net2011),
    .S(net604),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _14614_ (.A0(\core.registers[2][12] ),
    .A1(net990),
    .S(net604),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _14615_ (.A0(\core.registers[2][13] ),
    .A1(net985),
    .S(net605),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _14616_ (.A0(\core.registers[2][14] ),
    .A1(net978),
    .S(net604),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _14617_ (.A0(\core.registers[2][15] ),
    .A1(net981),
    .S(net605),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _14618_ (.A0(\core.registers[2][16] ),
    .A1(net1126),
    .S(net603),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _14619_ (.A0(\core.registers[2][17] ),
    .A1(net1129),
    .S(net603),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _14620_ (.A0(\core.registers[2][18] ),
    .A1(net1119),
    .S(net604),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _14621_ (.A0(\core.registers[2][19] ),
    .A1(net1122),
    .S(net603),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _14622_ (.A0(\core.registers[2][20] ),
    .A1(net1139),
    .S(net603),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _14623_ (.A0(\core.registers[2][21] ),
    .A1(net1143),
    .S(net603),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _14624_ (.A0(\core.registers[2][22] ),
    .A1(net1148),
    .S(net604),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _14625_ (.A0(\core.registers[2][23] ),
    .A1(net1152),
    .S(net603),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _14626_ (.A0(\core.registers[2][24] ),
    .A1(net1114),
    .S(net603),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _14627_ (.A0(\core.registers[2][25] ),
    .A1(net1109),
    .S(net603),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _14628_ (.A0(\core.registers[2][26] ),
    .A1(net1103),
    .S(net604),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _14629_ (.A0(\core.registers[2][27] ),
    .A1(net1107),
    .S(net603),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _14630_ (.A0(\core.registers[2][28] ),
    .A1(net1097),
    .S(net603),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _14631_ (.A0(\core.registers[2][29] ),
    .A1(net1092),
    .S(net605),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _14632_ (.A0(\core.registers[2][30] ),
    .A1(net1087),
    .S(net606),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _14633_ (.A0(\core.registers[2][31] ),
    .A1(net1090),
    .S(net605),
    .X(_00313_));
 sky130_fd_sc_hd__nor2_1 _14634_ (.A(_04512_),
    .B(_09098_),
    .Y(_09103_));
 sky130_fd_sc_hd__and3_4 _14635_ (.A(net679),
    .B(net1074),
    .C(_09103_),
    .X(_09104_));
 sky130_fd_sc_hd__mux2_1 _14636_ (.A0(\core.registers[28][0] ),
    .A1(net1036),
    .S(net601),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _14637_ (.A0(\core.registers[28][1] ),
    .A1(net1041),
    .S(net602),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _14638_ (.A0(\core.registers[28][2] ),
    .A1(net1047),
    .S(net602),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _14639_ (.A0(\core.registers[28][3] ),
    .A1(net1050),
    .S(net601),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _14640_ (.A0(\core.registers[28][4] ),
    .A1(net1055),
    .S(net602),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _14641_ (.A0(\core.registers[28][5] ),
    .A1(net1059),
    .S(net601),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _14642_ (.A0(\core.registers[28][6] ),
    .A1(net1064),
    .S(net601),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _14643_ (.A0(\core.registers[28][7] ),
    .A1(net1134),
    .S(net601),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _14644_ (.A0(\core.registers[28][8] ),
    .A1(net958),
    .S(net602),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _14645_ (.A0(\core.registers[28][9] ),
    .A1(net962),
    .S(net600),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _14646_ (.A0(\core.registers[28][10] ),
    .A1(net966),
    .S(net602),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _14647_ (.A0(\core.registers[28][11] ),
    .A1(net970),
    .S(net599),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _14648_ (.A0(\core.registers[28][12] ),
    .A1(net988),
    .S(net602),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _14649_ (.A0(\core.registers[28][13] ),
    .A1(net983),
    .S(net601),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _14650_ (.A0(\core.registers[28][14] ),
    .A1(net974),
    .S(net602),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _14651_ (.A0(\core.registers[28][15] ),
    .A1(net979),
    .S(net601),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(\core.registers[28][16] ),
    .A1(net1127),
    .S(net599),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _14653_ (.A0(\core.registers[28][17] ),
    .A1(net1131),
    .S(net599),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _14654_ (.A0(\core.registers[28][18] ),
    .A1(net1117),
    .S(net600),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _14655_ (.A0(\core.registers[28][19] ),
    .A1(net1122),
    .S(net600),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _14656_ (.A0(\core.registers[28][20] ),
    .A1(net1136),
    .S(net599),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _14657_ (.A0(\core.registers[28][21] ),
    .A1(net1140),
    .S(net599),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _14658_ (.A0(\core.registers[28][22] ),
    .A1(net1145),
    .S(net600),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _14659_ (.A0(\core.registers[28][23] ),
    .A1(net1149),
    .S(net599),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _14660_ (.A0(\core.registers[28][24] ),
    .A1(net1112),
    .S(net599),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _14661_ (.A0(\core.registers[28][25] ),
    .A1(net1110),
    .S(net599),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _14662_ (.A0(\core.registers[28][26] ),
    .A1(net1100),
    .S(net600),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _14663_ (.A0(\core.registers[28][27] ),
    .A1(net1104),
    .S(net599),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _14664_ (.A0(\core.registers[28][28] ),
    .A1(net1098),
    .S(net599),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _14665_ (.A0(\core.registers[28][29] ),
    .A1(net1095),
    .S(net601),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _14666_ (.A0(\core.registers[28][30] ),
    .A1(net1086),
    .S(net601),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _14667_ (.A0(\core.registers[28][31] ),
    .A1(net1091),
    .S(net601),
    .X(_00345_));
 sky130_fd_sc_hd__or3_2 _14668_ (.A(\core.csr.currentInstruction[9] ),
    .B(_04513_),
    .C(_04514_),
    .X(_09105_));
 sky130_fd_sc_hd__nor2_1 _14669_ (.A(_09093_),
    .B(_09105_),
    .Y(_09106_));
 sky130_fd_sc_hd__and3_4 _14670_ (.A(net680),
    .B(net1075),
    .C(_09106_),
    .X(_09107_));
 sky130_fd_sc_hd__mux2_1 _14671_ (.A0(\core.registers[27][0] ),
    .A1(net1036),
    .S(net598),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _14672_ (.A0(\core.registers[27][1] ),
    .A1(net1039),
    .S(net597),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _14673_ (.A0(\core.registers[27][2] ),
    .A1(net1043),
    .S(net597),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _14674_ (.A0(\core.registers[27][3] ),
    .A1(net1050),
    .S(net598),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _14675_ (.A0(\core.registers[27][4] ),
    .A1(net1056),
    .S(net598),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _14676_ (.A0(\core.registers[27][5] ),
    .A1(net1058),
    .S(net598),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _14677_ (.A0(\core.registers[27][6] ),
    .A1(net1061),
    .S(net597),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _14678_ (.A0(\core.registers[27][7] ),
    .A1(net1132),
    .S(net597),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _14679_ (.A0(\core.registers[27][8] ),
    .A1(net957),
    .S(net597),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _14680_ (.A0(\core.registers[27][9] ),
    .A1(net962),
    .S(net596),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _14681_ (.A0(\core.registers[27][10] ),
    .A1(net966),
    .S(net598),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _14682_ (.A0(\core.registers[27][11] ),
    .A1(net971),
    .S(net596),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _14683_ (.A0(\core.registers[27][12] ),
    .A1(net987),
    .S(net596),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _14684_ (.A0(\core.registers[27][13] ),
    .A1(net983),
    .S(net597),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _14685_ (.A0(\core.registers[27][14] ),
    .A1(net976),
    .S(net598),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _14686_ (.A0(\core.registers[27][15] ),
    .A1(net979),
    .S(net597),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _14687_ (.A0(\core.registers[27][16] ),
    .A1(net1127),
    .S(net595),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _14688_ (.A0(\core.registers[27][17] ),
    .A1(net1131),
    .S(net595),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _14689_ (.A0(\core.registers[27][18] ),
    .A1(net1117),
    .S(net595),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _14690_ (.A0(\core.registers[27][19] ),
    .A1(net1121),
    .S(net595),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _14691_ (.A0(\core.registers[27][20] ),
    .A1(net1137),
    .S(net595),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _14692_ (.A0(\core.registers[27][21] ),
    .A1(net1141),
    .S(net595),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _14693_ (.A0(\core.registers[27][22] ),
    .A1(net1145),
    .S(net596),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _14694_ (.A0(\core.registers[27][23] ),
    .A1(net1149),
    .S(net595),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _14695_ (.A0(\core.registers[27][24] ),
    .A1(net1113),
    .S(net595),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _14696_ (.A0(\core.registers[27][25] ),
    .A1(net1109),
    .S(net595),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _14697_ (.A0(\core.registers[27][26] ),
    .A1(net1100),
    .S(net596),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _14698_ (.A0(\core.registers[27][27] ),
    .A1(net1104),
    .S(net595),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _14699_ (.A0(\core.registers[27][28] ),
    .A1(net1098),
    .S(net596),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _14700_ (.A0(\core.registers[27][29] ),
    .A1(net1094),
    .S(net597),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _14701_ (.A0(\core.registers[27][30] ),
    .A1(net1084),
    .S(net597),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _14702_ (.A0(\core.registers[27][31] ),
    .A1(net1088),
    .S(net597),
    .X(_00377_));
 sky130_fd_sc_hd__nor2_1 _14703_ (.A(_09097_),
    .B(_09105_),
    .Y(_09108_));
 sky130_fd_sc_hd__and3_4 _14704_ (.A(net680),
    .B(net1075),
    .C(_09108_),
    .X(_09109_));
 sky130_fd_sc_hd__mux2_1 _14705_ (.A0(\core.registers[26][0] ),
    .A1(net1036),
    .S(net594),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _14706_ (.A0(\core.registers[26][1] ),
    .A1(net1039),
    .S(net593),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _14707_ (.A0(\core.registers[26][2] ),
    .A1(net1046),
    .S(net593),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _14708_ (.A0(\core.registers[26][3] ),
    .A1(net1051),
    .S(net594),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _14709_ (.A0(\core.registers[26][4] ),
    .A1(net1056),
    .S(net594),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _14710_ (.A0(\core.registers[26][5] ),
    .A1(net1058),
    .S(net594),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _14711_ (.A0(\core.registers[26][6] ),
    .A1(net1061),
    .S(net593),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _14712_ (.A0(\core.registers[26][7] ),
    .A1(net1132),
    .S(net593),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _14713_ (.A0(\core.registers[26][8] ),
    .A1(net957),
    .S(net593),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _14714_ (.A0(\core.registers[26][9] ),
    .A1(net962),
    .S(net592),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _14715_ (.A0(\core.registers[26][10] ),
    .A1(net966),
    .S(net594),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _14716_ (.A0(\core.registers[26][11] ),
    .A1(net971),
    .S(net594),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _14717_ (.A0(\core.registers[26][12] ),
    .A1(net987),
    .S(net592),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _14718_ (.A0(\core.registers[26][13] ),
    .A1(net983),
    .S(net593),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _14719_ (.A0(\core.registers[26][14] ),
    .A1(net976),
    .S(net594),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _14720_ (.A0(\core.registers[26][15] ),
    .A1(net980),
    .S(net593),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _14721_ (.A0(\core.registers[26][16] ),
    .A1(net1127),
    .S(net591),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _14722_ (.A0(\core.registers[26][17] ),
    .A1(net1131),
    .S(net591),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _14723_ (.A0(\core.registers[26][18] ),
    .A1(net1117),
    .S(net591),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _14724_ (.A0(\core.registers[26][19] ),
    .A1(net1121),
    .S(net591),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _14725_ (.A0(\core.registers[26][20] ),
    .A1(net1137),
    .S(net591),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _14726_ (.A0(\core.registers[26][21] ),
    .A1(net1141),
    .S(net591),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _14727_ (.A0(\core.registers[26][22] ),
    .A1(net1145),
    .S(net592),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _14728_ (.A0(\core.registers[26][23] ),
    .A1(net1149),
    .S(net591),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _14729_ (.A0(\core.registers[26][24] ),
    .A1(net1113),
    .S(net591),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _14730_ (.A0(\core.registers[26][25] ),
    .A1(net1109),
    .S(net591),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _14731_ (.A0(\core.registers[26][26] ),
    .A1(net1100),
    .S(net592),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _14732_ (.A0(\core.registers[26][27] ),
    .A1(net1104),
    .S(net591),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _14733_ (.A0(\core.registers[26][28] ),
    .A1(net1098),
    .S(net592),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _14734_ (.A0(\core.registers[26][29] ),
    .A1(net1094),
    .S(net593),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _14735_ (.A0(\core.registers[26][30] ),
    .A1(net1084),
    .S(net593),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _14736_ (.A0(\core.registers[26][31] ),
    .A1(net1088),
    .S(net593),
    .X(_00409_));
 sky130_fd_sc_hd__and3b_4 _14737_ (.A_N(\core.pipe0_fetch.currentPipeStall ),
    .B(_08639_),
    .C(net697),
    .X(_09110_));
 sky130_fd_sc_hd__nand2b_4 _14738_ (.A_N(\core.pipe0_fetch.currentPipeStall ),
    .B(net678),
    .Y(_09111_));
 sky130_fd_sc_hd__or2_1 _14739_ (.A(net450),
    .B(net658),
    .X(_09112_));
 sky130_fd_sc_hd__o211a_1 _14740_ (.A1(\core.csr.instruction_memoryAddress[0] ),
    .A2(net587),
    .B1(_09112_),
    .C1(net1893),
    .X(_00410_));
 sky130_fd_sc_hd__or2_1 _14741_ (.A(net461),
    .B(net658),
    .X(_09113_));
 sky130_fd_sc_hd__o211a_1 _14742_ (.A1(\core.csr.instruction_memoryAddress[1] ),
    .A2(net587),
    .B1(_09113_),
    .C1(net1893),
    .X(_00411_));
 sky130_fd_sc_hd__or2_1 _14743_ (.A(net472),
    .B(net660),
    .X(_09114_));
 sky130_fd_sc_hd__o211a_1 _14744_ (.A1(\core.csr.instruction_memoryAddress[2] ),
    .A2(net589),
    .B1(_09114_),
    .C1(net1913),
    .X(_00412_));
 sky130_fd_sc_hd__or2_1 _14745_ (.A(net475),
    .B(net661),
    .X(_09115_));
 sky130_fd_sc_hd__o211a_1 _14746_ (.A1(\core.csr.instruction_memoryAddress[3] ),
    .A2(net589),
    .B1(_09115_),
    .C1(net1914),
    .X(_00413_));
 sky130_fd_sc_hd__or2_1 _14747_ (.A(net476),
    .B(net660),
    .X(_09116_));
 sky130_fd_sc_hd__o211a_1 _14748_ (.A1(\core.csr.instruction_memoryAddress[4] ),
    .A2(net589),
    .B1(_09116_),
    .C1(net1913),
    .X(_00414_));
 sky130_fd_sc_hd__or2_1 _14749_ (.A(net477),
    .B(net660),
    .X(_09117_));
 sky130_fd_sc_hd__o211a_1 _14750_ (.A1(\core.csr.instruction_memoryAddress[5] ),
    .A2(net589),
    .B1(_09117_),
    .C1(net1913),
    .X(_00415_));
 sky130_fd_sc_hd__or2_1 _14751_ (.A(net478),
    .B(net660),
    .X(_09118_));
 sky130_fd_sc_hd__o211a_1 _14752_ (.A1(\core.csr.instruction_memoryAddress[6] ),
    .A2(net589),
    .B1(_09118_),
    .C1(net1931),
    .X(_00416_));
 sky130_fd_sc_hd__or2_1 _14753_ (.A(net479),
    .B(net660),
    .X(_09119_));
 sky130_fd_sc_hd__o211a_1 _14754_ (.A1(\core.csr.instruction_memoryAddress[7] ),
    .A2(net589),
    .B1(_09119_),
    .C1(net1930),
    .X(_00417_));
 sky130_fd_sc_hd__or2_1 _14755_ (.A(net480),
    .B(net660),
    .X(_09120_));
 sky130_fd_sc_hd__o211a_1 _14756_ (.A1(\core.csr.instruction_memoryAddress[8] ),
    .A2(net589),
    .B1(_09120_),
    .C1(net1931),
    .X(_00418_));
 sky130_fd_sc_hd__or2_1 _14757_ (.A(net481),
    .B(net660),
    .X(_09121_));
 sky130_fd_sc_hd__o211a_1 _14758_ (.A1(\core.csr.instruction_memoryAddress[9] ),
    .A2(net590),
    .B1(_09121_),
    .C1(net1913),
    .X(_00419_));
 sky130_fd_sc_hd__or2_1 _14759_ (.A(net451),
    .B(net660),
    .X(_09122_));
 sky130_fd_sc_hd__o211a_1 _14760_ (.A1(\core.csr.instruction_memoryAddress[10] ),
    .A2(net589),
    .B1(_09122_),
    .C1(net1915),
    .X(_00420_));
 sky130_fd_sc_hd__or2_1 _14761_ (.A(net452),
    .B(net660),
    .X(_09123_));
 sky130_fd_sc_hd__o211a_1 _14762_ (.A1(\core.csr.instruction_memoryAddress[11] ),
    .A2(net589),
    .B1(_09123_),
    .C1(net1915),
    .X(_00421_));
 sky130_fd_sc_hd__or2_1 _14763_ (.A(net453),
    .B(net660),
    .X(_09124_));
 sky130_fd_sc_hd__o211a_1 _14764_ (.A1(\core.csr.instruction_memoryAddress[12] ),
    .A2(net589),
    .B1(_09124_),
    .C1(net1915),
    .X(_00422_));
 sky130_fd_sc_hd__or2_1 _14765_ (.A(net454),
    .B(net661),
    .X(_09125_));
 sky130_fd_sc_hd__o211a_1 _14766_ (.A1(\core.csr.instruction_memoryAddress[13] ),
    .A2(net590),
    .B1(_09125_),
    .C1(net1909),
    .X(_00423_));
 sky130_fd_sc_hd__or2_1 _14767_ (.A(net455),
    .B(net661),
    .X(_09126_));
 sky130_fd_sc_hd__o211a_1 _14768_ (.A1(\core.csr.instruction_memoryAddress[14] ),
    .A2(net590),
    .B1(_09126_),
    .C1(net1910),
    .X(_00424_));
 sky130_fd_sc_hd__or2_1 _14769_ (.A(net456),
    .B(net661),
    .X(_09127_));
 sky130_fd_sc_hd__o211a_1 _14770_ (.A1(\core.csr.instruction_memoryAddress[15] ),
    .A2(net590),
    .B1(_09127_),
    .C1(net1910),
    .X(_00425_));
 sky130_fd_sc_hd__or2_1 _14771_ (.A(net457),
    .B(net661),
    .X(_09128_));
 sky130_fd_sc_hd__o211a_1 _14772_ (.A1(\core.csr.instruction_memoryAddress[16] ),
    .A2(net590),
    .B1(_09128_),
    .C1(net1910),
    .X(_00426_));
 sky130_fd_sc_hd__or2_1 _14773_ (.A(net458),
    .B(net661),
    .X(_09129_));
 sky130_fd_sc_hd__o211a_1 _14774_ (.A1(\core.csr.instruction_memoryAddress[17] ),
    .A2(net590),
    .B1(_09129_),
    .C1(net1909),
    .X(_00427_));
 sky130_fd_sc_hd__or2_1 _14775_ (.A(net459),
    .B(net659),
    .X(_09130_));
 sky130_fd_sc_hd__o211a_1 _14776_ (.A1(\core.csr.instruction_memoryAddress[18] ),
    .A2(net588),
    .B1(_09130_),
    .C1(net1909),
    .X(_00428_));
 sky130_fd_sc_hd__or2_1 _14777_ (.A(net460),
    .B(net659),
    .X(_09131_));
 sky130_fd_sc_hd__o211a_1 _14778_ (.A1(\core.csr.instruction_memoryAddress[19] ),
    .A2(net588),
    .B1(_09131_),
    .C1(net1899),
    .X(_00429_));
 sky130_fd_sc_hd__or2_1 _14779_ (.A(net462),
    .B(net659),
    .X(_09132_));
 sky130_fd_sc_hd__o211a_1 _14780_ (.A1(\core.csr.instruction_memoryAddress[20] ),
    .A2(net588),
    .B1(_09132_),
    .C1(net1900),
    .X(_00430_));
 sky130_fd_sc_hd__or2_1 _14781_ (.A(net463),
    .B(net658),
    .X(_09133_));
 sky130_fd_sc_hd__o211a_1 _14782_ (.A1(\core.csr.instruction_memoryAddress[21] ),
    .A2(net587),
    .B1(_09133_),
    .C1(net1893),
    .X(_00431_));
 sky130_fd_sc_hd__or2_1 _14783_ (.A(net464),
    .B(net658),
    .X(_09134_));
 sky130_fd_sc_hd__o211a_1 _14784_ (.A1(\core.csr.instruction_memoryAddress[22] ),
    .A2(net587),
    .B1(_09134_),
    .C1(net1886),
    .X(_00432_));
 sky130_fd_sc_hd__or2_1 _14785_ (.A(net465),
    .B(net658),
    .X(_09135_));
 sky130_fd_sc_hd__o211a_1 _14786_ (.A1(\core.csr.instruction_memoryAddress[23] ),
    .A2(net587),
    .B1(_09135_),
    .C1(net1893),
    .X(_00433_));
 sky130_fd_sc_hd__or2_1 _14787_ (.A(net466),
    .B(net658),
    .X(_09136_));
 sky130_fd_sc_hd__o211a_1 _14788_ (.A1(\core.csr.instruction_memoryAddress[24] ),
    .A2(net587),
    .B1(_09136_),
    .C1(net1893),
    .X(_00434_));
 sky130_fd_sc_hd__or2_1 _14789_ (.A(net467),
    .B(net658),
    .X(_09137_));
 sky130_fd_sc_hd__o211a_1 _14790_ (.A1(\core.csr.instruction_memoryAddress[25] ),
    .A2(net587),
    .B1(_09137_),
    .C1(net1899),
    .X(_00435_));
 sky130_fd_sc_hd__or2_1 _14791_ (.A(net468),
    .B(net659),
    .X(_09138_));
 sky130_fd_sc_hd__o211a_1 _14792_ (.A1(\core.csr.instruction_memoryAddress[26] ),
    .A2(net588),
    .B1(_09138_),
    .C1(net1899),
    .X(_00436_));
 sky130_fd_sc_hd__or2_1 _14793_ (.A(net469),
    .B(net659),
    .X(_09139_));
 sky130_fd_sc_hd__o211a_1 _14794_ (.A1(\core.csr.instruction_memoryAddress[27] ),
    .A2(net588),
    .B1(_09139_),
    .C1(net1899),
    .X(_00437_));
 sky130_fd_sc_hd__or2_1 _14795_ (.A(net470),
    .B(net658),
    .X(_09140_));
 sky130_fd_sc_hd__o211a_1 _14796_ (.A1(\core.csr.instruction_memoryAddress[28] ),
    .A2(net587),
    .B1(_09140_),
    .C1(net1887),
    .X(_00438_));
 sky130_fd_sc_hd__or2_1 _14797_ (.A(net471),
    .B(net659),
    .X(_09141_));
 sky130_fd_sc_hd__o211a_1 _14798_ (.A1(\core.csr.instruction_memoryAddress[29] ),
    .A2(net588),
    .B1(_09141_),
    .C1(net1891),
    .X(_00439_));
 sky130_fd_sc_hd__or2_1 _14799_ (.A(net473),
    .B(net658),
    .X(_09142_));
 sky130_fd_sc_hd__o211a_1 _14800_ (.A1(\core.csr.instruction_memoryAddress[30] ),
    .A2(net587),
    .B1(_09142_),
    .C1(net1887),
    .X(_00440_));
 sky130_fd_sc_hd__or2_1 _14801_ (.A(net474),
    .B(net658),
    .X(_09143_));
 sky130_fd_sc_hd__o211a_1 _14802_ (.A1(\core.csr.instruction_memoryAddress[31] ),
    .A2(net587),
    .B1(_09143_),
    .C1(net1889),
    .X(_00441_));
 sky130_fd_sc_hd__o21ai_1 _14803_ (.A1(net800),
    .A2(_07391_),
    .B1(net1773),
    .Y(_09144_));
 sky130_fd_sc_hd__o211a_1 _14804_ (.A1(\core.cancelStall ),
    .A2(net1773),
    .B1(net1908),
    .C1(_09144_),
    .X(_00442_));
 sky130_fd_sc_hd__and2_2 _14805_ (.A(net1326),
    .B(_07413_),
    .X(_09145_));
 sky130_fd_sc_hd__nand2_2 _14806_ (.A(net1327),
    .B(_07413_),
    .Y(_09146_));
 sky130_fd_sc_hd__and3_1 _14807_ (.A(net1326),
    .B(_07413_),
    .C(_07415_),
    .X(_09147_));
 sky130_fd_sc_hd__nand2_2 _14808_ (.A(_07415_),
    .B(_09145_),
    .Y(_09148_));
 sky130_fd_sc_hd__nand2_1 _14809_ (.A(_07491_),
    .B(net1174),
    .Y(_09149_));
 sky130_fd_sc_hd__o211a_4 _14810_ (.A1(_07494_),
    .A2(_09149_),
    .B1(net697),
    .C1(_08639_),
    .X(_09150_));
 sky130_fd_sc_hd__mux2_1 _14811_ (.A0(_05108_),
    .A1(_06639_),
    .S(net1308),
    .X(_09151_));
 sky130_fd_sc_hd__mux2_1 _14812_ (.A0(_05023_),
    .A1(_06562_),
    .S(net1308),
    .X(_09152_));
 sky130_fd_sc_hd__mux2_1 _14813_ (.A0(_09151_),
    .A1(_09152_),
    .S(net932),
    .X(_09153_));
 sky130_fd_sc_hd__mux2_1 _14814_ (.A0(_05187_),
    .A1(_06484_),
    .S(net1308),
    .X(_09154_));
 sky130_fd_sc_hd__mux2_1 _14815_ (.A0(_05276_),
    .A1(_06406_),
    .S(net1308),
    .X(_09155_));
 sky130_fd_sc_hd__mux2_1 _14816_ (.A0(_09154_),
    .A1(_09155_),
    .S(net932),
    .X(_09156_));
 sky130_fd_sc_hd__mux2_1 _14817_ (.A0(_09153_),
    .A1(_09156_),
    .S(net935),
    .X(_09157_));
 sky130_fd_sc_hd__mux2_1 _14818_ (.A0(_04771_),
    .A1(_05549_),
    .S(net1315),
    .X(_09158_));
 sky130_fd_sc_hd__mux2_1 _14819_ (.A0(_04693_),
    .A1(_06311_),
    .S(net1315),
    .X(_09159_));
 sky130_fd_sc_hd__mux2_1 _14820_ (.A0(_09158_),
    .A1(_09159_),
    .S(net934),
    .X(_09160_));
 sky130_fd_sc_hd__mux2_1 _14821_ (.A0(_04927_),
    .A1(_05331_),
    .S(net1315),
    .X(_09161_));
 sky130_fd_sc_hd__mux2_1 _14822_ (.A0(_04850_),
    .A1(_05452_),
    .S(net1315),
    .X(_09162_));
 sky130_fd_sc_hd__mux2_1 _14823_ (.A0(_09161_),
    .A1(_09162_),
    .S(net934),
    .X(_09163_));
 sky130_fd_sc_hd__mux2_1 _14824_ (.A0(_09160_),
    .A1(_09163_),
    .S(net935),
    .X(_09164_));
 sky130_fd_sc_hd__mux2_1 _14825_ (.A0(_09164_),
    .A1(_09157_),
    .S(net940),
    .X(_09165_));
 sky130_fd_sc_hd__mux2_1 _14826_ (.A0(_05795_),
    .A1(_07021_),
    .S(net1312),
    .X(_09166_));
 sky130_fd_sc_hd__mux2_1 _14827_ (.A0(_05880_),
    .A1(_06945_),
    .S(net1311),
    .X(_09167_));
 sky130_fd_sc_hd__mux2_1 _14828_ (.A0(_09166_),
    .A1(_09167_),
    .S(net933),
    .X(_09168_));
 sky130_fd_sc_hd__mux2_1 _14829_ (.A0(_05629_),
    .A1(_06788_),
    .S(net1310),
    .X(_09169_));
 sky130_fd_sc_hd__mux2_1 _14830_ (.A0(_05710_),
    .A1(_06866_),
    .S(net1310),
    .X(_09170_));
 sky130_fd_sc_hd__mux2_1 _14831_ (.A0(_09169_),
    .A1(_09170_),
    .S(net933),
    .X(_09171_));
 sky130_fd_sc_hd__mux2_1 _14832_ (.A0(_09168_),
    .A1(_09171_),
    .S(net936),
    .X(_09172_));
 sky130_fd_sc_hd__mux2_1 _14833_ (.A0(_05964_),
    .A1(_07108_),
    .S(net1311),
    .X(_09173_));
 sky130_fd_sc_hd__mux2_1 _14834_ (.A0(_06048_),
    .A1(_07191_),
    .S(net1311),
    .X(_09174_));
 sky130_fd_sc_hd__mux2_1 _14835_ (.A0(_09173_),
    .A1(_09174_),
    .S(net933),
    .X(_09175_));
 sky130_fd_sc_hd__mux2_1 _14836_ (.A0(_06227_),
    .A1(_07275_),
    .S(net1312),
    .X(_09176_));
 sky130_fd_sc_hd__mux2_1 _14837_ (.A0(_06133_),
    .A1(_07347_),
    .S(net1311),
    .X(_09177_));
 sky130_fd_sc_hd__mux2_1 _14838_ (.A0(_09176_),
    .A1(_09177_),
    .S(_06196_),
    .X(_09178_));
 sky130_fd_sc_hd__mux2_1 _14839_ (.A0(_09175_),
    .A1(_09178_),
    .S(_06101_),
    .X(_09179_));
 sky130_fd_sc_hd__mux2_1 _14840_ (.A0(_09179_),
    .A1(_09172_),
    .S(net940),
    .X(_09180_));
 sky130_fd_sc_hd__mux2_1 _14841_ (.A0(_09165_),
    .A1(_09180_),
    .S(net886),
    .X(_09181_));
 sky130_fd_sc_hd__mux2_1 _14842_ (.A0(_04850_),
    .A1(_05452_),
    .S(net1310),
    .X(_09182_));
 sky130_fd_sc_hd__mux2_1 _14843_ (.A0(_04927_),
    .A1(_05331_),
    .S(net1309),
    .X(_09183_));
 sky130_fd_sc_hd__mux2_1 _14844_ (.A0(_09182_),
    .A1(_09183_),
    .S(net932),
    .X(_09184_));
 sky130_fd_sc_hd__mux2_1 _14845_ (.A0(_04693_),
    .A1(_06311_),
    .S(net1310),
    .X(_09185_));
 sky130_fd_sc_hd__mux2_1 _14846_ (.A0(_04771_),
    .A1(_05549_),
    .S(net1310),
    .X(_09186_));
 sky130_fd_sc_hd__mux2_1 _14847_ (.A0(_09185_),
    .A1(_09186_),
    .S(net932),
    .X(_09187_));
 sky130_fd_sc_hd__mux2_1 _14848_ (.A0(_09184_),
    .A1(_09187_),
    .S(net936),
    .X(_09188_));
 sky130_fd_sc_hd__mux2_1 _14849_ (.A0(_05276_),
    .A1(_06406_),
    .S(net1313),
    .X(_09189_));
 sky130_fd_sc_hd__mux2_1 _14850_ (.A0(_05187_),
    .A1(_06484_),
    .S(net1313),
    .X(_09190_));
 sky130_fd_sc_hd__mux2_1 _14851_ (.A0(_09189_),
    .A1(_09190_),
    .S(net932),
    .X(_09191_));
 sky130_fd_sc_hd__mux2_1 _14852_ (.A0(_05023_),
    .A1(_06562_),
    .S(_07386_),
    .X(_09192_));
 sky130_fd_sc_hd__mux2_1 _14853_ (.A0(_05108_),
    .A1(_06639_),
    .S(_07386_),
    .X(_09193_));
 sky130_fd_sc_hd__mux2_1 _14854_ (.A0(_09192_),
    .A1(_09193_),
    .S(net932),
    .X(_09194_));
 sky130_fd_sc_hd__mux2_1 _14855_ (.A0(_09191_),
    .A1(_09194_),
    .S(net935),
    .X(_09195_));
 sky130_fd_sc_hd__mux2_1 _14856_ (.A0(_09195_),
    .A1(_09188_),
    .S(net940),
    .X(_09196_));
 sky130_fd_sc_hd__mux2_1 _14857_ (.A0(_05710_),
    .A1(_06866_),
    .S(net1314),
    .X(_09197_));
 sky130_fd_sc_hd__mux2_1 _14858_ (.A0(_05629_),
    .A1(_06788_),
    .S(net1314),
    .X(_09198_));
 sky130_fd_sc_hd__mux2_1 _14859_ (.A0(_09197_),
    .A1(_09198_),
    .S(net933),
    .X(_09199_));
 sky130_fd_sc_hd__mux2_1 _14860_ (.A0(_05879_),
    .A1(_06946_),
    .S(net1314),
    .X(_09200_));
 sky130_fd_sc_hd__mux2_2 _14861_ (.A0(_05795_),
    .A1(_07021_),
    .S(net1314),
    .X(_09201_));
 sky130_fd_sc_hd__inv_2 _14862_ (.A(_09201_),
    .Y(_09202_));
 sky130_fd_sc_hd__mux2_1 _14863_ (.A0(_09200_),
    .A1(_09202_),
    .S(net933),
    .X(_09203_));
 sky130_fd_sc_hd__inv_2 _14864_ (.A(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__mux2_1 _14865_ (.A0(_09199_),
    .A1(_09204_),
    .S(net936),
    .X(_09205_));
 sky130_fd_sc_hd__mux2_1 _14866_ (.A0(_06133_),
    .A1(_07347_),
    .S(net1314),
    .X(_09206_));
 sky130_fd_sc_hd__mux2_1 _14867_ (.A0(_06227_),
    .A1(_07275_),
    .S(net1314),
    .X(_09207_));
 sky130_fd_sc_hd__mux2_1 _14868_ (.A0(_09206_),
    .A1(_09207_),
    .S(net931),
    .X(_09208_));
 sky130_fd_sc_hd__mux2_1 _14869_ (.A0(_06047_),
    .A1(_07192_),
    .S(net1314),
    .X(_09209_));
 sky130_fd_sc_hd__mux2_1 _14870_ (.A0(_05963_),
    .A1(_07109_),
    .S(net1314),
    .X(_09210_));
 sky130_fd_sc_hd__mux2_1 _14871_ (.A0(_09209_),
    .A1(_09210_),
    .S(net933),
    .X(_09211_));
 sky130_fd_sc_hd__inv_2 _14872_ (.A(_09211_),
    .Y(_09212_));
 sky130_fd_sc_hd__mux2_1 _14873_ (.A0(_09208_),
    .A1(_09212_),
    .S(net885),
    .X(_09213_));
 sky130_fd_sc_hd__mux2_1 _14874_ (.A0(_09205_),
    .A1(_09213_),
    .S(net939),
    .X(_09214_));
 sky130_fd_sc_hd__mux2_1 _14875_ (.A0(_09196_),
    .A1(_09214_),
    .S(net944),
    .X(_09215_));
 sky130_fd_sc_hd__mux2_2 _14876_ (.A0(_09181_),
    .A1(_09215_),
    .S(net948),
    .X(_09216_));
 sky130_fd_sc_hd__and2_1 _14877_ (.A(_07374_),
    .B(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__nand2_1 _14878_ (.A(_06696_),
    .B(net1319),
    .Y(_09218_));
 sky130_fd_sc_hd__o31a_1 _14879_ (.A1(_04469_),
    .A2(_04475_),
    .A3(_04477_),
    .B1(_07488_),
    .X(_09219_));
 sky130_fd_sc_hd__nor2_1 _14880_ (.A(_04474_),
    .B(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__or2_1 _14881_ (.A(_04474_),
    .B(_09219_),
    .X(_09221_));
 sky130_fd_sc_hd__and3_4 _14882_ (.A(_07275_),
    .B(net1310),
    .C(net1014),
    .X(_09222_));
 sky130_fd_sc_hd__inv_2 _14883_ (.A(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__or2_2 _14884_ (.A(net947),
    .B(_09222_),
    .X(_09224_));
 sky130_fd_sc_hd__or2_4 _14885_ (.A(net945),
    .B(_09222_),
    .X(_09225_));
 sky130_fd_sc_hd__o21a_1 _14886_ (.A1(_06196_),
    .A2(net1014),
    .B1(_09176_),
    .X(_09226_));
 sky130_fd_sc_hd__mux2_1 _14887_ (.A0(_09222_),
    .A1(_09226_),
    .S(net936),
    .X(_09227_));
 sky130_fd_sc_hd__mux2_1 _14888_ (.A0(_09222_),
    .A1(_09227_),
    .S(net939),
    .X(_09228_));
 sky130_fd_sc_hd__o21a_2 _14889_ (.A1(net886),
    .A2(_09228_),
    .B1(_09225_),
    .X(_09229_));
 sky130_fd_sc_hd__o21ai_4 _14890_ (.A1(net950),
    .A2(_09229_),
    .B1(net825),
    .Y(_09230_));
 sky130_fd_sc_hd__o221a_1 _14891_ (.A1(_06695_),
    .A2(_07379_),
    .B1(net1308),
    .B2(_09230_),
    .C1(_09218_),
    .X(_09231_));
 sky130_fd_sc_hd__a32o_1 _14892_ (.A1(_04423_),
    .A2(_07361_),
    .A3(_07377_),
    .B1(_07373_),
    .B2(_04465_),
    .X(_09232_));
 sky130_fd_sc_hd__or3b_4 _14893_ (.A(_09232_),
    .B(_09217_),
    .C_N(_09231_),
    .X(_09233_));
 sky130_fd_sc_hd__nor2_4 _14894_ (.A(_04423_),
    .B(_09146_),
    .Y(_09234_));
 sky130_fd_sc_hd__nand2_1 _14895_ (.A(net1878),
    .B(_09145_),
    .Y(_09235_));
 sky130_fd_sc_hd__mux2_1 _14896_ (.A0(net1377),
    .A1(_06225_),
    .S(net1172),
    .X(_09236_));
 sky130_fd_sc_hd__nor2_2 _14897_ (.A(_04477_),
    .B(_09146_),
    .Y(_09237_));
 sky130_fd_sc_hd__nand2_1 _14898_ (.A(_04476_),
    .B(_09145_),
    .Y(_09238_));
 sky130_fd_sc_hd__nand2_1 _14899_ (.A(_07845_),
    .B(_07847_),
    .Y(_09239_));
 sky130_fd_sc_hd__a21o_2 _14900_ (.A1(_07863_),
    .A2(_07867_),
    .B1(net1789),
    .X(_09240_));
 sky130_fd_sc_hd__nor2_1 _14901_ (.A(_09239_),
    .B(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__or2_1 _14902_ (.A(_09239_),
    .B(_09240_),
    .X(_09242_));
 sky130_fd_sc_hd__a31oi_4 _14903_ (.A1(net1791),
    .A2(net1775),
    .A3(net1215),
    .B1(net1034),
    .Y(_09243_));
 sky130_fd_sc_hd__a31o_4 _14904_ (.A1(net1791),
    .A2(net1775),
    .A3(net1215),
    .B1(net1033),
    .X(_09244_));
 sky130_fd_sc_hd__mux2_1 _14905_ (.A0(_07851_),
    .A1(\core.pipe0_currentInstruction[28] ),
    .S(net1794),
    .X(_09245_));
 sky130_fd_sc_hd__and2b_1 _14906_ (.A_N(net1794),
    .B(_07850_),
    .X(_09246_));
 sky130_fd_sc_hd__a21o_1 _14907_ (.A1(net1794),
    .A2(\core.pipe0_currentInstruction[29] ),
    .B1(_09246_),
    .X(_09247_));
 sky130_fd_sc_hd__mux2_2 _14908_ (.A0(_07849_),
    .A1(\core.pipe0_currentInstruction[26] ),
    .S(net1793),
    .X(_09248_));
 sky130_fd_sc_hd__inv_2 _14909_ (.A(_09248_),
    .Y(_09249_));
 sky130_fd_sc_hd__or3_1 _14910_ (.A(_09245_),
    .B(_09247_),
    .C(_09248_),
    .X(_09250_));
 sky130_fd_sc_hd__mux2_2 _14911_ (.A0(_07848_),
    .A1(net1816),
    .S(net1793),
    .X(_09251_));
 sky130_fd_sc_hd__and2b_1 _14912_ (.A_N(net1794),
    .B(_07854_),
    .X(_09252_));
 sky130_fd_sc_hd__a21o_1 _14913_ (.A1(net1794),
    .A2(net1818),
    .B1(_09252_),
    .X(_09253_));
 sky130_fd_sc_hd__nand2_4 _14914_ (.A(_09251_),
    .B(_09253_),
    .Y(_09254_));
 sky130_fd_sc_hd__and2b_1 _14915_ (.A_N(net1792),
    .B(_07853_),
    .X(_09255_));
 sky130_fd_sc_hd__a21o_1 _14916_ (.A1(net1793),
    .A2(net1822),
    .B1(_09255_),
    .X(_09256_));
 sky130_fd_sc_hd__nor2_1 _14917_ (.A(net1793),
    .B(_07844_),
    .Y(_09257_));
 sky130_fd_sc_hd__a21o_2 _14918_ (.A1(net1793),
    .A2(net1752),
    .B1(_09257_),
    .X(_09258_));
 sky130_fd_sc_hd__nand2b_1 _14919_ (.A_N(_09256_),
    .B(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__or3_2 _14920_ (.A(_09250_),
    .B(_09254_),
    .C(_09259_),
    .X(_09260_));
 sky130_fd_sc_hd__and2b_1 _14921_ (.A_N(net1792),
    .B(_07852_),
    .X(_09261_));
 sky130_fd_sc_hd__a21o_4 _14922_ (.A1(net1793),
    .A2(\core.pipe0_currentInstruction[27] ),
    .B1(_09261_),
    .X(_09262_));
 sky130_fd_sc_hd__or2_4 _14923_ (.A(_09260_),
    .B(_09262_),
    .X(_09263_));
 sky130_fd_sc_hd__and2b_2 _14924_ (.A_N(net1790),
    .B(_07869_),
    .X(_09264_));
 sky130_fd_sc_hd__a21o_2 _14925_ (.A1(net1792),
    .A2(net1831),
    .B1(_09264_),
    .X(_09265_));
 sky130_fd_sc_hd__mux2_4 _14926_ (.A0(_07870_),
    .A1(net1837),
    .S(net1792),
    .X(_09266_));
 sky130_fd_sc_hd__nor2_8 _14927_ (.A(_09265_),
    .B(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__mux2_8 _14928_ (.A0(_07843_),
    .A1(net1849),
    .S(net1792),
    .X(_09268_));
 sky130_fd_sc_hd__inv_2 _14929_ (.A(_09268_),
    .Y(_09269_));
 sky130_fd_sc_hd__mux2_4 _14930_ (.A0(_07876_),
    .A1(net1851),
    .S(net1792),
    .X(_09270_));
 sky130_fd_sc_hd__nor2_4 _14931_ (.A(_09268_),
    .B(net1166),
    .Y(_09271_));
 sky130_fd_sc_hd__nand2_8 _14932_ (.A(_09267_),
    .B(_09271_),
    .Y(_09272_));
 sky130_fd_sc_hd__nor2_8 _14933_ (.A(_09263_),
    .B(_09272_),
    .Y(_09273_));
 sky130_fd_sc_hd__nand2b_4 _14934_ (.A_N(_09260_),
    .B(_09262_),
    .Y(_09274_));
 sky130_fd_sc_hd__nor2_8 _14935_ (.A(_09272_),
    .B(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__a22oi_2 _14936_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[32] ),
    .Y(_09276_));
 sky130_fd_sc_hd__and3_1 _14937_ (.A(net1004),
    .B(_09269_),
    .C(net1166),
    .X(_09277_));
 sky130_fd_sc_hd__nand2_2 _14938_ (.A(_09267_),
    .B(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__nor2_1 _14939_ (.A(_09263_),
    .B(net922),
    .Y(_09279_));
 sky130_fd_sc_hd__or2_4 _14940_ (.A(_09263_),
    .B(net922),
    .X(_09280_));
 sky130_fd_sc_hd__or3_4 _14941_ (.A(net1007),
    .B(_09260_),
    .C(_09272_),
    .X(_09281_));
 sky130_fd_sc_hd__nand2_4 _14942_ (.A(_09267_),
    .B(_09268_),
    .Y(_09282_));
 sky130_fd_sc_hd__nor2_2 _14943_ (.A(net1166),
    .B(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__or2_2 _14944_ (.A(net1166),
    .B(_09282_),
    .X(_09284_));
 sky130_fd_sc_hd__nor2_2 _14945_ (.A(_09263_),
    .B(_09284_),
    .Y(_09285_));
 sky130_fd_sc_hd__nor2_2 _14946_ (.A(_09274_),
    .B(_09284_),
    .Y(_09286_));
 sky130_fd_sc_hd__a22o_1 _14947_ (.A1(\core.csr.instretTimer.currentValue[0] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[32] ),
    .X(_09287_));
 sky130_fd_sc_hd__nor2_8 _14948_ (.A(_09274_),
    .B(net922),
    .Y(_09288_));
 sky130_fd_sc_hd__a221o_2 _14949_ (.A1(net1004),
    .A2(_09287_),
    .B1(net876),
    .B2(\core.csr.cycleTimer.currentValue[32] ),
    .C1(net884),
    .X(_09289_));
 sky130_fd_sc_hd__nand2_1 _14950_ (.A(_09245_),
    .B(_09247_),
    .Y(_09290_));
 sky130_fd_sc_hd__or4_2 _14951_ (.A(_09251_),
    .B(_09253_),
    .C(_09259_),
    .D(_09290_),
    .X(_09291_));
 sky130_fd_sc_hd__or3_4 _14952_ (.A(_09249_),
    .B(_09262_),
    .C(_09291_),
    .X(_09292_));
 sky130_fd_sc_hd__nor2_2 _14953_ (.A(net1007),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__and2_1 _14954_ (.A(_09283_),
    .B(_09293_),
    .X(_09294_));
 sky130_fd_sc_hd__and3_2 _14955_ (.A(_09267_),
    .B(_09268_),
    .C(net1166),
    .X(_09295_));
 sky130_fd_sc_hd__inv_2 _14956_ (.A(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__and2_1 _14957_ (.A(_09293_),
    .B(_09295_),
    .X(_09297_));
 sky130_fd_sc_hd__or3_1 _14958_ (.A(_09249_),
    .B(_09262_),
    .C(_09291_),
    .X(_09298_));
 sky130_fd_sc_hd__nor2_1 _14959_ (.A(net1007),
    .B(_09298_),
    .Y(_09299_));
 sky130_fd_sc_hd__and2b_1 _14960_ (.A_N(_09265_),
    .B(_09266_),
    .X(_09300_));
 sky130_fd_sc_hd__and2_4 _14961_ (.A(_09271_),
    .B(_09300_),
    .X(_09301_));
 sky130_fd_sc_hd__o21a_1 _14962_ (.A1(_09295_),
    .A2(_09301_),
    .B1(_09293_),
    .X(_09302_));
 sky130_fd_sc_hd__nor2_1 _14963_ (.A(net922),
    .B(_09292_),
    .Y(_09303_));
 sky130_fd_sc_hd__or2_2 _14964_ (.A(net922),
    .B(_09292_),
    .X(_09304_));
 sky130_fd_sc_hd__and3_1 _14965_ (.A(_09267_),
    .B(_09271_),
    .C(_09293_),
    .X(_09305_));
 sky130_fd_sc_hd__or3_4 _14966_ (.A(_09248_),
    .B(_09262_),
    .C(_09291_),
    .X(_09306_));
 sky130_fd_sc_hd__nand2_2 _14967_ (.A(_09277_),
    .B(_09300_),
    .Y(_09307_));
 sky130_fd_sc_hd__nor2_2 _14968_ (.A(_09306_),
    .B(_09307_),
    .Y(_09308_));
 sky130_fd_sc_hd__and3b_1 _14969_ (.A_N(_09306_),
    .B(net1004),
    .C(_09301_),
    .X(_09309_));
 sky130_fd_sc_hd__nor3_1 _14970_ (.A(net1007),
    .B(_09272_),
    .C(_09306_),
    .Y(_09310_));
 sky130_fd_sc_hd__or3_1 _14971_ (.A(net872),
    .B(_09309_),
    .C(_09310_),
    .X(_09311_));
 sky130_fd_sc_hd__or3_1 _14972_ (.A(_09302_),
    .B(_09308_),
    .C(_09311_),
    .X(_09312_));
 sky130_fd_sc_hd__or3_1 _14973_ (.A(_09248_),
    .B(_09262_),
    .C(_09290_),
    .X(_09313_));
 sky130_fd_sc_hd__or4_4 _14974_ (.A(_09254_),
    .B(_09256_),
    .C(_09258_),
    .D(_09313_),
    .X(_09314_));
 sky130_fd_sc_hd__nor2_1 _14975_ (.A(_09307_),
    .B(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__nor2_2 _14976_ (.A(net1007),
    .B(_09314_),
    .Y(_09316_));
 sky130_fd_sc_hd__inv_2 _14977_ (.A(_09316_),
    .Y(_09317_));
 sky130_fd_sc_hd__nand2_1 _14978_ (.A(_09301_),
    .B(_09316_),
    .Y(_09318_));
 sky130_fd_sc_hd__nor2_1 _14979_ (.A(net922),
    .B(_09314_),
    .Y(_09319_));
 sky130_fd_sc_hd__or3_1 _14980_ (.A(net1007),
    .B(_09260_),
    .C(_09284_),
    .X(_09320_));
 sky130_fd_sc_hd__or2_2 _14981_ (.A(_09256_),
    .B(_09313_),
    .X(_09321_));
 sky130_fd_sc_hd__or3_4 _14982_ (.A(_09254_),
    .B(_09258_),
    .C(_09321_),
    .X(_09322_));
 sky130_fd_sc_hd__nor2_1 _14983_ (.A(net922),
    .B(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__or2_2 _14984_ (.A(net1007),
    .B(_09322_),
    .X(_09324_));
 sky130_fd_sc_hd__inv_2 _14985_ (.A(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__and3_1 _14986_ (.A(net264),
    .B(_09283_),
    .C(_09325_),
    .X(_09326_));
 sky130_fd_sc_hd__nor2_1 _14987_ (.A(_09307_),
    .B(_09322_),
    .Y(_09327_));
 sky130_fd_sc_hd__nor2_1 _14988_ (.A(_09282_),
    .B(_09324_),
    .Y(_09328_));
 sky130_fd_sc_hd__a31o_1 _14989_ (.A1(net1),
    .A2(_09301_),
    .A3(_09325_),
    .B1(_09328_),
    .X(_09329_));
 sky130_fd_sc_hd__nand2_1 _14990_ (.A(_09283_),
    .B(_09299_),
    .Y(_09330_));
 sky130_fd_sc_hd__o21a_1 _14991_ (.A1(_09295_),
    .A2(_09301_),
    .B1(_09299_),
    .X(_09331_));
 sky130_fd_sc_hd__o221a_1 _14992_ (.A1(\core.csr.traps.mtval.csrReadData[0] ),
    .A2(_09296_),
    .B1(net868),
    .B2(\core.csr.traps.mip.csrReadData[0] ),
    .C1(_09331_),
    .X(_09332_));
 sky130_fd_sc_hd__mux2_1 _14993_ (.A0(\core.csr.traps.mcause.csrReadData[0] ),
    .A1(_09332_),
    .S(_09330_),
    .X(_09333_));
 sky130_fd_sc_hd__nand2_4 _14994_ (.A(net1004),
    .B(_09301_),
    .Y(_09334_));
 sky130_fd_sc_hd__nor2_1 _14995_ (.A(_09306_),
    .B(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__or2_4 _14996_ (.A(_09306_),
    .B(_09334_),
    .X(_09336_));
 sky130_fd_sc_hd__and3_1 _14997_ (.A(_09267_),
    .B(_09271_),
    .C(_09299_),
    .X(_09337_));
 sky130_fd_sc_hd__a221o_1 _14998_ (.A1(\core.csr.traps.mtvec.csrReadData[0] ),
    .A2(_09308_),
    .B1(_09337_),
    .B2(\core.csr.traps.mscratch.currentValue[0] ),
    .C1(net913),
    .X(_09338_));
 sky130_fd_sc_hd__or3_1 _14999_ (.A(net1007),
    .B(_09272_),
    .C(_09306_),
    .X(_09339_));
 sky130_fd_sc_hd__a211o_1 _15000_ (.A1(_09283_),
    .A2(_09299_),
    .B1(_09308_),
    .C1(_09331_),
    .X(_09340_));
 sky130_fd_sc_hd__o21bai_1 _15001_ (.A1(net922),
    .A2(_09298_),
    .B1_N(_09337_),
    .Y(_09341_));
 sky130_fd_sc_hd__o31a_1 _15002_ (.A1(net913),
    .A2(_09340_),
    .A3(_09341_),
    .B1(_09339_),
    .X(_09342_));
 sky130_fd_sc_hd__o221a_1 _15003_ (.A1(\core.csr.traps.mie.currentValue[0] ),
    .A2(net910),
    .B1(_09338_),
    .B2(_09333_),
    .C1(_09342_),
    .X(_09343_));
 sky130_fd_sc_hd__a211o_1 _15004_ (.A1(\core.csr.mconfigptr.currentValue[0] ),
    .A2(_09327_),
    .B1(_09329_),
    .C1(_09343_),
    .X(_09344_));
 sky130_fd_sc_hd__a211o_1 _15005_ (.A1(net280),
    .A2(net1166),
    .B1(_09282_),
    .C1(_09324_),
    .X(_09345_));
 sky130_fd_sc_hd__a211o_1 _15006_ (.A1(_09344_),
    .A2(_09345_),
    .B1(_09323_),
    .C1(_09326_),
    .X(_09346_));
 sky130_fd_sc_hd__o311a_1 _15007_ (.A1(net253),
    .A2(net922),
    .A3(_09322_),
    .B1(_09346_),
    .C1(_09320_),
    .X(_09347_));
 sky130_fd_sc_hd__o221ai_4 _15008_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(net880),
    .B1(_09289_),
    .B2(_09347_),
    .C1(_09281_),
    .Y(_09348_));
 sky130_fd_sc_hd__o21a_4 _15009_ (.A1(_09243_),
    .A2(_09276_),
    .B1(_09348_),
    .X(_09349_));
 sky130_fd_sc_hd__nor3_4 _15010_ (.A(_09254_),
    .B(_09258_),
    .C(_09321_),
    .Y(_09350_));
 sky130_fd_sc_hd__nand2b_4 _15011_ (.A_N(_09278_),
    .B(_09350_),
    .Y(_09351_));
 sky130_fd_sc_hd__or3b_4 _15012_ (.A(net1007),
    .B(_09282_),
    .C_N(_09350_),
    .X(_09352_));
 sky130_fd_sc_hd__nor2_4 _15013_ (.A(net1166),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__and4_1 _15014_ (.A(net1004),
    .B(_09269_),
    .C(net1166),
    .D(_09300_),
    .X(_09354_));
 sky130_fd_sc_hd__and2_1 _15015_ (.A(_09350_),
    .B(_09354_),
    .X(_09355_));
 sky130_fd_sc_hd__inv_2 _15016_ (.A(net855),
    .Y(_09356_));
 sky130_fd_sc_hd__o21bai_4 _15017_ (.A1(_09292_),
    .A2(_09334_),
    .B1_N(net868),
    .Y(_09357_));
 sky130_fd_sc_hd__and2b_1 _15018_ (.A_N(_09306_),
    .B(_09354_),
    .X(_09358_));
 sky130_fd_sc_hd__nand3_2 _15019_ (.A(net1004),
    .B(_09267_),
    .C(_09271_),
    .Y(_09359_));
 sky130_fd_sc_hd__nor2_1 _15020_ (.A(_09292_),
    .B(_09359_),
    .Y(_09360_));
 sky130_fd_sc_hd__and3_4 _15021_ (.A(net1003),
    .B(_09301_),
    .C(_09350_),
    .X(_09361_));
 sky130_fd_sc_hd__or4_4 _15022_ (.A(_09254_),
    .B(_09258_),
    .C(_09321_),
    .D(_09334_),
    .X(_09362_));
 sky130_fd_sc_hd__o21ai_1 _15023_ (.A1(net1169),
    .A2(_09349_),
    .B1(_09236_),
    .Y(_09363_));
 sky130_fd_sc_hd__o21ai_4 _15024_ (.A1(net1881),
    .A2(_04463_),
    .B1(_04477_),
    .Y(_09364_));
 sky130_fd_sc_hd__and2_1 _15025_ (.A(_07377_),
    .B(_07413_),
    .X(_09365_));
 sky130_fd_sc_hd__nand2_4 _15026_ (.A(_07377_),
    .B(_07413_),
    .Y(_09366_));
 sky130_fd_sc_hd__a21oi_1 _15027_ (.A1(_09236_),
    .A2(net1211),
    .B1(_09364_),
    .Y(_09367_));
 sky130_fd_sc_hd__nor2_1 _15028_ (.A(net1174),
    .B(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__a22o_1 _15029_ (.A1(net1274),
    .A2(_06697_),
    .B1(_09363_),
    .B2(_09368_),
    .X(_09369_));
 sky130_fd_sc_hd__a211o_1 _15030_ (.A1(net1080),
    .A2(_09233_),
    .B1(_09369_),
    .C1(net1183),
    .X(_09370_));
 sky130_fd_sc_hd__o21a_1 _15031_ (.A1(net450),
    .A2(net1184),
    .B1(_09370_),
    .X(_09371_));
 sky130_fd_sc_hd__a21oi_1 _15032_ (.A1(_07368_),
    .A2(net1080),
    .B1(net1288),
    .Y(_09372_));
 sky130_fd_sc_hd__o21ai_1 _15033_ (.A1(net831),
    .A2(_09372_),
    .B1(_09150_),
    .Y(_09373_));
 sky130_fd_sc_hd__o221a_1 _15034_ (.A1(\core.pipe1_resultRegister[0] ),
    .A2(net655),
    .B1(_09371_),
    .B2(_09373_),
    .C1(net1921),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_2 _15035_ (.A0(_09185_),
    .A1(_09198_),
    .S(_06196_),
    .X(_09374_));
 sky130_fd_sc_hd__mux2_1 _15036_ (.A0(_09197_),
    .A1(_09201_),
    .S(net931),
    .X(_09375_));
 sky130_fd_sc_hd__mux2_1 _15037_ (.A0(_09374_),
    .A1(_09375_),
    .S(net937),
    .X(_09376_));
 sky130_fd_sc_hd__mux2_1 _15038_ (.A0(_09200_),
    .A1(_09210_),
    .S(net931),
    .X(_09377_));
 sky130_fd_sc_hd__nor2_1 _15039_ (.A(net934),
    .B(_09206_),
    .Y(_09378_));
 sky130_fd_sc_hd__a211o_1 _15040_ (.A1(net934),
    .A2(_09209_),
    .B1(_09378_),
    .C1(net885),
    .X(_09379_));
 sky130_fd_sc_hd__o21ai_1 _15041_ (.A1(net937),
    .A2(_09377_),
    .B1(_09379_),
    .Y(_09380_));
 sky130_fd_sc_hd__mux2_1 _15042_ (.A0(_09376_),
    .A1(_09380_),
    .S(net942),
    .X(_09381_));
 sky130_fd_sc_hd__mux2_1 _15043_ (.A0(_09154_),
    .A1(_09190_),
    .S(net931),
    .X(_09382_));
 sky130_fd_sc_hd__mux2_1 _15044_ (.A0(_09189_),
    .A1(_09193_),
    .S(net931),
    .X(_09383_));
 sky130_fd_sc_hd__mux2_1 _15045_ (.A0(_09382_),
    .A1(_09383_),
    .S(net935),
    .X(_09384_));
 sky130_fd_sc_hd__mux2_1 _15046_ (.A0(_09183_),
    .A1(_09192_),
    .S(net932),
    .X(_09385_));
 sky130_fd_sc_hd__mux2_1 _15047_ (.A0(_09182_),
    .A1(_09186_),
    .S(net931),
    .X(_09386_));
 sky130_fd_sc_hd__mux2_1 _15048_ (.A0(_09385_),
    .A1(_09386_),
    .S(net936),
    .X(_09387_));
 sky130_fd_sc_hd__mux2_1 _15049_ (.A0(_09384_),
    .A1(_09387_),
    .S(net941),
    .X(_09388_));
 sky130_fd_sc_hd__mux2_1 _15050_ (.A0(_09381_),
    .A1(_09388_),
    .S(net887),
    .X(_09389_));
 sky130_fd_sc_hd__mux2_1 _15051_ (.A0(_09174_),
    .A1(_09177_),
    .S(net933),
    .X(_09390_));
 sky130_fd_sc_hd__mux2_1 _15052_ (.A0(_09226_),
    .A1(_09390_),
    .S(net937),
    .X(_09391_));
 sky130_fd_sc_hd__inv_2 _15053_ (.A(_09391_),
    .Y(_09392_));
 sky130_fd_sc_hd__mux2_1 _15054_ (.A0(_09167_),
    .A1(_09173_),
    .S(net933),
    .X(_09393_));
 sky130_fd_sc_hd__mux2_2 _15055_ (.A0(_09166_),
    .A1(_09170_),
    .S(net931),
    .X(_09394_));
 sky130_fd_sc_hd__mux2_1 _15056_ (.A0(_09393_),
    .A1(_09394_),
    .S(net937),
    .X(_09395_));
 sky130_fd_sc_hd__mux2_1 _15057_ (.A0(_09391_),
    .A1(_09395_),
    .S(net942),
    .X(_09396_));
 sky130_fd_sc_hd__mux2_1 _15058_ (.A0(_09152_),
    .A1(_09161_),
    .S(net932),
    .X(_09397_));
 sky130_fd_sc_hd__mux2_1 _15059_ (.A0(_09151_),
    .A1(_09155_),
    .S(net931),
    .X(_09398_));
 sky130_fd_sc_hd__mux2_1 _15060_ (.A0(_09397_),
    .A1(_09398_),
    .S(net935),
    .X(_09399_));
 sky130_fd_sc_hd__mux2_1 _15061_ (.A0(_09159_),
    .A1(_09169_),
    .S(net933),
    .X(_09400_));
 sky130_fd_sc_hd__mux2_2 _15062_ (.A0(_09158_),
    .A1(_09162_),
    .S(net931),
    .X(_09401_));
 sky130_fd_sc_hd__mux2_1 _15063_ (.A0(_09400_),
    .A1(_09401_),
    .S(net935),
    .X(_09402_));
 sky130_fd_sc_hd__mux2_1 _15064_ (.A0(_09402_),
    .A1(_09399_),
    .S(net941),
    .X(_09403_));
 sky130_fd_sc_hd__mux2_4 _15065_ (.A0(_09396_),
    .A1(_09403_),
    .S(net945),
    .X(_09404_));
 sky130_fd_sc_hd__mux2_4 _15066_ (.A0(_09389_),
    .A1(_09404_),
    .S(net949),
    .X(_09405_));
 sky130_fd_sc_hd__mux2_1 _15067_ (.A0(_09178_),
    .A1(_09222_),
    .S(_06101_),
    .X(_09406_));
 sky130_fd_sc_hd__mux2_1 _15068_ (.A0(_09222_),
    .A1(_09406_),
    .S(net942),
    .X(_09407_));
 sky130_fd_sc_hd__o21a_1 _15069_ (.A1(net886),
    .A2(_09407_),
    .B1(_09225_),
    .X(_09408_));
 sky130_fd_sc_hd__o21ai_4 _15070_ (.A1(net949),
    .A2(_09408_),
    .B1(net826),
    .Y(_09409_));
 sky130_fd_sc_hd__mux2_1 _15071_ (.A0(_07383_),
    .A1(net1322),
    .S(_06134_),
    .X(_09410_));
 sky130_fd_sc_hd__o22a_1 _15072_ (.A1(_06101_),
    .A2(_06133_),
    .B1(net1319),
    .B2(_09410_),
    .X(_09411_));
 sky130_fd_sc_hd__o21ai_1 _15073_ (.A1(net1310),
    .A2(_09409_),
    .B1(net1326),
    .Y(_09412_));
 sky130_fd_sc_hd__a211o_1 _15074_ (.A1(_07374_),
    .A2(_09405_),
    .B1(_09411_),
    .C1(_09412_),
    .X(_09413_));
 sky130_fd_sc_hd__nand2_1 _15075_ (.A(_06136_),
    .B(_06228_),
    .Y(_09414_));
 sky130_fd_sc_hd__nor2_1 _15076_ (.A(_07475_),
    .B(net1014),
    .Y(_09415_));
 sky130_fd_sc_hd__o211a_1 _15077_ (.A1(_06136_),
    .A2(_06228_),
    .B1(net1015),
    .C1(_09414_),
    .X(_09416_));
 sky130_fd_sc_hd__mux2_1 _15078_ (.A0(net1473),
    .A1(_06132_),
    .S(net1172),
    .X(_09417_));
 sky130_fd_sc_hd__a22o_1 _15079_ (.A1(\core.csr.cycleTimer.currentValue[1] ),
    .A2(net930),
    .B1(net926),
    .B2(\core.csr.cycleTimer.currentValue[33] ),
    .X(_09418_));
 sky130_fd_sc_hd__a22o_1 _15080_ (.A1(\core.csr.instretTimer.currentValue[1] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[33] ),
    .X(_09419_));
 sky130_fd_sc_hd__and2_1 _15081_ (.A(net281),
    .B(net1166),
    .X(_09420_));
 sky130_fd_sc_hd__mux2_1 _15082_ (.A0(\core.csr.traps.mip.csrReadData[1] ),
    .A1(\core.csr.traps.mtval.csrReadData[1] ),
    .S(net869),
    .X(_09421_));
 sky130_fd_sc_hd__a221o_1 _15083_ (.A1(\core.csr.traps.mcause.csrReadData[1] ),
    .A2(net872),
    .B1(net822),
    .B2(_09421_),
    .C1(net864),
    .X(_09422_));
 sky130_fd_sc_hd__o21a_1 _15084_ (.A1(\core.csr.trapReturnVector[1] ),
    .A2(net861),
    .B1(_09422_),
    .X(_09423_));
 sky130_fd_sc_hd__a221o_2 _15085_ (.A1(\core.csr.traps.mtvec.csrReadData[1] ),
    .A2(net905),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[1] ),
    .C1(_09423_),
    .X(_09424_));
 sky130_fd_sc_hd__mux2_1 _15086_ (.A0(\core.csr.traps.mie.currentValue[1] ),
    .A1(_09424_),
    .S(net909),
    .X(_09425_));
 sky130_fd_sc_hd__a221o_2 _15087_ (.A1(\core.csr.mconfigptr.currentValue[1] ),
    .A2(net855),
    .B1(_09361_),
    .B2(net2),
    .C1(_09425_),
    .X(_09426_));
 sky130_fd_sc_hd__mux2_1 _15088_ (.A0(_09420_),
    .A1(_09426_),
    .S(_09352_),
    .X(_09427_));
 sky130_fd_sc_hd__a21o_1 _15089_ (.A1(net271),
    .A2(net824),
    .B1(_09427_),
    .X(_09428_));
 sky130_fd_sc_hd__mux2_2 _15090_ (.A0(net255),
    .A1(_09428_),
    .S(_09351_),
    .X(_09429_));
 sky130_fd_sc_hd__a221o_1 _15091_ (.A1(\core.csr.cycleTimer.currentValue[33] ),
    .A2(net876),
    .B1(_09419_),
    .B2(net1004),
    .C1(_09429_),
    .X(_09430_));
 sky130_fd_sc_hd__mux2_2 _15092_ (.A0(\core.csr.cycleTimer.currentValue[1] ),
    .A1(_09430_),
    .S(net881),
    .X(_09431_));
 sky130_fd_sc_hd__a21oi_4 _15093_ (.A1(net1004),
    .A2(_09418_),
    .B1(_09431_),
    .Y(_09432_));
 sky130_fd_sc_hd__o21ai_1 _15094_ (.A1(net1169),
    .A2(_09432_),
    .B1(_09417_),
    .Y(_09433_));
 sky130_fd_sc_hd__and3_1 _15095_ (.A(net1326),
    .B(_07413_),
    .C(_09364_),
    .X(_09434_));
 sky130_fd_sc_hd__nand2_1 _15096_ (.A(_09145_),
    .B(_09364_),
    .Y(_09435_));
 sky130_fd_sc_hd__a21o_1 _15097_ (.A1(net1211),
    .A2(_09417_),
    .B1(net1208),
    .X(_09436_));
 sky130_fd_sc_hd__a32o_1 _15098_ (.A1(net1215),
    .A2(_09433_),
    .A3(_09436_),
    .B1(_07474_),
    .B2(net1274),
    .X(_09437_));
 sky130_fd_sc_hd__o31a_1 _15099_ (.A1(net1327),
    .A2(_09415_),
    .A3(_09416_),
    .B1(_09413_),
    .X(_09438_));
 sky130_fd_sc_hd__a21oi_1 _15100_ (.A1(net1080),
    .A2(_09438_),
    .B1(_09437_),
    .Y(_09439_));
 sky130_fd_sc_hd__o211a_1 _15101_ (.A1(net1184),
    .A2(_07405_),
    .B1(_09439_),
    .C1(net1284),
    .X(_09440_));
 sky130_fd_sc_hd__o21ai_1 _15102_ (.A1(_06102_),
    .A2(_09440_),
    .B1(net655),
    .Y(_09441_));
 sky130_fd_sc_hd__o211a_1 _15103_ (.A1(net1809),
    .A2(net655),
    .B1(_09441_),
    .C1(net1920),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _15104_ (.A0(_09168_),
    .A1(_09175_),
    .S(net885),
    .X(_09442_));
 sky130_fd_sc_hd__mux2_1 _15105_ (.A0(_09406_),
    .A1(_09442_),
    .S(net942),
    .X(_09443_));
 sky130_fd_sc_hd__mux2_1 _15106_ (.A0(_09153_),
    .A1(_09163_),
    .S(net885),
    .X(_09444_));
 sky130_fd_sc_hd__mux2_1 _15107_ (.A0(_09160_),
    .A1(_09171_),
    .S(net885),
    .X(_09445_));
 sky130_fd_sc_hd__mux2_1 _15108_ (.A0(_09445_),
    .A1(_09444_),
    .S(net941),
    .X(_09446_));
 sky130_fd_sc_hd__mux2_2 _15109_ (.A0(_09443_),
    .A1(_09446_),
    .S(net945),
    .X(_09447_));
 sky130_fd_sc_hd__mux2_1 _15110_ (.A0(_09184_),
    .A1(_09194_),
    .S(net885),
    .X(_09448_));
 sky130_fd_sc_hd__mux2_1 _15111_ (.A0(_09156_),
    .A1(_09191_),
    .S(net935),
    .X(_09449_));
 sky130_fd_sc_hd__mux2_1 _15112_ (.A0(_09449_),
    .A1(_09448_),
    .S(net941),
    .X(_09450_));
 sky130_fd_sc_hd__mux2_1 _15113_ (.A0(_09187_),
    .A1(_09199_),
    .S(net936),
    .X(_09451_));
 sky130_fd_sc_hd__nor2_1 _15114_ (.A(net937),
    .B(_09203_),
    .Y(_09452_));
 sky130_fd_sc_hd__o21ai_1 _15115_ (.A1(net885),
    .A2(_09211_),
    .B1(net942),
    .Y(_09453_));
 sky130_fd_sc_hd__o221a_1 _15116_ (.A1(net943),
    .A2(_09451_),
    .B1(_09452_),
    .B2(_09453_),
    .C1(net946),
    .X(_09454_));
 sky130_fd_sc_hd__a21o_1 _15117_ (.A1(net887),
    .A2(_09450_),
    .B1(_09454_),
    .X(_09455_));
 sky130_fd_sc_hd__mux2_4 _15118_ (.A0(_09447_),
    .A1(_09455_),
    .S(_05847_),
    .X(_09456_));
 sky130_fd_sc_hd__nand2_1 _15119_ (.A(_07374_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__mux2_1 _15120_ (.A0(_09223_),
    .A1(_09392_),
    .S(net942),
    .X(_09458_));
 sky130_fd_sc_hd__inv_2 _15121_ (.A(_09458_),
    .Y(_09459_));
 sky130_fd_sc_hd__o21ai_2 _15122_ (.A1(net887),
    .A2(_09459_),
    .B1(_09225_),
    .Y(_09460_));
 sky130_fd_sc_hd__a21bo_4 _15123_ (.A1(net947),
    .A2(_09460_),
    .B1_N(net826),
    .X(_09461_));
 sky130_fd_sc_hd__a21oi_1 _15124_ (.A1(_06050_),
    .A2(_07378_),
    .B1(net1330),
    .Y(_09462_));
 sky130_fd_sc_hd__o221a_1 _15125_ (.A1(_06053_),
    .A2(_07384_),
    .B1(net1311),
    .B2(_09461_),
    .C1(_09462_),
    .X(_09463_));
 sky130_fd_sc_hd__o211a_1 _15126_ (.A1(_06051_),
    .A2(_07381_),
    .B1(_09457_),
    .C1(_09463_),
    .X(_09464_));
 sky130_fd_sc_hd__nand2_1 _15127_ (.A(_08382_),
    .B(net1010),
    .Y(_09465_));
 sky130_fd_sc_hd__o211a_1 _15128_ (.A1(_06694_),
    .A2(net1010),
    .B1(_09465_),
    .C1(net1330),
    .X(_09466_));
 sky130_fd_sc_hd__mux2_1 _15129_ (.A0(net1439),
    .A1(_06046_),
    .S(net1172),
    .X(_09467_));
 sky130_fd_sc_hd__a22o_1 _15130_ (.A1(\core.csr.cycleTimer.currentValue[2] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[34] ),
    .X(_09468_));
 sky130_fd_sc_hd__a22o_1 _15131_ (.A1(\core.csr.instretTimer.currentValue[2] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[34] ),
    .X(_09469_));
 sky130_fd_sc_hd__mux2_1 _15132_ (.A0(\core.csr.traps.mip.csrReadData[2] ),
    .A1(\core.csr.traps.mtval.csrReadData[2] ),
    .S(net868),
    .X(_09470_));
 sky130_fd_sc_hd__and2_1 _15133_ (.A(net282),
    .B(net1166),
    .X(_09471_));
 sky130_fd_sc_hd__or2_4 _15134_ (.A(_09306_),
    .B(_09359_),
    .X(_09472_));
 sky130_fd_sc_hd__a221o_1 _15135_ (.A1(\core.csr.traps.mcause.csrReadData[2] ),
    .A2(net872),
    .B1(net822),
    .B2(_09470_),
    .C1(net864),
    .X(_09473_));
 sky130_fd_sc_hd__o21ba_1 _15136_ (.A1(\core.csr.trapReturnVector[2] ),
    .A2(net860),
    .B1_N(net902),
    .X(_09474_));
 sky130_fd_sc_hd__a221o_1 _15137_ (.A1(\core.csr.traps.mscratch.currentValue[2] ),
    .A2(net902),
    .B1(_09473_),
    .B2(_09474_),
    .C1(net905),
    .X(_09475_));
 sky130_fd_sc_hd__a21oi_1 _15138_ (.A1(_04394_),
    .A2(net905),
    .B1(net913),
    .Y(_09476_));
 sky130_fd_sc_hd__a22o_1 _15139_ (.A1(\core.csr.traps.mie.currentValue[2] ),
    .A2(net913),
    .B1(_09475_),
    .B2(_09476_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_4 _15140_ (.A0(\core.csr.traps.machineInterruptEnable ),
    .A1(_01961_),
    .S(_09472_),
    .X(_01962_));
 sky130_fd_sc_hd__a221o_1 _15141_ (.A1(\core.csr.mconfigptr.currentValue[2] ),
    .A2(net856),
    .B1(_09361_),
    .B2(net3),
    .C1(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _15142_ (.A0(_09471_),
    .A1(_01963_),
    .S(_09352_),
    .X(_01964_));
 sky130_fd_sc_hd__a21o_1 _15143_ (.A1(net272),
    .A2(net824),
    .B1(_01964_),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_2 _15144_ (.A0(net256),
    .A1(_01965_),
    .S(_09351_),
    .X(_01966_));
 sky130_fd_sc_hd__a221o_1 _15145_ (.A1(\core.csr.cycleTimer.currentValue[34] ),
    .A2(net876),
    .B1(_09469_),
    .B2(net1002),
    .C1(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_2 _15146_ (.A0(\core.csr.cycleTimer.currentValue[2] ),
    .A1(_01967_),
    .S(net880),
    .X(_01968_));
 sky130_fd_sc_hd__a21oi_4 _15147_ (.A1(net1002),
    .A2(_09468_),
    .B1(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__o21ai_2 _15148_ (.A1(net1170),
    .A2(_01969_),
    .B1(_09467_),
    .Y(_01970_));
 sky130_fd_sc_hd__a21o_1 _15149_ (.A1(net1211),
    .A2(_09467_),
    .B1(net1209),
    .X(_01971_));
 sky130_fd_sc_hd__a221o_2 _15150_ (.A1(_07399_),
    .A2(_07577_),
    .B1(_08382_),
    .B2(net1274),
    .C1(net1288),
    .X(_01972_));
 sky130_fd_sc_hd__a31oi_4 _15151_ (.A1(net1215),
    .A2(_01970_),
    .A3(_01971_),
    .B1(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__o31a_1 _15152_ (.A1(net1083),
    .A2(_09464_),
    .A3(_09466_),
    .B1(_01973_),
    .X(_01974_));
 sky130_fd_sc_hd__o21ai_1 _15153_ (.A1(_06016_),
    .A2(_01974_),
    .B1(net655),
    .Y(_01975_));
 sky130_fd_sc_hd__o211a_1 _15154_ (.A1(\core.pipe1_resultRegister[2] ),
    .A2(net655),
    .B1(_01975_),
    .C1(net1920),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _15155_ (.A0(_09390_),
    .A1(_09393_),
    .S(net937),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_2 _15156_ (.A0(_09227_),
    .A1(_01976_),
    .S(net939),
    .X(_01977_));
 sky130_fd_sc_hd__inv_2 _15157_ (.A(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__or2_1 _15158_ (.A(net885),
    .B(_09397_),
    .X(_01979_));
 sky130_fd_sc_hd__o21ai_1 _15159_ (.A1(net935),
    .A2(_09401_),
    .B1(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__mux2_1 _15160_ (.A0(_09394_),
    .A1(_09400_),
    .S(net935),
    .X(_01981_));
 sky130_fd_sc_hd__inv_2 _15161_ (.A(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__mux2_1 _15162_ (.A0(_01982_),
    .A1(_01980_),
    .S(net939),
    .X(_01983_));
 sky130_fd_sc_hd__inv_2 _15163_ (.A(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__mux2_2 _15164_ (.A0(_01978_),
    .A1(_01983_),
    .S(net944),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _15165_ (.A0(_09383_),
    .A1(_09385_),
    .S(net935),
    .X(_01986_));
 sky130_fd_sc_hd__inv_2 _15166_ (.A(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__mux2_1 _15167_ (.A0(_09382_),
    .A1(_09398_),
    .S(net885),
    .X(_01988_));
 sky130_fd_sc_hd__inv_2 _15168_ (.A(_01988_),
    .Y(_01989_));
 sky130_fd_sc_hd__mux2_1 _15169_ (.A0(_01988_),
    .A1(_01986_),
    .S(net939),
    .X(_01990_));
 sky130_fd_sc_hd__or2_1 _15170_ (.A(net936),
    .B(_09386_),
    .X(_01991_));
 sky130_fd_sc_hd__o21ai_1 _15171_ (.A1(net885),
    .A2(_09374_),
    .B1(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__or2_1 _15172_ (.A(net939),
    .B(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__o21ai_1 _15173_ (.A1(net937),
    .A2(_09375_),
    .B1(net942),
    .Y(_01994_));
 sky130_fd_sc_hd__a21o_1 _15174_ (.A1(net937),
    .A2(_09377_),
    .B1(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__nor2_1 _15175_ (.A(net944),
    .B(_01990_),
    .Y(_01996_));
 sky130_fd_sc_hd__a311o_1 _15176_ (.A1(net944),
    .A2(_01993_),
    .A3(_01995_),
    .B1(_01996_),
    .C1(net950),
    .X(_01997_));
 sky130_fd_sc_hd__o21a_1 _15177_ (.A1(net948),
    .A2(_01985_),
    .B1(_01997_),
    .X(_01998_));
 sky130_fd_sc_hd__o21ai_1 _15178_ (.A1(_05966_),
    .A2(_07384_),
    .B1(_07381_),
    .Y(_01999_));
 sky130_fd_sc_hd__a22o_1 _15179_ (.A1(_05966_),
    .A2(net1322),
    .B1(_01999_),
    .B2(_05967_),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _15180_ (.A0(_09222_),
    .A1(_09179_),
    .S(net940),
    .X(_02001_));
 sky130_fd_sc_hd__o21a_1 _15181_ (.A1(net886),
    .A2(_02001_),
    .B1(_09225_),
    .X(_02002_));
 sky130_fd_sc_hd__o21ai_1 _15182_ (.A1(net950),
    .A2(_02002_),
    .B1(net825),
    .Y(_02003_));
 sky130_fd_sc_hd__o22a_1 _15183_ (.A1(net1325),
    .A2(_01998_),
    .B1(_02003_),
    .B2(net1310),
    .X(_02004_));
 sky130_fd_sc_hd__and3b_1 _15184_ (.A_N(_02000_),
    .B(_02004_),
    .C(net1326),
    .X(_02005_));
 sky130_fd_sc_hd__or2_1 _15185_ (.A(_08394_),
    .B(net1015),
    .X(_02006_));
 sky130_fd_sc_hd__o211a_1 _15186_ (.A1(_06693_),
    .A2(net1010),
    .B1(_02006_),
    .C1(net1329),
    .X(_02007_));
 sky130_fd_sc_hd__or3_1 _15187_ (.A(net1083),
    .B(_02005_),
    .C(_02007_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _15188_ (.A0(net1492),
    .A1(_05962_),
    .S(net1172),
    .X(_02009_));
 sky130_fd_sc_hd__a22o_1 _15189_ (.A1(\core.csr.cycleTimer.currentValue[3] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[35] ),
    .X(_02010_));
 sky130_fd_sc_hd__a22o_1 _15190_ (.A1(\core.csr.instretTimer.currentValue[3] ),
    .A2(net919),
    .B1(net915),
    .B2(\core.csr.instretTimer.currentValue[35] ),
    .X(_02011_));
 sky130_fd_sc_hd__a21o_1 _15191_ (.A1(net283),
    .A2(_09270_),
    .B1(_09352_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _15192_ (.A0(\core.csr.traps.mip.csrReadData[3] ),
    .A1(\core.csr.traps.mtval.csrReadData[3] ),
    .S(net869),
    .X(_02013_));
 sky130_fd_sc_hd__a221o_1 _15193_ (.A1(\core.csr.traps.mcause.csrReadData[3] ),
    .A2(net872),
    .B1(net822),
    .B2(_02013_),
    .C1(net864),
    .X(_02014_));
 sky130_fd_sc_hd__o21a_1 _15194_ (.A1(\core.csr.trapReturnVector[3] ),
    .A2(net860),
    .B1(_02014_),
    .X(_02015_));
 sky130_fd_sc_hd__a221o_4 _15195_ (.A1(\core.csr.traps.mtvec.csrReadData[3] ),
    .A2(net905),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[3] ),
    .C1(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_1 _15196_ (.A0(\core.csr.traps.mie.currentValue[3] ),
    .A1(_02016_),
    .S(net910),
    .X(_02017_));
 sky130_fd_sc_hd__a32o_1 _15197_ (.A1(net1003),
    .A2(_09295_),
    .A3(_09350_),
    .B1(_09361_),
    .B2(net4),
    .X(_02018_));
 sky130_fd_sc_hd__a211o_2 _15198_ (.A1(\core.csr.mconfigptr.currentValue[3] ),
    .A2(net856),
    .B1(_02017_),
    .C1(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__a22o_1 _15199_ (.A1(net273),
    .A2(net824),
    .B1(_02012_),
    .B2(_02019_),
    .X(_02020_));
 sky130_fd_sc_hd__mux2_1 _15200_ (.A0(net257),
    .A1(_02020_),
    .S(_09351_),
    .X(_02021_));
 sky130_fd_sc_hd__a221o_1 _15201_ (.A1(\core.csr.cycleTimer.currentValue[35] ),
    .A2(net877),
    .B1(_02011_),
    .B2(net1002),
    .C1(_02021_),
    .X(_02022_));
 sky130_fd_sc_hd__mux2_2 _15202_ (.A0(\core.csr.cycleTimer.currentValue[3] ),
    .A1(_02022_),
    .S(net880),
    .X(_02023_));
 sky130_fd_sc_hd__a21oi_4 _15203_ (.A1(net1002),
    .A2(_02010_),
    .B1(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__o21ba_1 _15204_ (.A1(net1170),
    .A2(_02024_),
    .B1_N(_02009_),
    .X(_02025_));
 sky130_fd_sc_hd__o21a_1 _15205_ (.A1(_09366_),
    .A2(_02009_),
    .B1(net1165),
    .X(_02026_));
 sky130_fd_sc_hd__or3_1 _15206_ (.A(net1174),
    .B(_02025_),
    .C(_02026_),
    .X(_02027_));
 sky130_fd_sc_hd__o221a_1 _15207_ (.A1(net1185),
    .A2(_07568_),
    .B1(_08394_),
    .B2(_04480_),
    .C1(net1284),
    .X(_02028_));
 sky130_fd_sc_hd__and3_1 _15208_ (.A(_02008_),
    .B(_02027_),
    .C(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__o21ai_1 _15209_ (.A1(_05932_),
    .A2(_02029_),
    .B1(net656),
    .Y(_02030_));
 sky130_fd_sc_hd__o211a_1 _15210_ (.A1(\core.pipe1_resultRegister[3] ),
    .A2(net656),
    .B1(_02030_),
    .C1(net1926),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _15211_ (.A0(_09172_),
    .A1(_09164_),
    .S(net940),
    .X(_02031_));
 sky130_fd_sc_hd__mux2_4 _15212_ (.A0(_02001_),
    .A1(_02031_),
    .S(net945),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _15213_ (.A0(_09157_),
    .A1(_09195_),
    .S(net939),
    .X(_02033_));
 sky130_fd_sc_hd__or2_1 _15214_ (.A(net944),
    .B(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _15215_ (.A0(_09188_),
    .A1(_09205_),
    .S(net940),
    .X(_02035_));
 sky130_fd_sc_hd__o211a_1 _15216_ (.A1(net886),
    .A2(_02035_),
    .B1(_02034_),
    .C1(net948),
    .X(_02036_));
 sky130_fd_sc_hd__a21oi_4 _15217_ (.A1(net950),
    .A2(_02032_),
    .B1(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__or2_1 _15218_ (.A(net1324),
    .B(_02037_),
    .X(_02038_));
 sky130_fd_sc_hd__nor2_8 _15219_ (.A(net1326),
    .B(_07393_),
    .Y(_02039_));
 sky130_fd_sc_hd__or2_4 _15220_ (.A(net1326),
    .B(_07393_),
    .X(_02040_));
 sky130_fd_sc_hd__nor2_1 _15221_ (.A(_06692_),
    .B(net1011),
    .Y(_02041_));
 sky130_fd_sc_hd__a211o_1 _15222_ (.A1(_08421_),
    .A2(net1011),
    .B1(_02040_),
    .C1(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__o21a_2 _15223_ (.A1(net886),
    .A2(_01977_),
    .B1(_09225_),
    .X(_02043_));
 sky130_fd_sc_hd__o21ai_4 _15224_ (.A1(net950),
    .A2(_02043_),
    .B1(net825),
    .Y(_02044_));
 sky130_fd_sc_hd__a31o_1 _15225_ (.A1(_05846_),
    .A2(_05880_),
    .A3(net1322),
    .B1(net1319),
    .X(_02045_));
 sky130_fd_sc_hd__nand2_1 _15226_ (.A(_05882_),
    .B(_02045_),
    .Y(_02046_));
 sky130_fd_sc_hd__o221a_1 _15227_ (.A1(_05883_),
    .A2(_07384_),
    .B1(net1311),
    .B2(_02044_),
    .C1(_02042_),
    .X(_02047_));
 sky130_fd_sc_hd__a31o_1 _15228_ (.A1(_02038_),
    .A2(_02046_),
    .A3(_02047_),
    .B1(net1083),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _15229_ (.A0(_04645_),
    .A1(_05878_),
    .S(net1173),
    .X(_02049_));
 sky130_fd_sc_hd__a22o_1 _15230_ (.A1(\core.csr.cycleTimer.currentValue[4] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[36] ),
    .X(_02050_));
 sky130_fd_sc_hd__a22o_1 _15231_ (.A1(\core.csr.instretTimer.currentValue[4] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[36] ),
    .X(_02051_));
 sky130_fd_sc_hd__or2_1 _15232_ (.A(net5),
    .B(_09362_),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _15233_ (.A0(\core.csr.traps.mip.csrReadData[4] ),
    .A1(\core.csr.traps.mtval.csrReadData[4] ),
    .S(net869),
    .X(_02053_));
 sky130_fd_sc_hd__a221o_1 _15234_ (.A1(\core.csr.traps.mcause.csrReadData[4] ),
    .A2(net873),
    .B1(net823),
    .B2(_02053_),
    .C1(net864),
    .X(_02054_));
 sky130_fd_sc_hd__o21a_1 _15235_ (.A1(\core.csr.trapReturnVector[4] ),
    .A2(net860),
    .B1(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__a221o_1 _15236_ (.A1(\core.csr.traps.mtvec.csrReadData[4] ),
    .A2(net906),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[4] ),
    .C1(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _15237_ (.A0(\core.csr.traps.mie.currentValue[4] ),
    .A1(_02056_),
    .S(net910),
    .X(_02057_));
 sky130_fd_sc_hd__a211o_4 _15238_ (.A1(\core.csr.mconfigptr.currentValue[4] ),
    .A2(net855),
    .B1(_09361_),
    .C1(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__a22o_1 _15239_ (.A1(net274),
    .A2(net824),
    .B1(_02052_),
    .B2(_02058_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _15240_ (.A0(net258),
    .A1(_02059_),
    .S(_09351_),
    .X(_02060_));
 sky130_fd_sc_hd__a221o_1 _15241_ (.A1(\core.csr.cycleTimer.currentValue[36] ),
    .A2(net876),
    .B1(_02051_),
    .B2(net1003),
    .C1(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _15242_ (.A0(\core.csr.cycleTimer.currentValue[4] ),
    .A1(_02061_),
    .S(net880),
    .X(_02062_));
 sky130_fd_sc_hd__a21o_4 _15243_ (.A1(net1003),
    .A2(_02050_),
    .B1(_02062_),
    .X(_02063_));
 sky130_fd_sc_hd__a21oi_1 _15244_ (.A1(net1168),
    .A2(_02063_),
    .B1(_02049_),
    .Y(_02064_));
 sky130_fd_sc_hd__o21a_1 _15245_ (.A1(_09366_),
    .A2(_02049_),
    .B1(net1165),
    .X(_02065_));
 sky130_fd_sc_hd__or3_1 _15246_ (.A(net1174),
    .B(_02064_),
    .C(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__o221a_1 _15247_ (.A1(net1185),
    .A2(_07592_),
    .B1(_08421_),
    .B2(_04480_),
    .C1(net1284),
    .X(_02067_));
 sky130_fd_sc_hd__and3_1 _15248_ (.A(_02048_),
    .B(_02066_),
    .C(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__o21ai_2 _15249_ (.A1(_05848_),
    .A2(_02068_),
    .B1(_09150_),
    .Y(_02069_));
 sky130_fd_sc_hd__o211a_1 _15250_ (.A1(\core.pipe1_resultRegister[4] ),
    .A2(net656),
    .B1(_02069_),
    .C1(net1924),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _15251_ (.A0(_09387_),
    .A1(_09376_),
    .S(net942),
    .X(_02070_));
 sky130_fd_sc_hd__mux2_1 _15252_ (.A0(_09399_),
    .A1(_09384_),
    .S(net941),
    .X(_02071_));
 sky130_fd_sc_hd__or2_1 _15253_ (.A(net946),
    .B(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__mux2_1 _15254_ (.A0(_09395_),
    .A1(_09402_),
    .S(net942),
    .X(_02073_));
 sky130_fd_sc_hd__mux2_4 _15255_ (.A0(_09459_),
    .A1(_02073_),
    .S(net946),
    .X(_02074_));
 sky130_fd_sc_hd__o211a_1 _15256_ (.A1(net887),
    .A2(_02070_),
    .B1(_02072_),
    .C1(net947),
    .X(_02075_));
 sky130_fd_sc_hd__a21oi_2 _15257_ (.A1(net949),
    .A2(_02074_),
    .B1(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__or2_1 _15258_ (.A(net1324),
    .B(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__nor2_1 _15259_ (.A(_06691_),
    .B(net1011),
    .Y(_02078_));
 sky130_fd_sc_hd__a211o_1 _15260_ (.A1(_08435_),
    .A2(net1010),
    .B1(_02040_),
    .C1(_02078_),
    .X(_02079_));
 sky130_fd_sc_hd__o21a_1 _15261_ (.A1(net886),
    .A2(_09443_),
    .B1(_09225_),
    .X(_02080_));
 sky130_fd_sc_hd__o21ai_2 _15262_ (.A1(net949),
    .A2(_02080_),
    .B1(net826),
    .Y(_02081_));
 sky130_fd_sc_hd__a21oi_1 _15263_ (.A1(_05796_),
    .A2(net1322),
    .B1(net1319),
    .Y(_02082_));
 sky130_fd_sc_hd__nand2_1 _15264_ (.A(_05798_),
    .B(net1316),
    .Y(_02083_));
 sky130_fd_sc_hd__o221a_1 _15265_ (.A1(net1311),
    .A2(_02081_),
    .B1(_02082_),
    .B2(_05797_),
    .C1(_02079_),
    .X(_02084_));
 sky130_fd_sc_hd__a31o_1 _15266_ (.A1(_02077_),
    .A2(_02083_),
    .A3(_02084_),
    .B1(net1083),
    .X(_02085_));
 sky130_fd_sc_hd__nand2_1 _15267_ (.A(_05794_),
    .B(net1172),
    .Y(_02086_));
 sky130_fd_sc_hd__a22o_1 _15268_ (.A1(\core.csr.cycleTimer.currentValue[5] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[37] ),
    .X(_02087_));
 sky130_fd_sc_hd__a22o_1 _15269_ (.A1(\core.csr.instretTimer.currentValue[5] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[37] ),
    .X(_02088_));
 sky130_fd_sc_hd__or2_1 _15270_ (.A(net6),
    .B(_09362_),
    .X(_02089_));
 sky130_fd_sc_hd__mux2_1 _15271_ (.A0(\core.csr.traps.mip.csrReadData[5] ),
    .A1(\core.csr.traps.mtval.csrReadData[5] ),
    .S(net868),
    .X(_02090_));
 sky130_fd_sc_hd__a221o_1 _15272_ (.A1(\core.csr.traps.mcause.csrReadData[5] ),
    .A2(net872),
    .B1(net823),
    .B2(_02090_),
    .C1(net864),
    .X(_02091_));
 sky130_fd_sc_hd__o21a_1 _15273_ (.A1(\core.csr.trapReturnVector[5] ),
    .A2(net861),
    .B1(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__a221o_2 _15274_ (.A1(\core.csr.traps.mtvec.csrReadData[5] ),
    .A2(net906),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[5] ),
    .C1(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__mux2_1 _15275_ (.A0(\core.csr.traps.mie.currentValue[5] ),
    .A1(_02093_),
    .S(net909),
    .X(_02094_));
 sky130_fd_sc_hd__a211o_4 _15276_ (.A1(\core.csr.mconfigptr.currentValue[5] ),
    .A2(net855),
    .B1(_09361_),
    .C1(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__a22o_1 _15277_ (.A1(net275),
    .A2(net824),
    .B1(_02089_),
    .B2(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__mux2_1 _15278_ (.A0(net259),
    .A1(_02096_),
    .S(_09351_),
    .X(_02097_));
 sky130_fd_sc_hd__a221o_1 _15279_ (.A1(\core.csr.cycleTimer.currentValue[37] ),
    .A2(net876),
    .B1(_02088_),
    .B2(net1002),
    .C1(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__mux2_2 _15280_ (.A0(\core.csr.cycleTimer.currentValue[5] ),
    .A1(_02098_),
    .S(net880),
    .X(_02099_));
 sky130_fd_sc_hd__a21oi_4 _15281_ (.A1(net1003),
    .A2(_02087_),
    .B1(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__or2_1 _15282_ (.A(net1170),
    .B(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__nand2_1 _15283_ (.A(net1211),
    .B(_02086_),
    .Y(_02102_));
 sky130_fd_sc_hd__a221o_1 _15284_ (.A1(_02086_),
    .A2(_02101_),
    .B1(_02102_),
    .B2(net1165),
    .C1(net1174),
    .X(_02103_));
 sky130_fd_sc_hd__o221a_1 _15285_ (.A1(net1185),
    .A2(_07559_),
    .B1(_08435_),
    .B2(_04480_),
    .C1(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__a31o_1 _15286_ (.A1(net1284),
    .A2(_02085_),
    .A3(_02104_),
    .B1(_05764_),
    .X(_02105_));
 sky130_fd_sc_hd__nand2_1 _15287_ (.A(net656),
    .B(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__o211a_1 _15288_ (.A1(\core.pipe1_resultRegister[5] ),
    .A2(net656),
    .B1(_02106_),
    .C1(net1922),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _15289_ (.A0(_09442_),
    .A1(_09445_),
    .S(net941),
    .X(_02107_));
 sky130_fd_sc_hd__mux2_1 _15290_ (.A0(_09407_),
    .A1(_02107_),
    .S(net945),
    .X(_02108_));
 sky130_fd_sc_hd__mux2_1 _15291_ (.A0(_09444_),
    .A1(_09449_),
    .S(net941),
    .X(_02109_));
 sky130_fd_sc_hd__mux2_1 _15292_ (.A0(_09448_),
    .A1(_09451_),
    .S(net941),
    .X(_02110_));
 sky130_fd_sc_hd__mux2_1 _15293_ (.A0(_02109_),
    .A1(_02110_),
    .S(net945),
    .X(_02111_));
 sky130_fd_sc_hd__mux2_2 _15294_ (.A0(_02108_),
    .A1(_02111_),
    .S(net947),
    .X(_02112_));
 sky130_fd_sc_hd__o21a_1 _15295_ (.A1(net887),
    .A2(_09396_),
    .B1(_09225_),
    .X(_02113_));
 sky130_fd_sc_hd__o21ai_1 _15296_ (.A1(net949),
    .A2(_02113_),
    .B1(net826),
    .Y(_02114_));
 sky130_fd_sc_hd__inv_2 _15297_ (.A(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__a221o_1 _15298_ (.A1(_05711_),
    .A2(net1322),
    .B1(_07383_),
    .B2(_05713_),
    .C1(net1329),
    .X(_02116_));
 sky130_fd_sc_hd__a221o_1 _15299_ (.A1(_07374_),
    .A2(_02112_),
    .B1(_02115_),
    .B2(net1314),
    .C1(_02116_),
    .X(_02117_));
 sky130_fd_sc_hd__a21oi_1 _15300_ (.A1(_05712_),
    .A2(net1319),
    .B1(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__a21o_1 _15301_ (.A1(_08437_),
    .A2(net1010),
    .B1(net1326),
    .X(_02119_));
 sky130_fd_sc_hd__a21oi_1 _15302_ (.A1(_06688_),
    .A2(net1014),
    .B1(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__nand2_1 _15303_ (.A(_04479_),
    .B(_08437_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_1 _15304_ (.A(_05709_),
    .B(net1173),
    .Y(_02122_));
 sky130_fd_sc_hd__a22o_1 _15305_ (.A1(\core.csr.cycleTimer.currentValue[6] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[38] ),
    .X(_02123_));
 sky130_fd_sc_hd__a22o_1 _15306_ (.A1(\core.csr.instretTimer.currentValue[6] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[38] ),
    .X(_02124_));
 sky130_fd_sc_hd__a221o_1 _15307_ (.A1(\core.csr.cycleTimer.currentValue[38] ),
    .A2(net876),
    .B1(_02124_),
    .B2(net1002),
    .C1(net884),
    .X(_02125_));
 sky130_fd_sc_hd__and3_1 _15308_ (.A(\core.csr.traps.mcause.csrReadData[6] ),
    .B(_09283_),
    .C(_09293_),
    .X(_02126_));
 sky130_fd_sc_hd__mux2_1 _15309_ (.A0(\core.csr.traps.mip.csrReadData[6] ),
    .A1(\core.csr.traps.mtval.csrReadData[6] ),
    .S(net869),
    .X(_02127_));
 sky130_fd_sc_hd__a221o_1 _15310_ (.A1(\core.csr.trapReturnVector[6] ),
    .A2(net865),
    .B1(_02127_),
    .B2(_09302_),
    .C1(_02126_),
    .X(_02128_));
 sky130_fd_sc_hd__a211o_1 _15311_ (.A1(\core.csr.traps.mscratch.currentValue[6] ),
    .A2(_09305_),
    .B1(_09308_),
    .C1(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__a21oi_1 _15312_ (.A1(_04393_),
    .A2(_09308_),
    .B1(_09309_),
    .Y(_02130_));
 sky130_fd_sc_hd__a221o_1 _15313_ (.A1(\core.csr.traps.mie.currentValue[6] ),
    .A2(_09309_),
    .B1(_02129_),
    .B2(_02130_),
    .C1(_09310_),
    .X(_02131_));
 sky130_fd_sc_hd__or4_1 _15314_ (.A(\core.csr.traps.machinePreviousInterruptEnable ),
    .B(net1007),
    .C(_09272_),
    .D(_09306_),
    .X(_02132_));
 sky130_fd_sc_hd__o311a_1 _15315_ (.A1(net865),
    .A2(_09305_),
    .A3(_09312_),
    .B1(_02131_),
    .C1(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__a221o_1 _15316_ (.A1(\core.csr.mconfigptr.currentValue[6] ),
    .A2(_09315_),
    .B1(_09316_),
    .B2(_09301_),
    .C1(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__o221a_1 _15317_ (.A1(_09282_),
    .A2(_09317_),
    .B1(_09318_),
    .B2(net7),
    .C1(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__a311o_1 _15318_ (.A1(net276),
    .A2(_09283_),
    .A3(_09316_),
    .B1(_09319_),
    .C1(_02135_),
    .X(_02136_));
 sky130_fd_sc_hd__o311a_1 _15319_ (.A1(net260),
    .A2(_09278_),
    .A3(_09314_),
    .B1(_09320_),
    .C1(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__o221a_2 _15320_ (.A1(\core.csr.cycleTimer.currentValue[6] ),
    .A2(net880),
    .B1(_02125_),
    .B2(_02137_),
    .C1(_09281_),
    .X(_02138_));
 sky130_fd_sc_hd__a21oi_4 _15321_ (.A1(net1002),
    .A2(_02123_),
    .B1(_02138_),
    .Y(_02139_));
 sky130_fd_sc_hd__or3_2 _15322_ (.A(net873),
    .B(net913),
    .C(net906),
    .X(_02140_));
 sky130_fd_sc_hd__or3_2 _15323_ (.A(net865),
    .B(net823),
    .C(net902),
    .X(_02141_));
 sky130_fd_sc_hd__o21a_1 _15324_ (.A1(net1170),
    .A2(_02139_),
    .B1(_02122_),
    .X(_02142_));
 sky130_fd_sc_hd__a21oi_1 _15325_ (.A1(net1211),
    .A2(_02122_),
    .B1(net1209),
    .Y(_02143_));
 sky130_fd_sc_hd__or3_1 _15326_ (.A(net1083),
    .B(_02118_),
    .C(_02120_),
    .X(_02144_));
 sky130_fd_sc_hd__o311a_1 _15327_ (.A1(net1174),
    .A2(_02142_),
    .A3(_02143_),
    .B1(_02144_),
    .C1(_02121_),
    .X(_02145_));
 sky130_fd_sc_hd__o211a_1 _15328_ (.A1(net1184),
    .A2(_07551_),
    .B1(_02145_),
    .C1(net1284),
    .X(_02146_));
 sky130_fd_sc_hd__o21ai_2 _15329_ (.A1(_05679_),
    .A2(_02146_),
    .B1(net657),
    .Y(_02147_));
 sky130_fd_sc_hd__o211a_1 _15330_ (.A1(\core.pipe1_resultRegister[6] ),
    .A2(net656),
    .B1(_02147_),
    .C1(net1926),
    .X(_00449_));
 sky130_fd_sc_hd__nand2_1 _15331_ (.A(_05628_),
    .B(net1173),
    .Y(_02148_));
 sky130_fd_sc_hd__a22o_1 _15332_ (.A1(\core.csr.cycleTimer.currentValue[7] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[39] ),
    .X(_02149_));
 sky130_fd_sc_hd__a22o_1 _15333_ (.A1(\core.csr.instretTimer.currentValue[7] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[39] ),
    .X(_02150_));
 sky130_fd_sc_hd__or2_1 _15334_ (.A(net8),
    .B(_09362_),
    .X(_02151_));
 sky130_fd_sc_hd__mux2_1 _15335_ (.A0(\core.csr.traps.mip.csrReadData[7] ),
    .A1(\core.csr.traps.mtval.csrReadData[7] ),
    .S(net868),
    .X(_02152_));
 sky130_fd_sc_hd__a221o_1 _15336_ (.A1(\core.csr.traps.mcause.csrReadData[7] ),
    .A2(net872),
    .B1(net823),
    .B2(_02152_),
    .C1(net864),
    .X(_02153_));
 sky130_fd_sc_hd__o21a_1 _15337_ (.A1(\core.csr.trapReturnVector[7] ),
    .A2(net861),
    .B1(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__a221o_4 _15338_ (.A1(\core.csr.traps.mtvec.csrReadData[7] ),
    .A2(net905),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[7] ),
    .C1(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__mux2_1 _15339_ (.A0(\core.csr.traps.mie.currentValue[7] ),
    .A1(_02155_),
    .S(net909),
    .X(_02156_));
 sky130_fd_sc_hd__a211o_4 _15340_ (.A1(\core.csr.mconfigptr.currentValue[7] ),
    .A2(net855),
    .B1(_09361_),
    .C1(_02156_),
    .X(_02157_));
 sky130_fd_sc_hd__a22o_1 _15341_ (.A1(net277),
    .A2(net824),
    .B1(_02151_),
    .B2(_02157_),
    .X(_02158_));
 sky130_fd_sc_hd__mux2_1 _15342_ (.A0(net261),
    .A1(_02158_),
    .S(_09351_),
    .X(_02159_));
 sky130_fd_sc_hd__a221o_1 _15343_ (.A1(\core.csr.cycleTimer.currentValue[39] ),
    .A2(net876),
    .B1(_02150_),
    .B2(net1002),
    .C1(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__mux2_2 _15344_ (.A0(\core.csr.cycleTimer.currentValue[7] ),
    .A1(_02160_),
    .S(net880),
    .X(_02161_));
 sky130_fd_sc_hd__a21oi_4 _15345_ (.A1(net1002),
    .A2(_02149_),
    .B1(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hd__o21a_1 _15346_ (.A1(net1170),
    .A2(_02162_),
    .B1(_02148_),
    .X(_02163_));
 sky130_fd_sc_hd__a21oi_1 _15347_ (.A1(net1212),
    .A2(_02148_),
    .B1(net1209),
    .Y(_02164_));
 sky130_fd_sc_hd__o32a_1 _15348_ (.A1(net1174),
    .A2(_02163_),
    .A3(_02164_),
    .B1(_07542_),
    .B2(net1185),
    .X(_02165_));
 sky130_fd_sc_hd__o211a_1 _15349_ (.A1(_04480_),
    .A2(_08462_),
    .B1(_02165_),
    .C1(net1284),
    .X(_02166_));
 sky130_fd_sc_hd__o21ai_1 _15350_ (.A1(_08462_),
    .A2(net1015),
    .B1(net1329),
    .Y(_02167_));
 sky130_fd_sc_hd__a21oi_1 _15351_ (.A1(_06684_),
    .A2(net1014),
    .B1(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__mux2_1 _15352_ (.A0(_01976_),
    .A1(_01981_),
    .S(net939),
    .X(_02169_));
 sky130_fd_sc_hd__mux2_2 _15353_ (.A0(_09228_),
    .A1(_02169_),
    .S(net944),
    .X(_02170_));
 sky130_fd_sc_hd__inv_2 _15354_ (.A(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__mux2_1 _15355_ (.A0(_01980_),
    .A1(_01989_),
    .S(net939),
    .X(_02172_));
 sky130_fd_sc_hd__inv_2 _15356_ (.A(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__mux2_1 _15357_ (.A0(_01987_),
    .A1(_01992_),
    .S(net939),
    .X(_02174_));
 sky130_fd_sc_hd__mux2_1 _15358_ (.A0(_02172_),
    .A1(_02174_),
    .S(net944),
    .X(_02175_));
 sky130_fd_sc_hd__mux2_1 _15359_ (.A0(_02171_),
    .A1(_02175_),
    .S(net948),
    .X(_02176_));
 sky130_fd_sc_hd__o21a_1 _15360_ (.A1(_05630_),
    .A2(_07384_),
    .B1(_07381_),
    .X(_02177_));
 sky130_fd_sc_hd__o2bb2a_1 _15361_ (.A1_N(_05630_),
    .A2_N(net1322),
    .B1(_02177_),
    .B2(_05631_),
    .X(_02178_));
 sky130_fd_sc_hd__o21ai_1 _15362_ (.A1(net886),
    .A2(_09180_),
    .B1(_09225_),
    .Y(_02179_));
 sky130_fd_sc_hd__a21bo_1 _15363_ (.A1(net948),
    .A2(_02179_),
    .B1_N(net825),
    .X(_02180_));
 sky130_fd_sc_hd__o22a_2 _15364_ (.A1(net1324),
    .A2(_02176_),
    .B1(_02180_),
    .B2(net1309),
    .X(_02181_));
 sky130_fd_sc_hd__and3_1 _15365_ (.A(net1327),
    .B(_02178_),
    .C(_02181_),
    .X(_02182_));
 sky130_fd_sc_hd__o31a_1 _15366_ (.A1(net1083),
    .A2(_02168_),
    .A3(_02182_),
    .B1(_02166_),
    .X(_02183_));
 sky130_fd_sc_hd__o21ai_1 _15367_ (.A1(_05598_),
    .A2(_02183_),
    .B1(net655),
    .Y(_02184_));
 sky130_fd_sc_hd__o211a_1 _15368_ (.A1(\core.pipe1_resultRegister[7] ),
    .A2(net655),
    .B1(_02184_),
    .C1(net1921),
    .X(_00450_));
 sky130_fd_sc_hd__or2_1 _15369_ (.A(_08464_),
    .B(net1014),
    .X(_02185_));
 sky130_fd_sc_hd__o211a_1 _15370_ (.A1(_06687_),
    .A2(net1010),
    .B1(_02185_),
    .C1(net1329),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _15371_ (.A0(_09165_),
    .A1(_09196_),
    .S(net945),
    .X(_02187_));
 sky130_fd_sc_hd__inv_2 _15372_ (.A(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__mux2_1 _15373_ (.A0(_02179_),
    .A1(_02188_),
    .S(net948),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _15374_ (.A0(_07384_),
    .A1(_07379_),
    .S(_06312_),
    .X(_02190_));
 sky130_fd_sc_hd__a21oi_1 _15375_ (.A1(_07381_),
    .A2(_02190_),
    .B1(_06313_),
    .Y(_02191_));
 sky130_fd_sc_hd__o21ai_2 _15376_ (.A1(net950),
    .A2(_02170_),
    .B1(net825),
    .Y(_02192_));
 sky130_fd_sc_hd__o22a_1 _15377_ (.A1(net1324),
    .A2(_02189_),
    .B1(_02192_),
    .B2(net1309),
    .X(_02193_));
 sky130_fd_sc_hd__or3b_1 _15378_ (.A(_02186_),
    .B(_02191_),
    .C_N(_02193_),
    .X(_02194_));
 sky130_fd_sc_hd__o21ai_1 _15379_ (.A1(net1184),
    .A2(_07685_),
    .B1(net1282),
    .Y(_02195_));
 sky130_fd_sc_hd__nand2_1 _15380_ (.A(_06310_),
    .B(net1173),
    .Y(_02196_));
 sky130_fd_sc_hd__a22o_1 _15381_ (.A1(\core.csr.cycleTimer.currentValue[8] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[40] ),
    .X(_02197_));
 sky130_fd_sc_hd__a22o_1 _15382_ (.A1(\core.csr.instretTimer.currentValue[8] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[40] ),
    .X(_02198_));
 sky130_fd_sc_hd__or2_1 _15383_ (.A(\core.csr.traps.mie.currentValue[8] ),
    .B(net909),
    .X(_02199_));
 sky130_fd_sc_hd__o21ai_2 _15384_ (.A1(net922),
    .A2(_09306_),
    .B1(_09356_),
    .Y(_02200_));
 sky130_fd_sc_hd__mux2_1 _15385_ (.A0(\core.csr.traps.mip.csrReadData[8] ),
    .A1(\core.csr.traps.mtval.csrReadData[8] ),
    .S(net868),
    .X(_02201_));
 sky130_fd_sc_hd__a221o_1 _15386_ (.A1(\core.csr.traps.mcause.csrReadData[8] ),
    .A2(net872),
    .B1(net822),
    .B2(_02201_),
    .C1(net864),
    .X(_02202_));
 sky130_fd_sc_hd__o21a_2 _15387_ (.A1(\core.csr.trapReturnVector[8] ),
    .A2(net860),
    .B1(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _15388_ (.A0(_02203_),
    .A1(\core.csr.traps.mscratch.currentValue[8] ),
    .S(net902),
    .X(_02204_));
 sky130_fd_sc_hd__a211o_1 _15389_ (.A1(\core.csr.traps.mtvec.csrReadData[8] ),
    .A2(net906),
    .B1(_02204_),
    .C1(net913),
    .X(_02205_));
 sky130_fd_sc_hd__a31o_2 _15390_ (.A1(_09472_),
    .A2(_02199_),
    .A3(_02205_),
    .B1(_02200_),
    .X(_02206_));
 sky130_fd_sc_hd__o211a_1 _15391_ (.A1(\core.csr.mconfigptr.currentValue[8] ),
    .A2(_09356_),
    .B1(_09362_),
    .C1(_09352_),
    .X(_02207_));
 sky130_fd_sc_hd__a22o_1 _15392_ (.A1(net278),
    .A2(net824),
    .B1(_02206_),
    .B2(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__mux2_1 _15393_ (.A0(net262),
    .A1(_02208_),
    .S(_09351_),
    .X(_02209_));
 sky130_fd_sc_hd__a221o_1 _15394_ (.A1(\core.csr.cycleTimer.currentValue[40] ),
    .A2(net876),
    .B1(_02198_),
    .B2(net1003),
    .C1(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_2 _15395_ (.A0(\core.csr.cycleTimer.currentValue[8] ),
    .A1(_02210_),
    .S(net881),
    .X(_02211_));
 sky130_fd_sc_hd__a21oi_4 _15396_ (.A1(net1002),
    .A2(_02197_),
    .B1(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__o21ai_1 _15397_ (.A1(net1170),
    .A2(_02212_),
    .B1(_02196_),
    .Y(_02213_));
 sky130_fd_sc_hd__a21o_1 _15398_ (.A1(net1211),
    .A2(_02196_),
    .B1(net1209),
    .X(_02214_));
 sky130_fd_sc_hd__a32o_1 _15399_ (.A1(net1215),
    .A2(_02213_),
    .A3(_02214_),
    .B1(_08464_),
    .B2(net1274),
    .X(_02215_));
 sky130_fd_sc_hd__a211o_1 _15400_ (.A1(net1080),
    .A2(_02194_),
    .B1(_02195_),
    .C1(_02215_),
    .X(_02216_));
 sky130_fd_sc_hd__o21ai_2 _15401_ (.A1(net480),
    .A2(net1284),
    .B1(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_1 _15402_ (.A(net656),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__o211a_1 _15403_ (.A1(\core.pipe1_resultRegister[8] ),
    .A2(net656),
    .B1(_02218_),
    .C1(net1925),
    .X(_00451_));
 sky130_fd_sc_hd__o21a_1 _15404_ (.A1(_08489_),
    .A2(net1014),
    .B1(net1329),
    .X(_02219_));
 sky130_fd_sc_hd__o21ai_1 _15405_ (.A1(_06686_),
    .A2(net1010),
    .B1(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__o21ai_1 _15406_ (.A1(net949),
    .A2(_02108_),
    .B1(net826),
    .Y(_02221_));
 sky130_fd_sc_hd__mux2_1 _15407_ (.A0(_09388_),
    .A1(_09403_),
    .S(net887),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_2 _15408_ (.A0(_02113_),
    .A1(_02222_),
    .S(net947),
    .X(_02223_));
 sky130_fd_sc_hd__nand2_1 _15409_ (.A(_07374_),
    .B(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__mux2_1 _15410_ (.A0(_07384_),
    .A1(_07379_),
    .S(_05550_),
    .X(_02225_));
 sky130_fd_sc_hd__a22o_1 _15411_ (.A1(_05512_),
    .A2(_05548_),
    .B1(_07381_),
    .B2(_02225_),
    .X(_02226_));
 sky130_fd_sc_hd__o2111a_1 _15412_ (.A1(net1310),
    .A2(_02221_),
    .B1(_02224_),
    .C1(_02226_),
    .D1(net1079),
    .X(_02227_));
 sky130_fd_sc_hd__nand2_1 _15413_ (.A(_05547_),
    .B(net1172),
    .Y(_02228_));
 sky130_fd_sc_hd__a22o_1 _15414_ (.A1(\core.csr.cycleTimer.currentValue[9] ),
    .A2(net930),
    .B1(net926),
    .B2(\core.csr.cycleTimer.currentValue[41] ),
    .X(_02229_));
 sky130_fd_sc_hd__a22o_1 _15415_ (.A1(\core.csr.instretTimer.currentValue[9] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[41] ),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_1 _15416_ (.A0(\core.csr.traps.mip.csrReadData[9] ),
    .A1(\core.csr.traps.mtval.csrReadData[9] ),
    .S(net868),
    .X(_02231_));
 sky130_fd_sc_hd__a221o_1 _15417_ (.A1(\core.csr.traps.mcause.csrReadData[9] ),
    .A2(net872),
    .B1(net822),
    .B2(_02231_),
    .C1(net864),
    .X(_02232_));
 sky130_fd_sc_hd__o21a_1 _15418_ (.A1(\core.csr.trapReturnVector[9] ),
    .A2(net860),
    .B1(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__a221o_4 _15419_ (.A1(\core.csr.traps.mtvec.csrReadData[9] ),
    .A2(net905),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[9] ),
    .C1(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__mux2_1 _15420_ (.A0(\core.csr.traps.mie.currentValue[9] ),
    .A1(_02234_),
    .S(net909),
    .X(_02235_));
 sky130_fd_sc_hd__a221o_1 _15421_ (.A1(net279),
    .A2(net824),
    .B1(net855),
    .B2(\core.csr.mconfigptr.currentValue[9] ),
    .C1(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_1 _15422_ (.A0(net263),
    .A1(_02236_),
    .S(_09351_),
    .X(_02237_));
 sky130_fd_sc_hd__a221o_1 _15423_ (.A1(\core.csr.cycleTimer.currentValue[41] ),
    .A2(net876),
    .B1(_02230_),
    .B2(net1005),
    .C1(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_2 _15424_ (.A0(\core.csr.cycleTimer.currentValue[9] ),
    .A1(_02238_),
    .S(net880),
    .X(_02239_));
 sky130_fd_sc_hd__a21oi_4 _15425_ (.A1(net1004),
    .A2(_02229_),
    .B1(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__o21ai_1 _15426_ (.A1(net1169),
    .A2(_02240_),
    .B1(_02228_),
    .Y(_02241_));
 sky130_fd_sc_hd__a21o_1 _15427_ (.A1(net1211),
    .A2(_02228_),
    .B1(net1208),
    .X(_02242_));
 sky130_fd_sc_hd__a32o_1 _15428_ (.A1(net1215),
    .A2(_02241_),
    .A3(_02242_),
    .B1(_08489_),
    .B2(net1274),
    .X(_02243_));
 sky130_fd_sc_hd__a2bb2o_1 _15429_ (.A1_N(net1080),
    .A2_N(_02243_),
    .B1(_02227_),
    .B2(_02220_),
    .X(_02244_));
 sky130_fd_sc_hd__o211a_1 _15430_ (.A1(net1184),
    .A2(_07694_),
    .B1(_02244_),
    .C1(net1281),
    .X(_02245_));
 sky130_fd_sc_hd__o21ai_4 _15431_ (.A1(_05513_),
    .A2(_02245_),
    .B1(net657),
    .Y(_02246_));
 sky130_fd_sc_hd__o211a_1 _15432_ (.A1(\core.pipe1_resultRegister[9] ),
    .A2(net655),
    .B1(_02246_),
    .C1(net1921),
    .X(_00452_));
 sky130_fd_sc_hd__and3_1 _15433_ (.A(_06676_),
    .B(_06679_),
    .C(net1014),
    .X(_02247_));
 sky130_fd_sc_hd__a21o_1 _15434_ (.A1(_08503_),
    .A2(net1010),
    .B1(net1326),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _15435_ (.A0(_09446_),
    .A1(_09450_),
    .S(net945),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_4 _15436_ (.A0(_02080_),
    .A1(_02249_),
    .S(net947),
    .X(_02250_));
 sky130_fd_sc_hd__nand2_1 _15437_ (.A(_07374_),
    .B(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__o21ai_4 _15438_ (.A1(net949),
    .A2(_02074_),
    .B1(net825),
    .Y(_02252_));
 sky130_fd_sc_hd__a221oi_1 _15439_ (.A1(_05453_),
    .A2(net1322),
    .B1(_07383_),
    .B2(_05455_),
    .C1(net1329),
    .Y(_02253_));
 sky130_fd_sc_hd__o211a_1 _15440_ (.A1(net1311),
    .A2(_02252_),
    .B1(_02253_),
    .C1(_02251_),
    .X(_02254_));
 sky130_fd_sc_hd__a21bo_1 _15441_ (.A1(_05454_),
    .A2(net1319),
    .B1_N(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(net1274),
    .B(_08503_),
    .Y(_02256_));
 sky130_fd_sc_hd__nand2_1 _15443_ (.A(_05451_),
    .B(net1172),
    .Y(_02257_));
 sky130_fd_sc_hd__a22o_1 _15444_ (.A1(\core.csr.cycleTimer.currentValue[10] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[42] ),
    .X(_02258_));
 sky130_fd_sc_hd__a22o_1 _15445_ (.A1(\core.csr.instretTimer.currentValue[10] ),
    .A2(net918),
    .B1(net914),
    .B2(\core.csr.instretTimer.currentValue[42] ),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _15446_ (.A0(\core.csr.traps.mip.csrReadData[10] ),
    .A1(\core.csr.traps.mtval.csrReadData[10] ),
    .S(net868),
    .X(_02260_));
 sky130_fd_sc_hd__a221o_1 _15447_ (.A1(\core.csr.traps.mcause.csrReadData[10] ),
    .A2(net872),
    .B1(net822),
    .B2(_02260_),
    .C1(net864),
    .X(_02261_));
 sky130_fd_sc_hd__o21a_1 _15448_ (.A1(\core.csr.trapReturnVector[10] ),
    .A2(net860),
    .B1(_02261_),
    .X(_02262_));
 sky130_fd_sc_hd__a221o_4 _15449_ (.A1(\core.csr.traps.mtvec.csrReadData[10] ),
    .A2(net905),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[10] ),
    .C1(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _15450_ (.A0(\core.csr.traps.mie.currentValue[10] ),
    .A1(_02263_),
    .S(net909),
    .X(_02264_));
 sky130_fd_sc_hd__a221o_1 _15451_ (.A1(net265),
    .A2(net824),
    .B1(net855),
    .B2(\core.csr.mconfigptr.currentValue[10] ),
    .C1(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _15452_ (.A0(net254),
    .A1(_02265_),
    .S(_09351_),
    .X(_02266_));
 sky130_fd_sc_hd__a221o_1 _15453_ (.A1(\core.csr.cycleTimer.currentValue[42] ),
    .A2(net876),
    .B1(_02259_),
    .B2(net1003),
    .C1(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_2 _15454_ (.A0(\core.csr.cycleTimer.currentValue[10] ),
    .A1(_02267_),
    .S(net880),
    .X(_02268_));
 sky130_fd_sc_hd__a21oi_4 _15455_ (.A1(net1003),
    .A2(_02258_),
    .B1(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__o21a_1 _15456_ (.A1(net1169),
    .A2(_02269_),
    .B1(_02257_),
    .X(_02270_));
 sky130_fd_sc_hd__a21oi_1 _15457_ (.A1(net1211),
    .A2(_02257_),
    .B1(net1209),
    .Y(_02271_));
 sky130_fd_sc_hd__o211ai_1 _15458_ (.A1(_02247_),
    .A2(_02248_),
    .B1(_02255_),
    .C1(net1080),
    .Y(_02272_));
 sky130_fd_sc_hd__o311a_1 _15459_ (.A1(_09148_),
    .A2(_02270_),
    .A3(_02271_),
    .B1(_02272_),
    .C1(_02256_),
    .X(_02273_));
 sky130_fd_sc_hd__o211a_1 _15460_ (.A1(net1184),
    .A2(_07674_),
    .B1(_02273_),
    .C1(net1281),
    .X(_02274_));
 sky130_fd_sc_hd__o21ai_4 _15461_ (.A1(_05422_),
    .A2(_02274_),
    .B1(net657),
    .Y(_02275_));
 sky130_fd_sc_hd__o211a_1 _15462_ (.A1(\core.pipe1_resultRegister[10] ),
    .A2(net656),
    .B1(_02275_),
    .C1(net1920),
    .X(_00453_));
 sky130_fd_sc_hd__a21o_1 _15463_ (.A1(_06677_),
    .A2(_06678_),
    .B1(net1010),
    .X(_02276_));
 sky130_fd_sc_hd__o21a_1 _15464_ (.A1(_08367_),
    .A2(net1014),
    .B1(_02039_),
    .X(_02277_));
 sky130_fd_sc_hd__nand2_1 _15465_ (.A(_02276_),
    .B(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__mux2_1 _15466_ (.A0(_01984_),
    .A1(_01990_),
    .S(net944),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_4 _15467_ (.A0(_02043_),
    .A1(_02279_),
    .S(net948),
    .X(_02280_));
 sky130_fd_sc_hd__nand2_1 _15468_ (.A(_07374_),
    .B(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__o21ai_4 _15469_ (.A1(net950),
    .A2(_02032_),
    .B1(net825),
    .Y(_02282_));
 sky130_fd_sc_hd__o221a_1 _15470_ (.A1(_05369_),
    .A2(_07384_),
    .B1(net1309),
    .B2(_02282_),
    .C1(_02281_),
    .X(_02283_));
 sky130_fd_sc_hd__o221a_1 _15471_ (.A1(_05367_),
    .A2(_07379_),
    .B1(_07381_),
    .B2(_05365_),
    .C1(_02278_),
    .X(_02284_));
 sky130_fd_sc_hd__a21oi_1 _15472_ (.A1(_02283_),
    .A2(_02284_),
    .B1(net1083),
    .Y(_02285_));
 sky130_fd_sc_hd__nand2_1 _15473_ (.A(_05330_),
    .B(net1172),
    .Y(_02286_));
 sky130_fd_sc_hd__a21o_1 _15474_ (.A1(net1211),
    .A2(_02286_),
    .B1(_09364_),
    .X(_02287_));
 sky130_fd_sc_hd__a22o_1 _15475_ (.A1(\core.csr.cycleTimer.currentValue[11] ),
    .A2(net929),
    .B1(net925),
    .B2(\core.csr.cycleTimer.currentValue[43] ),
    .X(_02288_));
 sky130_fd_sc_hd__a22o_1 _15476_ (.A1(\core.csr.instretTimer.currentValue[11] ),
    .A2(net919),
    .B1(net915),
    .B2(\core.csr.instretTimer.currentValue[43] ),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _15477_ (.A0(\core.csr.traps.mip.csrReadData[11] ),
    .A1(\core.csr.traps.mtval.csrReadData[11] ),
    .S(net868),
    .X(_02290_));
 sky130_fd_sc_hd__a221o_1 _15478_ (.A1(\core.csr.traps.mcause.csrReadData[11] ),
    .A2(net872),
    .B1(net822),
    .B2(_02290_),
    .C1(net864),
    .X(_02291_));
 sky130_fd_sc_hd__o21a_1 _15479_ (.A1(\core.csr.trapReturnVector[11] ),
    .A2(net860),
    .B1(_02291_),
    .X(_02292_));
 sky130_fd_sc_hd__a221o_4 _15480_ (.A1(\core.csr.traps.mtvec.csrReadData[11] ),
    .A2(net905),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[11] ),
    .C1(_02292_),
    .X(_02293_));
 sky130_fd_sc_hd__mux2_1 _15481_ (.A0(\core.csr.traps.mie.currentValue[11] ),
    .A1(_02293_),
    .S(net909),
    .X(_02294_));
 sky130_fd_sc_hd__a22o_1 _15482_ (.A1(net266),
    .A2(net824),
    .B1(_02289_),
    .B2(net1005),
    .X(_02295_));
 sky130_fd_sc_hd__a211o_1 _15483_ (.A1(\core.csr.mconfigptr.currentValue[11] ),
    .A2(net856),
    .B1(_02294_),
    .C1(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__a211o_1 _15484_ (.A1(\core.csr.cycleTimer.currentValue[43] ),
    .A2(net877),
    .B1(_02296_),
    .C1(net884),
    .X(_02297_));
 sky130_fd_sc_hd__o21a_1 _15485_ (.A1(\core.csr.cycleTimer.currentValue[11] ),
    .A2(net880),
    .B1(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__a21oi_4 _15486_ (.A1(net1003),
    .A2(_02288_),
    .B1(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__o21ai_1 _15487_ (.A1(net1169),
    .A2(_02299_),
    .B1(_02286_),
    .Y(_02300_));
 sky130_fd_sc_hd__o21ai_1 _15488_ (.A1(net1184),
    .A2(_07666_),
    .B1(net1281),
    .Y(_02301_));
 sky130_fd_sc_hd__a31o_1 _15489_ (.A1(net1214),
    .A2(_02287_),
    .A3(_02300_),
    .B1(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__a211o_1 _15490_ (.A1(net1274),
    .A2(_08367_),
    .B1(_02285_),
    .C1(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__o21ai_4 _15491_ (.A1(net452),
    .A2(net1281),
    .B1(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__nand2_1 _15492_ (.A(net655),
    .B(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__o211a_1 _15493_ (.A1(\core.pipe1_resultRegister[11] ),
    .A2(net655),
    .B1(_02305_),
    .C1(net1920),
    .X(_00454_));
 sky130_fd_sc_hd__or2_1 _15494_ (.A(_08333_),
    .B(net1014),
    .X(_02306_));
 sky130_fd_sc_hd__o211a_1 _15495_ (.A1(_06681_),
    .A2(net1010),
    .B1(_02306_),
    .C1(net1329),
    .X(_02307_));
 sky130_fd_sc_hd__a21o_1 _15496_ (.A1(net944),
    .A2(_02033_),
    .B1(net950),
    .X(_02308_));
 sky130_fd_sc_hd__a21o_1 _15497_ (.A1(net886),
    .A2(_02031_),
    .B1(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__o21ai_2 _15498_ (.A1(net948),
    .A2(_02002_),
    .B1(_02309_),
    .Y(_02310_));
 sky130_fd_sc_hd__a21bo_1 _15499_ (.A1(net948),
    .A2(_01985_),
    .B1_N(net825),
    .X(_02311_));
 sky130_fd_sc_hd__mux2_1 _15500_ (.A0(net1322),
    .A1(net1316),
    .S(_05025_),
    .X(_02312_));
 sky130_fd_sc_hd__o21ai_1 _15501_ (.A1(net1319),
    .A2(_02312_),
    .B1(_05024_),
    .Y(_02313_));
 sky130_fd_sc_hd__o211a_1 _15502_ (.A1(net1309),
    .A2(_02311_),
    .B1(_02313_),
    .C1(net1079),
    .X(_02314_));
 sky130_fd_sc_hd__o21ai_1 _15503_ (.A1(net1324),
    .A2(_02310_),
    .B1(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__nand2_1 _15504_ (.A(_05022_),
    .B(net1172),
    .Y(_02316_));
 sky130_fd_sc_hd__a21o_1 _15505_ (.A1(net1211),
    .A2(_02316_),
    .B1(_09364_),
    .X(_02317_));
 sky130_fd_sc_hd__a22o_1 _15506_ (.A1(\core.csr.cycleTimer.currentValue[12] ),
    .A2(net930),
    .B1(net926),
    .B2(\core.csr.cycleTimer.currentValue[44] ),
    .X(_02318_));
 sky130_fd_sc_hd__a22o_1 _15507_ (.A1(\core.csr.instretTimer.currentValue[12] ),
    .A2(net919),
    .B1(net915),
    .B2(\core.csr.instretTimer.currentValue[44] ),
    .X(_02319_));
 sky130_fd_sc_hd__mux2_1 _15508_ (.A0(\core.csr.traps.mip.csrReadData[12] ),
    .A1(\core.csr.traps.mtval.csrReadData[12] ),
    .S(net868),
    .X(_02320_));
 sky130_fd_sc_hd__a221o_1 _15509_ (.A1(\core.csr.traps.mcause.csrReadData[12] ),
    .A2(net871),
    .B1(net822),
    .B2(_02320_),
    .C1(net863),
    .X(_02321_));
 sky130_fd_sc_hd__o21a_1 _15510_ (.A1(\core.csr.trapReturnVector[12] ),
    .A2(net860),
    .B1(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__a221o_4 _15511_ (.A1(\core.csr.traps.mtvec.csrReadData[12] ),
    .A2(net905),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[12] ),
    .C1(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _15512_ (.A0(\core.csr.traps.mie.currentValue[12] ),
    .A1(_02323_),
    .S(net909),
    .X(_02324_));
 sky130_fd_sc_hd__a22o_1 _15513_ (.A1(net267),
    .A2(_09353_),
    .B1(_02319_),
    .B2(net1005),
    .X(_02325_));
 sky130_fd_sc_hd__a211o_1 _15514_ (.A1(\core.csr.mconfigptr.currentValue[12] ),
    .A2(net856),
    .B1(_02324_),
    .C1(_02325_),
    .X(_02326_));
 sky130_fd_sc_hd__a211o_1 _15515_ (.A1(\core.csr.cycleTimer.currentValue[44] ),
    .A2(net877),
    .B1(_02326_),
    .C1(net884),
    .X(_02327_));
 sky130_fd_sc_hd__o21a_1 _15516_ (.A1(\core.csr.cycleTimer.currentValue[12] ),
    .A2(net881),
    .B1(_02327_),
    .X(_02328_));
 sky130_fd_sc_hd__a21oi_4 _15517_ (.A1(net1006),
    .A2(_02318_),
    .B1(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__o21ai_1 _15518_ (.A1(net1169),
    .A2(_02329_),
    .B1(_02316_),
    .Y(_02330_));
 sky130_fd_sc_hd__a32o_1 _15519_ (.A1(net1214),
    .A2(_02317_),
    .A3(_02330_),
    .B1(_08333_),
    .B2(net1274),
    .X(_02331_));
 sky130_fd_sc_hd__o22a_1 _15520_ (.A1(_02307_),
    .A2(_02315_),
    .B1(_02331_),
    .B2(net1080),
    .X(_02332_));
 sky130_fd_sc_hd__o21ai_1 _15521_ (.A1(net1184),
    .A2(_07641_),
    .B1(net1281),
    .Y(_02333_));
 sky130_fd_sc_hd__o22a_1 _15522_ (.A1(net1281),
    .A2(_08333_),
    .B1(_02332_),
    .B2(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__a21oi_1 _15523_ (.A1(net1881),
    .A2(net1258),
    .B1(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hd__nand2_1 _15524_ (.A(net657),
    .B(_02335_),
    .Y(_02336_));
 sky130_fd_sc_hd__o211a_1 _15525_ (.A1(\core.pipe1_resultRegister[12] ),
    .A2(net657),
    .B1(_02336_),
    .C1(net1908),
    .X(_00455_));
 sky130_fd_sc_hd__nor2_2 _15526_ (.A(net1229),
    .B(net1079),
    .Y(_02337_));
 sky130_fd_sc_hd__nand2_1 _15527_ (.A(net1227),
    .B(net1082),
    .Y(_02338_));
 sky130_fd_sc_hd__nand2_1 _15528_ (.A(_05107_),
    .B(net1172),
    .Y(_02339_));
 sky130_fd_sc_hd__a21o_1 _15529_ (.A1(net1212),
    .A2(_02339_),
    .B1(net1208),
    .X(_02340_));
 sky130_fd_sc_hd__a22o_1 _15530_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(net930),
    .B1(net926),
    .B2(\core.csr.cycleTimer.currentValue[45] ),
    .X(_02341_));
 sky130_fd_sc_hd__a22o_1 _15531_ (.A1(\core.csr.instretTimer.currentValue[13] ),
    .A2(net919),
    .B1(net915),
    .B2(\core.csr.instretTimer.currentValue[45] ),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _15532_ (.A0(\core.csr.traps.mip.csrReadData[13] ),
    .A1(\core.csr.traps.mtval.csrReadData[13] ),
    .S(net867),
    .X(_02343_));
 sky130_fd_sc_hd__a221o_1 _15533_ (.A1(\core.csr.traps.mcause.csrReadData[13] ),
    .A2(net871),
    .B1(net822),
    .B2(_02343_),
    .C1(net863),
    .X(_02344_));
 sky130_fd_sc_hd__o21a_1 _15534_ (.A1(\core.csr.trapReturnVector[13] ),
    .A2(net860),
    .B1(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__a221o_4 _15535_ (.A1(\core.csr.traps.mtvec.csrReadData[13] ),
    .A2(net904),
    .B1(net900),
    .B2(\core.csr.traps.mscratch.currentValue[13] ),
    .C1(_02345_),
    .X(_02346_));
 sky130_fd_sc_hd__mux2_1 _15536_ (.A0(\core.csr.traps.mie.currentValue[13] ),
    .A1(_02346_),
    .S(net909),
    .X(_02347_));
 sky130_fd_sc_hd__a22o_1 _15537_ (.A1(net268),
    .A2(_09353_),
    .B1(_02342_),
    .B2(net1005),
    .X(_02348_));
 sky130_fd_sc_hd__a211o_1 _15538_ (.A1(\core.csr.mconfigptr.currentValue[13] ),
    .A2(net855),
    .B1(_02347_),
    .C1(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__a211o_1 _15539_ (.A1(\core.csr.cycleTimer.currentValue[45] ),
    .A2(net877),
    .B1(_02349_),
    .C1(net884),
    .X(_02350_));
 sky130_fd_sc_hd__o21a_1 _15540_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(net881),
    .B1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__a21oi_4 _15541_ (.A1(net1005),
    .A2(_02341_),
    .B1(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__o21ai_1 _15542_ (.A1(net1169),
    .A2(_02352_),
    .B1(_02339_),
    .Y(_02353_));
 sky130_fd_sc_hd__a32o_1 _15543_ (.A1(net1214),
    .A2(_02340_),
    .A3(_02353_),
    .B1(_08332_),
    .B2(net1273),
    .X(_02354_));
 sky130_fd_sc_hd__or2_1 _15544_ (.A(net1030),
    .B(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__nand2_1 _15545_ (.A(net946),
    .B(_02071_),
    .Y(_02356_));
 sky130_fd_sc_hd__a21oi_1 _15546_ (.A1(net886),
    .A2(_02073_),
    .B1(net949),
    .Y(_02357_));
 sky130_fd_sc_hd__a22o_2 _15547_ (.A1(net949),
    .A2(_09460_),
    .B1(_02356_),
    .B2(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__o21ai_4 _15548_ (.A1(net949),
    .A2(_09447_),
    .B1(net826),
    .Y(_02359_));
 sky130_fd_sc_hd__mux2_1 _15549_ (.A0(net1320),
    .A1(net1316),
    .S(_05110_),
    .X(_02360_));
 sky130_fd_sc_hd__o21ai_1 _15550_ (.A1(net1319),
    .A2(_02360_),
    .B1(_05109_),
    .Y(_02361_));
 sky130_fd_sc_hd__and2_1 _15551_ (.A(_06703_),
    .B(net1013),
    .X(_02362_));
 sky130_fd_sc_hd__a211o_1 _15552_ (.A1(_08332_),
    .A2(net1011),
    .B1(net1207),
    .C1(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__o211a_1 _15553_ (.A1(net1323),
    .A2(_02358_),
    .B1(_02361_),
    .C1(net1327),
    .X(_02364_));
 sky130_fd_sc_hd__o21ai_1 _15554_ (.A1(net1308),
    .A2(_02359_),
    .B1(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__a21o_1 _15555_ (.A1(_02363_),
    .A2(_02365_),
    .B1(net1082),
    .X(_02366_));
 sky130_fd_sc_hd__a21o_1 _15556_ (.A1(_02355_),
    .A2(_02366_),
    .B1(net1295),
    .X(_02367_));
 sky130_fd_sc_hd__o21a_1 _15557_ (.A1(net1186),
    .A2(_07653_),
    .B1(_02367_),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _15558_ (.A0(_08332_),
    .A1(_02368_),
    .S(net1281),
    .X(_02369_));
 sky130_fd_sc_hd__a21bo_1 _15559_ (.A1(net1880),
    .A2(net1258),
    .B1_N(net657),
    .X(_02370_));
 sky130_fd_sc_hd__o221a_1 _15560_ (.A1(\core.pipe1_resultRegister[13] ),
    .A2(net657),
    .B1(_02369_),
    .B2(_02370_),
    .C1(net1908),
    .X(_00456_));
 sky130_fd_sc_hd__nand2_1 _15561_ (.A(_05275_),
    .B(net1171),
    .Y(_02371_));
 sky130_fd_sc_hd__a21o_1 _15562_ (.A1(net1212),
    .A2(_02371_),
    .B1(net1208),
    .X(_02372_));
 sky130_fd_sc_hd__a22o_1 _15563_ (.A1(\core.csr.cycleTimer.currentValue[14] ),
    .A2(net930),
    .B1(net926),
    .B2(\core.csr.cycleTimer.currentValue[46] ),
    .X(_02373_));
 sky130_fd_sc_hd__a22o_1 _15564_ (.A1(\core.csr.instretTimer.currentValue[14] ),
    .A2(net919),
    .B1(net915),
    .B2(\core.csr.instretTimer.currentValue[46] ),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _15565_ (.A0(\core.csr.traps.mip.csrReadData[14] ),
    .A1(\core.csr.traps.mtval.csrReadData[14] ),
    .S(net867),
    .X(_02375_));
 sky130_fd_sc_hd__a221o_1 _15566_ (.A1(\core.csr.traps.mcause.csrReadData[14] ),
    .A2(net871),
    .B1(net822),
    .B2(_02375_),
    .C1(net863),
    .X(_02376_));
 sky130_fd_sc_hd__o21a_1 _15567_ (.A1(\core.csr.trapReturnVector[14] ),
    .A2(net860),
    .B1(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__a221o_4 _15568_ (.A1(\core.csr.traps.mtvec.csrReadData[14] ),
    .A2(net905),
    .B1(net901),
    .B2(\core.csr.traps.mscratch.currentValue[14] ),
    .C1(_02377_),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _15569_ (.A0(\core.csr.traps.mie.currentValue[14] ),
    .A1(_02378_),
    .S(net909),
    .X(_02379_));
 sky130_fd_sc_hd__a22o_1 _15570_ (.A1(net269),
    .A2(_09353_),
    .B1(_02374_),
    .B2(net1005),
    .X(_02380_));
 sky130_fd_sc_hd__a211o_1 _15571_ (.A1(\core.csr.mconfigptr.currentValue[14] ),
    .A2(net855),
    .B1(_02379_),
    .C1(_02380_),
    .X(_02381_));
 sky130_fd_sc_hd__a211o_1 _15572_ (.A1(\core.csr.cycleTimer.currentValue[46] ),
    .A2(net877),
    .B1(_02381_),
    .C1(net884),
    .X(_02382_));
 sky130_fd_sc_hd__o21a_1 _15573_ (.A1(\core.csr.cycleTimer.currentValue[14] ),
    .A2(net881),
    .B1(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__a21oi_4 _15574_ (.A1(net1005),
    .A2(_02373_),
    .B1(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__o21ai_1 _15575_ (.A1(net1169),
    .A2(_02384_),
    .B1(_02371_),
    .Y(_02385_));
 sky130_fd_sc_hd__a32o_1 _15576_ (.A1(net1214),
    .A2(_02372_),
    .A3(_02385_),
    .B1(_08331_),
    .B2(net1273),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _15577_ (.A0(_02107_),
    .A1(_02109_),
    .S(net945),
    .X(_02387_));
 sky130_fd_sc_hd__mux2_4 _15578_ (.A0(_09408_),
    .A1(_02387_),
    .S(net947),
    .X(_02388_));
 sky130_fd_sc_hd__o21ai_4 _15579_ (.A1(net950),
    .A2(_09404_),
    .B1(net825),
    .Y(_02389_));
 sky130_fd_sc_hd__mux2_1 _15580_ (.A0(net1321),
    .A1(net1316),
    .S(_05278_),
    .X(_02390_));
 sky130_fd_sc_hd__o21a_1 _15581_ (.A1(net1317),
    .A2(_02390_),
    .B1(_05277_),
    .X(_02391_));
 sky130_fd_sc_hd__nand2_1 _15582_ (.A(_06709_),
    .B(net1013),
    .Y(_02392_));
 sky130_fd_sc_hd__a21oi_1 _15583_ (.A1(_08331_),
    .A2(net1009),
    .B1(net1207),
    .Y(_02393_));
 sky130_fd_sc_hd__a21oi_1 _15584_ (.A1(_07374_),
    .A2(_02388_),
    .B1(_02391_),
    .Y(_02394_));
 sky130_fd_sc_hd__o211a_1 _15585_ (.A1(net1308),
    .A2(_02389_),
    .B1(_02394_),
    .C1(net1327),
    .X(_02395_));
 sky130_fd_sc_hd__a21oi_2 _15586_ (.A1(_02392_),
    .A2(_02393_),
    .B1(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__o22a_1 _15587_ (.A1(net1030),
    .A2(_02386_),
    .B1(_02396_),
    .B2(net1082),
    .X(_02397_));
 sky130_fd_sc_hd__o2bb2a_1 _15588_ (.A1_N(net1183),
    .A2_N(_07630_),
    .B1(_02397_),
    .B2(net1295),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _15589_ (.A0(_08331_),
    .A1(_02398_),
    .S(net1281),
    .X(_02399_));
 sky130_fd_sc_hd__a21oi_1 _15590_ (.A1(net1878),
    .A2(net1258),
    .B1(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__nand2_1 _15591_ (.A(net657),
    .B(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__o211a_1 _15592_ (.A1(\core.pipe1_resultRegister[14] ),
    .A2(net657),
    .B1(_02401_),
    .C1(net1908),
    .X(_00457_));
 sky130_fd_sc_hd__nand2_1 _15593_ (.A(_05186_),
    .B(net1173),
    .Y(_02402_));
 sky130_fd_sc_hd__a21o_1 _15594_ (.A1(net1212),
    .A2(_02402_),
    .B1(net1208),
    .X(_02403_));
 sky130_fd_sc_hd__a22o_1 _15595_ (.A1(\core.csr.cycleTimer.currentValue[15] ),
    .A2(net930),
    .B1(net926),
    .B2(\core.csr.cycleTimer.currentValue[47] ),
    .X(_02404_));
 sky130_fd_sc_hd__a22o_1 _15596_ (.A1(\core.csr.instretTimer.currentValue[15] ),
    .A2(net919),
    .B1(net915),
    .B2(\core.csr.instretTimer.currentValue[47] ),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _15597_ (.A0(\core.csr.traps.mip.csrReadData[15] ),
    .A1(\core.csr.traps.mtval.csrReadData[15] ),
    .S(net867),
    .X(_02406_));
 sky130_fd_sc_hd__a221o_1 _15598_ (.A1(\core.csr.traps.mcause.csrReadData[15] ),
    .A2(net871),
    .B1(net821),
    .B2(_02406_),
    .C1(net863),
    .X(_02407_));
 sky130_fd_sc_hd__o21a_1 _15599_ (.A1(\core.csr.trapReturnVector[15] ),
    .A2(net859),
    .B1(_02407_),
    .X(_02408_));
 sky130_fd_sc_hd__a221o_4 _15600_ (.A1(\core.csr.traps.mtvec.csrReadData[15] ),
    .A2(net904),
    .B1(net900),
    .B2(\core.csr.traps.mscratch.currentValue[15] ),
    .C1(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _15601_ (.A0(\core.csr.traps.mie.currentValue[15] ),
    .A1(_02409_),
    .S(net910),
    .X(_02410_));
 sky130_fd_sc_hd__a22o_1 _15602_ (.A1(net270),
    .A2(_09353_),
    .B1(_02405_),
    .B2(net1005),
    .X(_02411_));
 sky130_fd_sc_hd__a211o_1 _15603_ (.A1(\core.csr.mconfigptr.currentValue[15] ),
    .A2(net855),
    .B1(_02410_),
    .C1(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__a211o_1 _15604_ (.A1(\core.csr.cycleTimer.currentValue[47] ),
    .A2(net877),
    .B1(_02412_),
    .C1(net884),
    .X(_02413_));
 sky130_fd_sc_hd__o21a_1 _15605_ (.A1(\core.csr.cycleTimer.currentValue[15] ),
    .A2(net881),
    .B1(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__a21oi_4 _15606_ (.A1(net1005),
    .A2(_02404_),
    .B1(_02414_),
    .Y(_02415_));
 sky130_fd_sc_hd__o21ai_1 _15607_ (.A1(net1169),
    .A2(_02415_),
    .B1(_02402_),
    .Y(_02416_));
 sky130_fd_sc_hd__a31o_1 _15608_ (.A1(net1214),
    .A2(_02403_),
    .A3(_02416_),
    .B1(net1030),
    .X(_02417_));
 sky130_fd_sc_hd__a21o_1 _15609_ (.A1(net1273),
    .A2(_08330_),
    .B1(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__o21ai_2 _15610_ (.A1(net950),
    .A2(_09181_),
    .B1(net825),
    .Y(_02419_));
 sky130_fd_sc_hd__mux2_1 _15611_ (.A0(_02169_),
    .A1(_02173_),
    .S(net944),
    .X(_02420_));
 sky130_fd_sc_hd__mux2_2 _15612_ (.A0(_09229_),
    .A1(_02420_),
    .S(net948),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _15613_ (.A0(net1321),
    .A1(net1316),
    .S(_05188_),
    .X(_02422_));
 sky130_fd_sc_hd__o22a_1 _15614_ (.A1(_05157_),
    .A2(_05187_),
    .B1(net1318),
    .B2(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__a2bb2o_1 _15615_ (.A1_N(net1308),
    .A2_N(_02419_),
    .B1(_02421_),
    .B2(_07374_),
    .X(_02424_));
 sky130_fd_sc_hd__o41a_1 _15616_ (.A1(net1328),
    .A2(net1082),
    .A3(_02423_),
    .A4(_02424_),
    .B1(_02418_),
    .X(_02425_));
 sky130_fd_sc_hd__a21o_1 _15617_ (.A1(_08330_),
    .A2(net1009),
    .B1(net1207),
    .X(_02426_));
 sky130_fd_sc_hd__a211o_1 _15618_ (.A1(_06670_),
    .A2(net1013),
    .B1(_02426_),
    .C1(net1081),
    .X(_02427_));
 sky130_fd_sc_hd__a21oi_1 _15619_ (.A1(_02425_),
    .A2(_02427_),
    .B1(net1294),
    .Y(_02428_));
 sky130_fd_sc_hd__a21oi_1 _15620_ (.A1(net1183),
    .A2(_07615_),
    .B1(_02428_),
    .Y(_02429_));
 sky130_fd_sc_hd__mux2_1 _15621_ (.A0(_08330_),
    .A1(_02429_),
    .S(net1280),
    .X(_02430_));
 sky130_fd_sc_hd__a21bo_1 _15622_ (.A1(\core.pipe0_currentInstruction[15] ),
    .A2(net1258),
    .B1_N(net654),
    .X(_02431_));
 sky130_fd_sc_hd__o221a_1 _15623_ (.A1(\core.pipe1_resultRegister[15] ),
    .A2(net654),
    .B1(_02430_),
    .B2(_02431_),
    .C1(net1908),
    .X(_00458_));
 sky130_fd_sc_hd__a21o_1 _15624_ (.A1(_08329_),
    .A2(net1009),
    .B1(net1207),
    .X(_02432_));
 sky130_fd_sc_hd__a21oi_1 _15625_ (.A1(_06705_),
    .A2(net1013),
    .B1(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__nand2_1 _15626_ (.A(net1313),
    .B(_02421_),
    .Y(_02434_));
 sky130_fd_sc_hd__a221oi_1 _15627_ (.A1(_06487_),
    .A2(net1321),
    .B1(net1316),
    .B2(_06488_),
    .C1(net1330),
    .Y(_02435_));
 sky130_fd_sc_hd__o221a_1 _15628_ (.A1(_06485_),
    .A2(_07381_),
    .B1(_02419_),
    .B2(net1323),
    .C1(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__a21oi_1 _15629_ (.A1(_02434_),
    .A2(_02436_),
    .B1(_02433_),
    .Y(_02437_));
 sky130_fd_sc_hd__or2_1 _15630_ (.A(_06482_),
    .B(_09234_),
    .X(_02438_));
 sky130_fd_sc_hd__a22o_1 _15631_ (.A1(\core.csr.cycleTimer.currentValue[16] ),
    .A2(net928),
    .B1(net924),
    .B2(\core.csr.cycleTimer.currentValue[48] ),
    .X(_02439_));
 sky130_fd_sc_hd__a22o_4 _15632_ (.A1(\core.csr.instretTimer.currentValue[16] ),
    .A2(net919),
    .B1(net915),
    .B2(\core.csr.instretTimer.currentValue[48] ),
    .X(_02440_));
 sky130_fd_sc_hd__o21ai_4 _15633_ (.A1(_02140_),
    .A2(_02141_),
    .B1(_09472_),
    .Y(_02441_));
 sky130_fd_sc_hd__o21ba_1 _15634_ (.A1(\core.csr.traps.mie.currentValue[16] ),
    .A2(net908),
    .B1_N(net819),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _15635_ (.A0(\core.csr.traps.mip.csrReadData[16] ),
    .A1(\core.csr.traps.mtval.csrReadData[16] ),
    .S(net867),
    .X(_02443_));
 sky130_fd_sc_hd__a221o_1 _15636_ (.A1(\core.csr.traps.mcause.csrReadData[16] ),
    .A2(net871),
    .B1(net821),
    .B2(_02443_),
    .C1(net863),
    .X(_02444_));
 sky130_fd_sc_hd__o21a_1 _15637_ (.A1(\core.csr.trapReturnVector[16] ),
    .A2(net859),
    .B1(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__a221o_1 _15638_ (.A1(\core.csr.traps.mtvec.csrReadData[16] ),
    .A2(net904),
    .B1(net900),
    .B2(\core.csr.traps.mscratch.currentValue[16] ),
    .C1(_02445_),
    .X(_02446_));
 sky130_fd_sc_hd__o21a_2 _15639_ (.A1(net912),
    .A2(_02446_),
    .B1(_02442_),
    .X(_02447_));
 sky130_fd_sc_hd__a221o_1 _15640_ (.A1(\core.csr.mconfigptr.currentValue[16] ),
    .A2(net856),
    .B1(_02440_),
    .B2(net1001),
    .C1(_02447_),
    .X(_02448_));
 sky130_fd_sc_hd__a211o_1 _15641_ (.A1(\core.csr.cycleTimer.currentValue[48] ),
    .A2(net875),
    .B1(_02448_),
    .C1(net883),
    .X(_02449_));
 sky130_fd_sc_hd__o21a_1 _15642_ (.A1(\core.csr.cycleTimer.currentValue[16] ),
    .A2(net879),
    .B1(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__a21oi_4 _15643_ (.A1(net1006),
    .A2(_02439_),
    .B1(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__o21ai_1 _15644_ (.A1(net1169),
    .A2(_02451_),
    .B1(_02438_),
    .Y(_02452_));
 sky130_fd_sc_hd__a21o_1 _15645_ (.A1(net1212),
    .A2(_02438_),
    .B1(net1208),
    .X(_02453_));
 sky130_fd_sc_hd__a32o_1 _15646_ (.A1(net1214),
    .A2(_02452_),
    .A3(_02453_),
    .B1(_08329_),
    .B2(net1272),
    .X(_02454_));
 sky130_fd_sc_hd__o22a_1 _15647_ (.A1(net1081),
    .A2(_02437_),
    .B1(_02454_),
    .B2(net1029),
    .X(_02455_));
 sky130_fd_sc_hd__o22a_1 _15648_ (.A1(net1186),
    .A2(_07767_),
    .B1(_02455_),
    .B2(net1294),
    .X(_02456_));
 sky130_fd_sc_hd__a22o_1 _15649_ (.A1(net1871),
    .A2(net1258),
    .B1(_08329_),
    .B2(net1286),
    .X(_02457_));
 sky130_fd_sc_hd__or3b_1 _15650_ (.A(_02456_),
    .B(_02457_),
    .C_N(net653),
    .X(_02458_));
 sky130_fd_sc_hd__o211a_1 _15651_ (.A1(\core.pipe1_resultRegister[16] ),
    .A2(net653),
    .B1(_02458_),
    .C1(net1907),
    .X(_00459_));
 sky130_fd_sc_hd__and3_1 _15652_ (.A(_06663_),
    .B(_06707_),
    .C(net1012),
    .X(_02459_));
 sky130_fd_sc_hd__a21o_1 _15653_ (.A1(_08328_),
    .A2(net1009),
    .B1(net1207),
    .X(_02460_));
 sky130_fd_sc_hd__nor2_1 _15654_ (.A(net1323),
    .B(_02389_),
    .Y(_02461_));
 sky130_fd_sc_hd__a221o_1 _15655_ (.A1(_06409_),
    .A2(net1321),
    .B1(net1316),
    .B2(_06410_),
    .C1(net1328),
    .X(_02462_));
 sky130_fd_sc_hd__a21o_1 _15656_ (.A1(net1313),
    .A2(_02388_),
    .B1(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__a211o_1 _15657_ (.A1(_06407_),
    .A2(net1318),
    .B1(_02461_),
    .C1(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__o21a_1 _15658_ (.A1(_02459_),
    .A2(_02460_),
    .B1(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__and2_1 _15659_ (.A(_06405_),
    .B(net1173),
    .X(_02466_));
 sky130_fd_sc_hd__a22o_1 _15660_ (.A1(\core.csr.cycleTimer.currentValue[17] ),
    .A2(net928),
    .B1(net924),
    .B2(\core.csr.cycleTimer.currentValue[49] ),
    .X(_02467_));
 sky130_fd_sc_hd__or2_1 _15661_ (.A(\core.csr.cycleTimer.currentValue[17] ),
    .B(net879),
    .X(_02468_));
 sky130_fd_sc_hd__a22o_4 _15662_ (.A1(\core.csr.instretTimer.currentValue[17] ),
    .A2(net920),
    .B1(net916),
    .B2(\core.csr.instretTimer.currentValue[49] ),
    .X(_02469_));
 sky130_fd_sc_hd__o21ba_1 _15663_ (.A1(\core.csr.traps.mie.currentValue[17] ),
    .A2(net908),
    .B1_N(net819),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _15664_ (.A0(\core.csr.traps.mip.csrReadData[17] ),
    .A1(\core.csr.traps.mtval.csrReadData[17] ),
    .S(net867),
    .X(_02471_));
 sky130_fd_sc_hd__a221o_1 _15665_ (.A1(\core.csr.traps.mcause.csrReadData[17] ),
    .A2(net871),
    .B1(net821),
    .B2(_02471_),
    .C1(net863),
    .X(_02472_));
 sky130_fd_sc_hd__o21a_1 _15666_ (.A1(\core.csr.trapReturnVector[17] ),
    .A2(net859),
    .B1(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__a221o_1 _15667_ (.A1(\core.csr.traps.mtvec.csrReadData[17] ),
    .A2(net904),
    .B1(net900),
    .B2(\core.csr.traps.mscratch.currentValue[17] ),
    .C1(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__o21a_2 _15668_ (.A1(net912),
    .A2(_02474_),
    .B1(_02470_),
    .X(_02475_));
 sky130_fd_sc_hd__a221o_1 _15669_ (.A1(\core.csr.mconfigptr.currentValue[17] ),
    .A2(net857),
    .B1(_02469_),
    .B2(_09244_),
    .C1(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__a211o_1 _15670_ (.A1(\core.csr.cycleTimer.currentValue[49] ),
    .A2(net875),
    .B1(_02476_),
    .C1(net883),
    .X(_02477_));
 sky130_fd_sc_hd__a22o_4 _15671_ (.A1(net1001),
    .A2(_02467_),
    .B1(_02468_),
    .B2(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__a21o_1 _15672_ (.A1(net1168),
    .A2(_02478_),
    .B1(_02466_),
    .X(_02479_));
 sky130_fd_sc_hd__o21ai_1 _15673_ (.A1(_09366_),
    .A2(_02466_),
    .B1(net1165),
    .Y(_02480_));
 sky130_fd_sc_hd__a32o_1 _15674_ (.A1(net1214),
    .A2(_02479_),
    .A3(_02480_),
    .B1(_08328_),
    .B2(net1273),
    .X(_02481_));
 sky130_fd_sc_hd__o22a_1 _15675_ (.A1(net1081),
    .A2(_02465_),
    .B1(_02481_),
    .B2(net1030),
    .X(_02482_));
 sky130_fd_sc_hd__o22a_1 _15676_ (.A1(net1186),
    .A2(_07758_),
    .B1(_02482_),
    .B2(net1294),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _15677_ (.A0(_08328_),
    .A1(_02483_),
    .S(net1280),
    .X(_02484_));
 sky130_fd_sc_hd__a21bo_1 _15678_ (.A1(net1867),
    .A2(_07493_),
    .B1_N(net653),
    .X(_02485_));
 sky130_fd_sc_hd__o221a_1 _15679_ (.A1(\core.pipe1_resultRegister[17] ),
    .A2(net653),
    .B1(_02484_),
    .B2(_02485_),
    .C1(net1906),
    .X(_00460_));
 sky130_fd_sc_hd__a21o_1 _15680_ (.A1(_08327_),
    .A2(net1009),
    .B1(net1207),
    .X(_02486_));
 sky130_fd_sc_hd__a21oi_1 _15681_ (.A1(_06665_),
    .A2(net1012),
    .B1(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__a221o_1 _15682_ (.A1(_06642_),
    .A2(net1320),
    .B1(net1317),
    .B2(_06640_),
    .C1(net1328),
    .X(_02488_));
 sky130_fd_sc_hd__a21oi_1 _15683_ (.A1(_06643_),
    .A2(net1372),
    .B1(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hd__o22a_2 _15684_ (.A1(net1308),
    .A2(_02358_),
    .B1(_02359_),
    .B2(net1323),
    .X(_02490_));
 sky130_fd_sc_hd__a21oi_2 _15685_ (.A1(_02489_),
    .A2(_02490_),
    .B1(_02487_),
    .Y(_02491_));
 sky130_fd_sc_hd__nor2_1 _15686_ (.A(_06637_),
    .B(_09234_),
    .Y(_02492_));
 sky130_fd_sc_hd__a22o_1 _15687_ (.A1(\core.csr.cycleTimer.currentValue[18] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[50] ),
    .X(_02493_));
 sky130_fd_sc_hd__or2_1 _15688_ (.A(\core.csr.cycleTimer.currentValue[18] ),
    .B(net878),
    .X(_02494_));
 sky130_fd_sc_hd__a22o_4 _15689_ (.A1(\core.csr.instretTimer.currentValue[18] ),
    .A2(net919),
    .B1(net915),
    .B2(\core.csr.instretTimer.currentValue[50] ),
    .X(_02495_));
 sky130_fd_sc_hd__o21ba_1 _15690_ (.A1(\core.csr.traps.mie.currentValue[18] ),
    .A2(net908),
    .B1_N(net818),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _15691_ (.A0(\core.csr.traps.mip.csrReadData[18] ),
    .A1(\core.csr.traps.mtval.csrReadData[18] ),
    .S(net867),
    .X(_02497_));
 sky130_fd_sc_hd__a221o_1 _15692_ (.A1(\core.csr.traps.mcause.csrReadData[18] ),
    .A2(net871),
    .B1(net821),
    .B2(_02497_),
    .C1(net863),
    .X(_02498_));
 sky130_fd_sc_hd__o21a_1 _15693_ (.A1(\core.csr.trapReturnVector[18] ),
    .A2(net859),
    .B1(_02498_),
    .X(_02499_));
 sky130_fd_sc_hd__a221o_1 _15694_ (.A1(\core.csr.traps.mtvec.csrReadData[18] ),
    .A2(net904),
    .B1(net900),
    .B2(\core.csr.traps.mscratch.currentValue[18] ),
    .C1(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__o21a_1 _15695_ (.A1(net912),
    .A2(_02500_),
    .B1(_02496_),
    .X(_02501_));
 sky130_fd_sc_hd__a221o_1 _15696_ (.A1(\core.csr.mconfigptr.currentValue[18] ),
    .A2(net854),
    .B1(_02495_),
    .B2(net1000),
    .C1(_02501_),
    .X(_02502_));
 sky130_fd_sc_hd__a211o_1 _15697_ (.A1(\core.csr.cycleTimer.currentValue[50] ),
    .A2(net874),
    .B1(_02502_),
    .C1(net882),
    .X(_02503_));
 sky130_fd_sc_hd__a22o_4 _15698_ (.A1(net999),
    .A2(_02493_),
    .B1(_02494_),
    .B2(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__a21o_1 _15699_ (.A1(net1168),
    .A2(_02504_),
    .B1(_02492_),
    .X(_02505_));
 sky130_fd_sc_hd__o21ai_1 _15700_ (.A1(net1210),
    .A2(_02492_),
    .B1(net1164),
    .Y(_02506_));
 sky130_fd_sc_hd__a32o_1 _15701_ (.A1(net1213),
    .A2(_02505_),
    .A3(_02506_),
    .B1(_08327_),
    .B2(net1272),
    .X(_02507_));
 sky130_fd_sc_hd__o22a_1 _15702_ (.A1(net1081),
    .A2(_02491_),
    .B1(_02507_),
    .B2(net1029),
    .X(_02508_));
 sky130_fd_sc_hd__o22a_1 _15703_ (.A1(net1186),
    .A2(_07747_),
    .B1(_02508_),
    .B2(net1294),
    .X(_02509_));
 sky130_fd_sc_hd__a22o_1 _15704_ (.A1(\core.pipe0_currentInstruction[18] ),
    .A2(net1257),
    .B1(_08327_),
    .B2(net1286),
    .X(_02510_));
 sky130_fd_sc_hd__or3b_1 _15705_ (.A(_02509_),
    .B(_02510_),
    .C_N(net653),
    .X(_02511_));
 sky130_fd_sc_hd__o211a_1 _15706_ (.A1(\core.pipe1_resultRegister[18] ),
    .A2(net653),
    .B1(_02511_),
    .C1(net1906),
    .X(_00461_));
 sky130_fd_sc_hd__a21o_1 _15707_ (.A1(_08326_),
    .A2(net1008),
    .B1(net1207),
    .X(_02512_));
 sky130_fd_sc_hd__a21oi_1 _15708_ (.A1(_06795_),
    .A2(net1012),
    .B1(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__a221o_1 _15709_ (.A1(_06563_),
    .A2(net1320),
    .B1(net1317),
    .B2(_06564_),
    .C1(net1328),
    .X(_02514_));
 sky130_fd_sc_hd__a21oi_1 _15710_ (.A1(_06565_),
    .A2(net1372),
    .B1(_02514_),
    .Y(_02515_));
 sky130_fd_sc_hd__o22a_2 _15711_ (.A1(net1309),
    .A2(_02310_),
    .B1(_02311_),
    .B2(net1324),
    .X(_02516_));
 sky130_fd_sc_hd__a21oi_2 _15712_ (.A1(_02515_),
    .A2(_02516_),
    .B1(_02513_),
    .Y(_02517_));
 sky130_fd_sc_hd__nor2_1 _15713_ (.A(_06560_),
    .B(_09234_),
    .Y(_02518_));
 sky130_fd_sc_hd__a22o_1 _15714_ (.A1(\core.csr.cycleTimer.currentValue[19] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[51] ),
    .X(_02519_));
 sky130_fd_sc_hd__or2_1 _15715_ (.A(\core.csr.cycleTimer.currentValue[19] ),
    .B(net878),
    .X(_02520_));
 sky130_fd_sc_hd__a22o_1 _15716_ (.A1(\core.csr.instretTimer.currentValue[19] ),
    .A2(net921),
    .B1(net917),
    .B2(\core.csr.instretTimer.currentValue[51] ),
    .X(_02521_));
 sky130_fd_sc_hd__o21ba_1 _15717_ (.A1(\core.csr.traps.mie.currentValue[19] ),
    .A2(net907),
    .B1_N(net819),
    .X(_02522_));
 sky130_fd_sc_hd__mux2_1 _15718_ (.A0(\core.csr.traps.mip.csrReadData[19] ),
    .A1(\core.csr.traps.mtval.csrReadData[19] ),
    .S(net867),
    .X(_02523_));
 sky130_fd_sc_hd__a221o_1 _15719_ (.A1(\core.csr.traps.mcause.csrReadData[19] ),
    .A2(net873),
    .B1(net821),
    .B2(_02523_),
    .C1(net865),
    .X(_02524_));
 sky130_fd_sc_hd__o21a_1 _15720_ (.A1(\core.csr.trapReturnVector[19] ),
    .A2(net859),
    .B1(_02524_),
    .X(_02525_));
 sky130_fd_sc_hd__a221o_1 _15721_ (.A1(\core.csr.traps.mtvec.csrReadData[19] ),
    .A2(net904),
    .B1(net900),
    .B2(\core.csr.traps.mscratch.currentValue[19] ),
    .C1(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__o21a_1 _15722_ (.A1(net911),
    .A2(_02526_),
    .B1(_02522_),
    .X(_02527_));
 sky130_fd_sc_hd__a221o_1 _15723_ (.A1(\core.csr.mconfigptr.currentValue[19] ),
    .A2(net854),
    .B1(_02521_),
    .B2(net1000),
    .C1(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__a211o_1 _15724_ (.A1(\core.csr.cycleTimer.currentValue[51] ),
    .A2(net874),
    .B1(_02528_),
    .C1(net882),
    .X(_02529_));
 sky130_fd_sc_hd__a22o_4 _15725_ (.A1(net1000),
    .A2(_02519_),
    .B1(_02520_),
    .B2(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__a21o_1 _15726_ (.A1(net1167),
    .A2(_02530_),
    .B1(_02518_),
    .X(_02531_));
 sky130_fd_sc_hd__o21ai_1 _15727_ (.A1(net1210),
    .A2(_02518_),
    .B1(net1164),
    .Y(_02532_));
 sky130_fd_sc_hd__a32o_1 _15728_ (.A1(net1213),
    .A2(_02531_),
    .A3(_02532_),
    .B1(_08326_),
    .B2(net1272),
    .X(_02533_));
 sky130_fd_sc_hd__o22a_1 _15729_ (.A1(net1081),
    .A2(_02517_),
    .B1(_02533_),
    .B2(net1029),
    .X(_02534_));
 sky130_fd_sc_hd__o22a_1 _15730_ (.A1(net1186),
    .A2(_07736_),
    .B1(_02534_),
    .B2(net1293),
    .X(_02535_));
 sky130_fd_sc_hd__a22o_1 _15731_ (.A1(net1855),
    .A2(net1257),
    .B1(_08326_),
    .B2(net1285),
    .X(_02536_));
 sky130_fd_sc_hd__or3b_1 _15732_ (.A(_02535_),
    .B(_02536_),
    .C_N(net651),
    .X(_02537_));
 sky130_fd_sc_hd__o211a_1 _15733_ (.A1(\core.pipe1_resultRegister[19] ),
    .A2(net654),
    .B1(_02537_),
    .C1(net1892),
    .X(_00462_));
 sky130_fd_sc_hd__and3_1 _15734_ (.A(_06657_),
    .B(_06708_),
    .C(net1012),
    .X(_02538_));
 sky130_fd_sc_hd__o21ai_1 _15735_ (.A1(_08324_),
    .A2(net1012),
    .B1(_02039_),
    .Y(_02539_));
 sky130_fd_sc_hd__nor2_1 _15736_ (.A(net1323),
    .B(_02282_),
    .Y(_02540_));
 sky130_fd_sc_hd__a221o_1 _15737_ (.A1(_06655_),
    .A2(net1320),
    .B1(net1317),
    .B2(_06653_),
    .C1(net1328),
    .X(_02541_));
 sky130_fd_sc_hd__a21o_1 _15738_ (.A1(_06656_),
    .A2(net1372),
    .B1(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__a211o_1 _15739_ (.A1(net1313),
    .A2(_02280_),
    .B1(_02540_),
    .C1(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__o21ai_1 _15740_ (.A1(_02538_),
    .A2(_02539_),
    .B1(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__and2_1 _15741_ (.A(_04926_),
    .B(net1171),
    .X(_02545_));
 sky130_fd_sc_hd__a22o_1 _15742_ (.A1(\core.csr.cycleTimer.currentValue[20] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[52] ),
    .X(_02546_));
 sky130_fd_sc_hd__or2_1 _15743_ (.A(\core.csr.cycleTimer.currentValue[20] ),
    .B(net878),
    .X(_02547_));
 sky130_fd_sc_hd__a22o_1 _15744_ (.A1(\core.csr.instretTimer.currentValue[20] ),
    .A2(net921),
    .B1(net917),
    .B2(\core.csr.instretTimer.currentValue[52] ),
    .X(_02548_));
 sky130_fd_sc_hd__o21ba_1 _15745_ (.A1(\core.csr.traps.mie.currentValue[20] ),
    .A2(net907),
    .B1_N(net818),
    .X(_02549_));
 sky130_fd_sc_hd__mux2_1 _15746_ (.A0(\core.csr.traps.mip.csrReadData[20] ),
    .A1(\core.csr.traps.mtval.csrReadData[20] ),
    .S(net866),
    .X(_02550_));
 sky130_fd_sc_hd__a221o_1 _15747_ (.A1(\core.csr.traps.mcause.csrReadData[20] ),
    .A2(net870),
    .B1(net820),
    .B2(_02550_),
    .C1(net862),
    .X(_02551_));
 sky130_fd_sc_hd__o21a_1 _15748_ (.A1(\core.csr.trapReturnVector[20] ),
    .A2(net858),
    .B1(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__a221o_1 _15749_ (.A1(\core.csr.traps.mtvec.csrReadData[20] ),
    .A2(net903),
    .B1(net899),
    .B2(\core.csr.traps.mscratch.currentValue[20] ),
    .C1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__o21a_2 _15750_ (.A1(net911),
    .A2(_02553_),
    .B1(_02549_),
    .X(_02554_));
 sky130_fd_sc_hd__a221o_1 _15751_ (.A1(\core.csr.mconfigptr.currentValue[20] ),
    .A2(net854),
    .B1(_02548_),
    .B2(net999),
    .C1(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__a211o_1 _15752_ (.A1(\core.csr.cycleTimer.currentValue[52] ),
    .A2(net874),
    .B1(_02555_),
    .C1(net882),
    .X(_02556_));
 sky130_fd_sc_hd__a22o_4 _15753_ (.A1(net1000),
    .A2(_02546_),
    .B1(_02547_),
    .B2(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__a21oi_1 _15754_ (.A1(net1167),
    .A2(_02557_),
    .B1(_02545_),
    .Y(_02558_));
 sky130_fd_sc_hd__o21a_1 _15755_ (.A1(net1210),
    .A2(_02545_),
    .B1(net1164),
    .X(_02559_));
 sky130_fd_sc_hd__o32a_1 _15756_ (.A1(net1174),
    .A2(_02558_),
    .A3(_02559_),
    .B1(_08324_),
    .B2(_04480_),
    .X(_02560_));
 sky130_fd_sc_hd__a22o_1 _15757_ (.A1(net1079),
    .A2(_02544_),
    .B1(_02560_),
    .B2(_02337_),
    .X(_02561_));
 sky130_fd_sc_hd__a22o_1 _15758_ (.A1(net1182),
    .A2(_07723_),
    .B1(_02561_),
    .B2(net1290),
    .X(_02562_));
 sky130_fd_sc_hd__o2bb2a_1 _15759_ (.A1_N(net1852),
    .A2_N(net1257),
    .B1(_08324_),
    .B2(net1277),
    .X(_02563_));
 sky130_fd_sc_hd__nand3_1 _15760_ (.A(net651),
    .B(_02562_),
    .C(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__o211a_1 _15761_ (.A1(\core.pipe1_resultRegister[20] ),
    .A2(net652),
    .B1(_02564_),
    .C1(net1891),
    .X(_00463_));
 sky130_fd_sc_hd__nand2_1 _15762_ (.A(_08323_),
    .B(net1008),
    .Y(_02565_));
 sky130_fd_sc_hd__nand3_1 _15763_ (.A(_06671_),
    .B(_06672_),
    .C(net1012),
    .Y(_02566_));
 sky130_fd_sc_hd__a221o_2 _15764_ (.A1(_04853_),
    .A2(net1320),
    .B1(net1317),
    .B2(_04851_),
    .C1(net1328),
    .X(_02567_));
 sky130_fd_sc_hd__a221o_1 _15765_ (.A1(_04854_),
    .A2(net1372),
    .B1(net1313),
    .B2(_02250_),
    .C1(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__o21ba_1 _15766_ (.A1(net1323),
    .A2(_02252_),
    .B1_N(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__a31o_1 _15767_ (.A1(_02039_),
    .A2(_02565_),
    .A3(_02566_),
    .B1(_02569_),
    .X(_02570_));
 sky130_fd_sc_hd__and2_1 _15768_ (.A(_04849_),
    .B(net1171),
    .X(_02571_));
 sky130_fd_sc_hd__a22o_1 _15769_ (.A1(\core.csr.cycleTimer.currentValue[21] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[53] ),
    .X(_02572_));
 sky130_fd_sc_hd__or2_1 _15770_ (.A(\core.csr.cycleTimer.currentValue[21] ),
    .B(net878),
    .X(_02573_));
 sky130_fd_sc_hd__a22o_1 _15771_ (.A1(\core.csr.instretTimer.currentValue[21] ),
    .A2(net921),
    .B1(net917),
    .B2(\core.csr.instretTimer.currentValue[53] ),
    .X(_02574_));
 sky130_fd_sc_hd__o21ba_1 _15772_ (.A1(\core.csr.traps.mie.currentValue[21] ),
    .A2(net907),
    .B1_N(net818),
    .X(_02575_));
 sky130_fd_sc_hd__mux2_1 _15773_ (.A0(\core.csr.traps.mip.csrReadData[21] ),
    .A1(\core.csr.traps.mtval.csrReadData[21] ),
    .S(net866),
    .X(_02576_));
 sky130_fd_sc_hd__a221o_1 _15774_ (.A1(\core.csr.traps.mcause.csrReadData[21] ),
    .A2(net870),
    .B1(net820),
    .B2(_02576_),
    .C1(net862),
    .X(_02577_));
 sky130_fd_sc_hd__o21a_1 _15775_ (.A1(\core.csr.trapReturnVector[21] ),
    .A2(net858),
    .B1(_02577_),
    .X(_02578_));
 sky130_fd_sc_hd__a221o_1 _15776_ (.A1(\core.csr.traps.mtvec.csrReadData[21] ),
    .A2(net903),
    .B1(net899),
    .B2(\core.csr.traps.mscratch.currentValue[21] ),
    .C1(_02578_),
    .X(_02579_));
 sky130_fd_sc_hd__o21a_2 _15777_ (.A1(net911),
    .A2(_02579_),
    .B1(_02575_),
    .X(_02580_));
 sky130_fd_sc_hd__a221o_1 _15778_ (.A1(\core.csr.mconfigptr.currentValue[21] ),
    .A2(net854),
    .B1(_02574_),
    .B2(net999),
    .C1(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__a211o_1 _15779_ (.A1(\core.csr.cycleTimer.currentValue[53] ),
    .A2(net874),
    .B1(_02581_),
    .C1(net882),
    .X(_02582_));
 sky130_fd_sc_hd__a22o_4 _15780_ (.A1(net1000),
    .A2(_02572_),
    .B1(_02573_),
    .B2(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__a21o_1 _15781_ (.A1(net1167),
    .A2(_02583_),
    .B1(_02571_),
    .X(_02584_));
 sky130_fd_sc_hd__o21ai_1 _15782_ (.A1(net1210),
    .A2(_02571_),
    .B1(net1164),
    .Y(_02585_));
 sky130_fd_sc_hd__a32o_1 _15783_ (.A1(net1213),
    .A2(_02584_),
    .A3(_02585_),
    .B1(_08323_),
    .B2(net1272),
    .X(_02586_));
 sky130_fd_sc_hd__o2bb2a_1 _15784_ (.A1_N(net1079),
    .A2_N(_02570_),
    .B1(_02586_),
    .B2(net1029),
    .X(_02587_));
 sky130_fd_sc_hd__o2bb2a_1 _15785_ (.A1_N(net1182),
    .A2_N(_07712_),
    .B1(_02587_),
    .B2(net1292),
    .X(_02588_));
 sky130_fd_sc_hd__a22o_1 _15786_ (.A1(\core.pipe0_currentInstruction[21] ),
    .A2(net1257),
    .B1(_08323_),
    .B2(net1285),
    .X(_02589_));
 sky130_fd_sc_hd__or3b_1 _15787_ (.A(_02588_),
    .B(_02589_),
    .C_N(net652),
    .X(_02590_));
 sky130_fd_sc_hd__o211a_1 _15788_ (.A1(\core.pipe1_resultRegister[21] ),
    .A2(net652),
    .B1(_02590_),
    .C1(net1888),
    .X(_00464_));
 sky130_fd_sc_hd__and3_1 _15789_ (.A(_06659_),
    .B(_06674_),
    .C(net1012),
    .X(_02591_));
 sky130_fd_sc_hd__o21ai_1 _15790_ (.A1(_08322_),
    .A2(net1012),
    .B1(_02039_),
    .Y(_02592_));
 sky130_fd_sc_hd__a221o_1 _15791_ (.A1(_04774_),
    .A2(net1320),
    .B1(net1317),
    .B2(_04773_),
    .C1(net1328),
    .X(_02593_));
 sky130_fd_sc_hd__a2bb2o_2 _15792_ (.A1_N(net1324),
    .A2_N(_02221_),
    .B1(_02223_),
    .B2(net1315),
    .X(_02594_));
 sky130_fd_sc_hd__a211o_1 _15793_ (.A1(_04777_),
    .A2(net1372),
    .B1(_02593_),
    .C1(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__o21ai_1 _15794_ (.A1(_02591_),
    .A2(_02592_),
    .B1(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__nand2_1 _15795_ (.A(_04770_),
    .B(net1171),
    .Y(_02597_));
 sky130_fd_sc_hd__a22o_1 _15796_ (.A1(\core.csr.cycleTimer.currentValue[22] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[54] ),
    .X(_02598_));
 sky130_fd_sc_hd__or2_1 _15797_ (.A(\core.csr.cycleTimer.currentValue[22] ),
    .B(net878),
    .X(_02599_));
 sky130_fd_sc_hd__a22o_1 _15798_ (.A1(\core.csr.instretTimer.currentValue[22] ),
    .A2(net921),
    .B1(net917),
    .B2(\core.csr.instretTimer.currentValue[54] ),
    .X(_02600_));
 sky130_fd_sc_hd__o21ba_1 _15799_ (.A1(\core.csr.traps.mie.currentValue[22] ),
    .A2(net907),
    .B1_N(net818),
    .X(_02601_));
 sky130_fd_sc_hd__mux2_1 _15800_ (.A0(\core.csr.traps.mip.csrReadData[22] ),
    .A1(\core.csr.traps.mtval.csrReadData[22] ),
    .S(net866),
    .X(_02602_));
 sky130_fd_sc_hd__a221o_1 _15801_ (.A1(\core.csr.traps.mcause.csrReadData[22] ),
    .A2(net870),
    .B1(net820),
    .B2(_02602_),
    .C1(net862),
    .X(_02603_));
 sky130_fd_sc_hd__o21a_1 _15802_ (.A1(\core.csr.trapReturnVector[22] ),
    .A2(net858),
    .B1(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__a221o_1 _15803_ (.A1(\core.csr.traps.mtvec.csrReadData[22] ),
    .A2(net903),
    .B1(net899),
    .B2(\core.csr.traps.mscratch.currentValue[22] ),
    .C1(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__o21a_2 _15804_ (.A1(net911),
    .A2(_02605_),
    .B1(_02601_),
    .X(_02606_));
 sky130_fd_sc_hd__a221o_2 _15805_ (.A1(\core.csr.mconfigptr.currentValue[22] ),
    .A2(net854),
    .B1(_02600_),
    .B2(net999),
    .C1(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__a211o_1 _15806_ (.A1(\core.csr.cycleTimer.currentValue[54] ),
    .A2(net874),
    .B1(_02607_),
    .C1(net882),
    .X(_02608_));
 sky130_fd_sc_hd__a22o_4 _15807_ (.A1(net999),
    .A2(_02598_),
    .B1(_02599_),
    .B2(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__a21boi_1 _15808_ (.A1(net1167),
    .A2(_02609_),
    .B1_N(_02597_),
    .Y(_02610_));
 sky130_fd_sc_hd__a21oi_1 _15809_ (.A1(net1212),
    .A2(_02597_),
    .B1(net1208),
    .Y(_02611_));
 sky130_fd_sc_hd__o32a_1 _15810_ (.A1(net1174),
    .A2(_02610_),
    .A3(_02611_),
    .B1(_08322_),
    .B2(_04480_),
    .X(_02612_));
 sky130_fd_sc_hd__a22o_1 _15811_ (.A1(net1079),
    .A2(_02596_),
    .B1(_02612_),
    .B2(_02337_),
    .X(_02613_));
 sky130_fd_sc_hd__a22o_1 _15812_ (.A1(net1182),
    .A2(_07716_),
    .B1(_02613_),
    .B2(net1290),
    .X(_02614_));
 sky130_fd_sc_hd__o2bb2a_1 _15813_ (.A1_N(\core.pipe0_currentInstruction[22] ),
    .A2_N(net1257),
    .B1(_08322_),
    .B2(net1276),
    .X(_02615_));
 sky130_fd_sc_hd__nand3_1 _15814_ (.A(net651),
    .B(_02614_),
    .C(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__o211a_1 _15815_ (.A1(\core.pipe1_resultRegister[22] ),
    .A2(net652),
    .B1(_02616_),
    .C1(net1888),
    .X(_00465_));
 sky130_fd_sc_hd__nand2_1 _15816_ (.A(_08321_),
    .B(net1008),
    .Y(_02617_));
 sky130_fd_sc_hd__o211a_1 _15817_ (.A1(_06661_),
    .A2(net1008),
    .B1(_02039_),
    .C1(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__a221o_1 _15818_ (.A1(_04696_),
    .A2(net1320),
    .B1(net1317),
    .B2(_04694_),
    .C1(net1328),
    .X(_02619_));
 sky130_fd_sc_hd__a21oi_1 _15819_ (.A1(_04697_),
    .A2(net1372),
    .B1(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__o22a_2 _15820_ (.A1(net1309),
    .A2(_02189_),
    .B1(_02192_),
    .B2(net1324),
    .X(_02621_));
 sky130_fd_sc_hd__a21oi_1 _15821_ (.A1(_02620_),
    .A2(_02621_),
    .B1(_02618_),
    .Y(_02622_));
 sky130_fd_sc_hd__and2_1 _15822_ (.A(_04692_),
    .B(net1171),
    .X(_02623_));
 sky130_fd_sc_hd__a22o_1 _15823_ (.A1(\core.csr.cycleTimer.currentValue[23] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[55] ),
    .X(_02624_));
 sky130_fd_sc_hd__or2_1 _15824_ (.A(\core.csr.cycleTimer.currentValue[23] ),
    .B(net878),
    .X(_02625_));
 sky130_fd_sc_hd__a22o_1 _15825_ (.A1(\core.csr.instretTimer.currentValue[23] ),
    .A2(net921),
    .B1(net917),
    .B2(\core.csr.instretTimer.currentValue[55] ),
    .X(_02626_));
 sky130_fd_sc_hd__o21ba_1 _15826_ (.A1(\core.csr.traps.mie.currentValue[23] ),
    .A2(net907),
    .B1_N(net818),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _15827_ (.A0(\core.csr.traps.mip.csrReadData[23] ),
    .A1(\core.csr.traps.mtval.csrReadData[23] ),
    .S(net866),
    .X(_02628_));
 sky130_fd_sc_hd__a221o_1 _15828_ (.A1(\core.csr.traps.mcause.csrReadData[23] ),
    .A2(net870),
    .B1(net820),
    .B2(_02628_),
    .C1(net862),
    .X(_02629_));
 sky130_fd_sc_hd__o21a_1 _15829_ (.A1(\core.csr.trapReturnVector[23] ),
    .A2(net858),
    .B1(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__a221o_1 _15830_ (.A1(\core.csr.traps.mtvec.csrReadData[23] ),
    .A2(net903),
    .B1(net899),
    .B2(\core.csr.traps.mscratch.currentValue[23] ),
    .C1(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__o21a_2 _15831_ (.A1(net911),
    .A2(_02631_),
    .B1(_02627_),
    .X(_02632_));
 sky130_fd_sc_hd__a221o_2 _15832_ (.A1(\core.csr.mconfigptr.currentValue[23] ),
    .A2(net854),
    .B1(_02626_),
    .B2(net999),
    .C1(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__a211o_1 _15833_ (.A1(\core.csr.cycleTimer.currentValue[55] ),
    .A2(net874),
    .B1(_02633_),
    .C1(net882),
    .X(_02634_));
 sky130_fd_sc_hd__a22o_4 _15834_ (.A1(net1000),
    .A2(_02624_),
    .B1(_02625_),
    .B2(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__a21o_1 _15835_ (.A1(net1167),
    .A2(_02635_),
    .B1(_02623_),
    .X(_02636_));
 sky130_fd_sc_hd__o21ai_1 _15836_ (.A1(net1210),
    .A2(_02623_),
    .B1(net1164),
    .Y(_02637_));
 sky130_fd_sc_hd__a32o_1 _15837_ (.A1(net1213),
    .A2(_02636_),
    .A3(_02637_),
    .B1(_08321_),
    .B2(net1272),
    .X(_02638_));
 sky130_fd_sc_hd__o22a_1 _15838_ (.A1(net1081),
    .A2(_02622_),
    .B1(_02638_),
    .B2(net1029),
    .X(_02639_));
 sky130_fd_sc_hd__o2bb2a_1 _15839_ (.A1_N(net1182),
    .A2_N(_07729_),
    .B1(_02639_),
    .B2(net1292),
    .X(_02640_));
 sky130_fd_sc_hd__a22o_1 _15840_ (.A1(net1831),
    .A2(net1257),
    .B1(_08321_),
    .B2(net1285),
    .X(_02641_));
 sky130_fd_sc_hd__or3b_2 _15841_ (.A(_02640_),
    .B(_02641_),
    .C_N(net651),
    .X(_02642_));
 sky130_fd_sc_hd__o211a_1 _15842_ (.A1(\core.pipe1_resultRegister[23] ),
    .A2(net652),
    .B1(_02642_),
    .C1(net1890),
    .X(_00466_));
 sky130_fd_sc_hd__nand2_1 _15843_ (.A(_08342_),
    .B(net1008),
    .Y(_02643_));
 sky130_fd_sc_hd__o211a_1 _15844_ (.A1(_06793_),
    .A2(net1008),
    .B1(_02039_),
    .C1(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__a21oi_1 _15845_ (.A1(_06790_),
    .A2(net1320),
    .B1(net1317),
    .Y(_02645_));
 sky130_fd_sc_hd__o22a_1 _15846_ (.A1(_06792_),
    .A2(_07384_),
    .B1(_02645_),
    .B2(_06789_),
    .X(_02646_));
 sky130_fd_sc_hd__o22a_2 _15847_ (.A1(net1309),
    .A2(_02176_),
    .B1(_02180_),
    .B2(net1324),
    .X(_02647_));
 sky130_fd_sc_hd__a31o_1 _15848_ (.A1(net1327),
    .A2(_02646_),
    .A3(_02647_),
    .B1(_02644_),
    .X(_02648_));
 sky130_fd_sc_hd__nand2_1 _15849_ (.A(_06787_),
    .B(net1171),
    .Y(_02649_));
 sky130_fd_sc_hd__a22o_1 _15850_ (.A1(\core.csr.cycleTimer.currentValue[24] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[56] ),
    .X(_02650_));
 sky130_fd_sc_hd__or2_1 _15851_ (.A(\core.csr.cycleTimer.currentValue[24] ),
    .B(net878),
    .X(_02651_));
 sky130_fd_sc_hd__a22o_1 _15852_ (.A1(\core.csr.instretTimer.currentValue[24] ),
    .A2(net921),
    .B1(net917),
    .B2(\core.csr.instretTimer.currentValue[56] ),
    .X(_02652_));
 sky130_fd_sc_hd__o21ba_1 _15853_ (.A1(\core.csr.traps.mie.currentValue[24] ),
    .A2(net907),
    .B1_N(net818),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _15854_ (.A0(\core.csr.traps.mip.csrReadData[24] ),
    .A1(\core.csr.traps.mtval.csrReadData[24] ),
    .S(net866),
    .X(_02654_));
 sky130_fd_sc_hd__a221o_1 _15855_ (.A1(\core.csr.traps.mcause.csrReadData[24] ),
    .A2(net870),
    .B1(net820),
    .B2(_02654_),
    .C1(net862),
    .X(_02655_));
 sky130_fd_sc_hd__o21a_1 _15856_ (.A1(\core.csr.trapReturnVector[24] ),
    .A2(net858),
    .B1(_02655_),
    .X(_02656_));
 sky130_fd_sc_hd__a221o_1 _15857_ (.A1(\core.csr.traps.mtvec.csrReadData[24] ),
    .A2(net903),
    .B1(net899),
    .B2(\core.csr.traps.mscratch.currentValue[24] ),
    .C1(_02656_),
    .X(_02657_));
 sky130_fd_sc_hd__o21a_2 _15858_ (.A1(net911),
    .A2(_02657_),
    .B1(_02653_),
    .X(_02658_));
 sky130_fd_sc_hd__a221o_2 _15859_ (.A1(\core.csr.mconfigptr.currentValue[24] ),
    .A2(net854),
    .B1(_02652_),
    .B2(net999),
    .C1(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__a211o_1 _15860_ (.A1(\core.csr.cycleTimer.currentValue[56] ),
    .A2(net874),
    .B1(_02659_),
    .C1(net882),
    .X(_02660_));
 sky130_fd_sc_hd__a22o_4 _15861_ (.A1(net1000),
    .A2(_02650_),
    .B1(_02651_),
    .B2(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__a21bo_1 _15862_ (.A1(net1167),
    .A2(_02661_),
    .B1_N(_02649_),
    .X(_02662_));
 sky130_fd_sc_hd__a21o_1 _15863_ (.A1(net1212),
    .A2(_02649_),
    .B1(net1208),
    .X(_02663_));
 sky130_fd_sc_hd__a32o_1 _15864_ (.A1(net1213),
    .A2(_02662_),
    .A3(_02663_),
    .B1(_08342_),
    .B2(net1272),
    .X(_02664_));
 sky130_fd_sc_hd__o2bb2a_1 _15865_ (.A1_N(net1079),
    .A2_N(_02648_),
    .B1(_02664_),
    .B2(net1029),
    .X(_02665_));
 sky130_fd_sc_hd__o2bb2a_1 _15866_ (.A1_N(net1182),
    .A2_N(_07785_),
    .B1(_02665_),
    .B2(net1292),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _15867_ (.A0(_08342_),
    .A1(_02666_),
    .S(net1276),
    .X(_02667_));
 sky130_fd_sc_hd__a21bo_1 _15868_ (.A1(net1825),
    .A2(net1257),
    .B1_N(net652),
    .X(_02668_));
 sky130_fd_sc_hd__o221a_1 _15869_ (.A1(\core.pipe1_resultRegister[24] ),
    .A2(net652),
    .B1(_02667_),
    .B2(_02668_),
    .C1(net1890),
    .X(_00467_));
 sky130_fd_sc_hd__and2_1 _15870_ (.A(_06865_),
    .B(net1171),
    .X(_02669_));
 sky130_fd_sc_hd__a22o_1 _15871_ (.A1(\core.csr.cycleTimer.currentValue[25] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[57] ),
    .X(_02670_));
 sky130_fd_sc_hd__or2_1 _15872_ (.A(\core.csr.cycleTimer.currentValue[25] ),
    .B(net878),
    .X(_02671_));
 sky130_fd_sc_hd__a22o_1 _15873_ (.A1(\core.csr.instretTimer.currentValue[25] ),
    .A2(net921),
    .B1(net917),
    .B2(\core.csr.instretTimer.currentValue[57] ),
    .X(_02672_));
 sky130_fd_sc_hd__o21ba_1 _15874_ (.A1(\core.csr.traps.mie.currentValue[25] ),
    .A2(net907),
    .B1_N(net818),
    .X(_02673_));
 sky130_fd_sc_hd__mux2_1 _15875_ (.A0(\core.csr.traps.mip.csrReadData[25] ),
    .A1(\core.csr.traps.mtval.csrReadData[25] ),
    .S(net866),
    .X(_02674_));
 sky130_fd_sc_hd__a221o_1 _15876_ (.A1(\core.csr.traps.mcause.csrReadData[25] ),
    .A2(net870),
    .B1(net821),
    .B2(_02674_),
    .C1(net862),
    .X(_02675_));
 sky130_fd_sc_hd__o21a_1 _15877_ (.A1(\core.csr.trapReturnVector[25] ),
    .A2(net859),
    .B1(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__a221o_1 _15878_ (.A1(\core.csr.traps.mtvec.csrReadData[25] ),
    .A2(net903),
    .B1(net899),
    .B2(\core.csr.traps.mscratch.currentValue[25] ),
    .C1(_02676_),
    .X(_02677_));
 sky130_fd_sc_hd__o21a_1 _15879_ (.A1(net911),
    .A2(_02677_),
    .B1(_02673_),
    .X(_02678_));
 sky130_fd_sc_hd__a221o_2 _15880_ (.A1(\core.csr.mconfigptr.currentValue[25] ),
    .A2(net854),
    .B1(_02672_),
    .B2(net999),
    .C1(_02678_),
    .X(_02679_));
 sky130_fd_sc_hd__a211o_1 _15881_ (.A1(\core.csr.cycleTimer.currentValue[57] ),
    .A2(net874),
    .B1(_02679_),
    .C1(net882),
    .X(_02680_));
 sky130_fd_sc_hd__a22o_4 _15882_ (.A1(net1000),
    .A2(_02670_),
    .B1(_02671_),
    .B2(_02680_),
    .X(_02681_));
 sky130_fd_sc_hd__a21o_1 _15883_ (.A1(net1167),
    .A2(_02681_),
    .B1(_02669_),
    .X(_02682_));
 sky130_fd_sc_hd__o21ai_1 _15884_ (.A1(net1210),
    .A2(_02669_),
    .B1(net1164),
    .Y(_02683_));
 sky130_fd_sc_hd__a31o_1 _15885_ (.A1(net1213),
    .A2(_02682_),
    .A3(_02683_),
    .B1(net1029),
    .X(_02684_));
 sky130_fd_sc_hd__a21o_1 _15886_ (.A1(net1272),
    .A2(_08341_),
    .B1(_02684_),
    .X(_02685_));
 sky130_fd_sc_hd__mux2_1 _15887_ (.A0(net1316),
    .A1(net1320),
    .S(_06868_),
    .X(_02686_));
 sky130_fd_sc_hd__o22a_4 _15888_ (.A1(_06836_),
    .A2(_06866_),
    .B1(net1317),
    .B2(_02686_),
    .X(_02687_));
 sky130_fd_sc_hd__a221o_4 _15889_ (.A1(net1314),
    .A2(_02112_),
    .B1(_02115_),
    .B2(_07374_),
    .C1(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__or3_1 _15890_ (.A(net1328),
    .B(net1081),
    .C(_02688_),
    .X(_02689_));
 sky130_fd_sc_hd__a21o_1 _15891_ (.A1(_08341_),
    .A2(net1008),
    .B1(net1207),
    .X(_02690_));
 sky130_fd_sc_hd__a211o_1 _15892_ (.A1(_06873_),
    .A2(net1013),
    .B1(_02690_),
    .C1(net1081),
    .X(_02691_));
 sky130_fd_sc_hd__and3_1 _15893_ (.A(_02685_),
    .B(_02689_),
    .C(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__o2bb2a_1 _15894_ (.A1_N(net1182),
    .A2_N(_07796_),
    .B1(_02692_),
    .B2(net1292),
    .X(_02693_));
 sky130_fd_sc_hd__mux2_1 _15895_ (.A0(_08341_),
    .A1(_02693_),
    .S(net1276),
    .X(_02694_));
 sky130_fd_sc_hd__a21bo_1 _15896_ (.A1(net1822),
    .A2(net1257),
    .B1_N(net652),
    .X(_02695_));
 sky130_fd_sc_hd__o221a_1 _15897_ (.A1(\core.pipe1_resultRegister[25] ),
    .A2(net652),
    .B1(_02694_),
    .B2(_02695_),
    .C1(net1892),
    .X(_00468_));
 sky130_fd_sc_hd__nand2_1 _15898_ (.A(_08340_),
    .B(net1008),
    .Y(_02696_));
 sky130_fd_sc_hd__o211a_1 _15899_ (.A1(_07120_),
    .A2(net1008),
    .B1(_02039_),
    .C1(_02696_),
    .X(_02697_));
 sky130_fd_sc_hd__o221a_1 _15900_ (.A1(_07023_),
    .A2(_07379_),
    .B1(_07381_),
    .B2(_07022_),
    .C1(net1327),
    .X(_02698_));
 sky130_fd_sc_hd__o22a_2 _15901_ (.A1(net1311),
    .A2(_02076_),
    .B1(_02081_),
    .B2(net1324),
    .X(_02699_));
 sky130_fd_sc_hd__o211a_1 _15902_ (.A1(_07024_),
    .A2(_07369_),
    .B1(_02698_),
    .C1(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__nor2_1 _15903_ (.A(_02697_),
    .B(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__nand2_1 _15904_ (.A(_07020_),
    .B(net1171),
    .Y(_02702_));
 sky130_fd_sc_hd__a22o_1 _15905_ (.A1(\core.csr.cycleTimer.currentValue[26] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[58] ),
    .X(_02703_));
 sky130_fd_sc_hd__or2_1 _15906_ (.A(\core.csr.cycleTimer.currentValue[26] ),
    .B(net879),
    .X(_02704_));
 sky130_fd_sc_hd__a22o_1 _15907_ (.A1(\core.csr.instretTimer.currentValue[26] ),
    .A2(net921),
    .B1(net917),
    .B2(\core.csr.instretTimer.currentValue[58] ),
    .X(_02705_));
 sky130_fd_sc_hd__o21ba_1 _15908_ (.A1(\core.csr.traps.mie.currentValue[26] ),
    .A2(net907),
    .B1_N(net818),
    .X(_02706_));
 sky130_fd_sc_hd__mux2_1 _15909_ (.A0(\core.csr.traps.mip.csrReadData[26] ),
    .A1(\core.csr.traps.mtval.csrReadData[26] ),
    .S(net866),
    .X(_02707_));
 sky130_fd_sc_hd__a221o_1 _15910_ (.A1(\core.csr.traps.mcause.csrReadData[26] ),
    .A2(net871),
    .B1(net820),
    .B2(_02707_),
    .C1(net863),
    .X(_02708_));
 sky130_fd_sc_hd__o21a_1 _15911_ (.A1(\core.csr.trapReturnVector[26] ),
    .A2(net858),
    .B1(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__a221o_1 _15912_ (.A1(\core.csr.traps.mtvec.csrReadData[26] ),
    .A2(net904),
    .B1(net900),
    .B2(\core.csr.traps.mscratch.currentValue[26] ),
    .C1(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__o21a_1 _15913_ (.A1(net912),
    .A2(_02710_),
    .B1(_02706_),
    .X(_02711_));
 sky130_fd_sc_hd__a221o_4 _15914_ (.A1(\core.csr.mconfigptr.currentValue[26] ),
    .A2(net854),
    .B1(_02705_),
    .B2(net999),
    .C1(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__a211o_1 _15915_ (.A1(\core.csr.cycleTimer.currentValue[58] ),
    .A2(net875),
    .B1(_02712_),
    .C1(net883),
    .X(_02713_));
 sky130_fd_sc_hd__a22o_4 _15916_ (.A1(net1001),
    .A2(_02703_),
    .B1(_02704_),
    .B2(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__a21bo_1 _15917_ (.A1(net1167),
    .A2(_02714_),
    .B1_N(_02702_),
    .X(_02715_));
 sky130_fd_sc_hd__a21o_1 _15918_ (.A1(net1212),
    .A2(_02702_),
    .B1(net1208),
    .X(_02716_));
 sky130_fd_sc_hd__a32o_1 _15919_ (.A1(net1213),
    .A2(_02715_),
    .A3(_02716_),
    .B1(_08340_),
    .B2(net1272),
    .X(_02717_));
 sky130_fd_sc_hd__o22a_1 _15920_ (.A1(net1081),
    .A2(_02701_),
    .B1(_02717_),
    .B2(net1029),
    .X(_02718_));
 sky130_fd_sc_hd__o2bb2a_1 _15921_ (.A1_N(net1182),
    .A2_N(_07801_),
    .B1(_02718_),
    .B2(net1292),
    .X(_02719_));
 sky130_fd_sc_hd__a22o_1 _15922_ (.A1(net1821),
    .A2(net1258),
    .B1(_08340_),
    .B2(net1286),
    .X(_02720_));
 sky130_fd_sc_hd__or3b_1 _15923_ (.A(_02719_),
    .B(_02720_),
    .C_N(net651),
    .X(_02721_));
 sky130_fd_sc_hd__o211a_1 _15924_ (.A1(\core.pipe1_resultRegister[26] ),
    .A2(net651),
    .B1(_02721_),
    .C1(net1892),
    .X(_00469_));
 sky130_fd_sc_hd__nand2_1 _15925_ (.A(_08339_),
    .B(net1008),
    .Y(_02722_));
 sky130_fd_sc_hd__o21ai_1 _15926_ (.A1(_07200_),
    .A2(_07201_),
    .B1(net1013),
    .Y(_02723_));
 sky130_fd_sc_hd__o221a_1 _15927_ (.A1(_06948_),
    .A2(_07379_),
    .B1(_07384_),
    .B2(_06950_),
    .C1(net1327),
    .X(_02724_));
 sky130_fd_sc_hd__o221a_1 _15928_ (.A1(net1308),
    .A2(_02037_),
    .B1(_02044_),
    .B2(net1323),
    .C1(_02724_),
    .X(_02725_));
 sky130_fd_sc_hd__o21a_1 _15929_ (.A1(_06947_),
    .A2(_07381_),
    .B1(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__a31o_1 _15930_ (.A1(_02039_),
    .A2(_02722_),
    .A3(_02723_),
    .B1(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__nor2_1 _15931_ (.A(_06943_),
    .B(_09234_),
    .Y(_02728_));
 sky130_fd_sc_hd__a22o_1 _15932_ (.A1(\core.csr.cycleTimer.currentValue[27] ),
    .A2(net928),
    .B1(net924),
    .B2(\core.csr.cycleTimer.currentValue[59] ),
    .X(_02729_));
 sky130_fd_sc_hd__or2_1 _15933_ (.A(\core.csr.cycleTimer.currentValue[27] ),
    .B(net879),
    .X(_02730_));
 sky130_fd_sc_hd__a22o_1 _15934_ (.A1(\core.csr.instretTimer.currentValue[27] ),
    .A2(net921),
    .B1(net917),
    .B2(\core.csr.instretTimer.currentValue[59] ),
    .X(_02731_));
 sky130_fd_sc_hd__o21ba_1 _15935_ (.A1(\core.csr.traps.mie.currentValue[27] ),
    .A2(net908),
    .B1_N(net819),
    .X(_02732_));
 sky130_fd_sc_hd__mux2_1 _15936_ (.A0(\core.csr.traps.mip.csrReadData[27] ),
    .A1(\core.csr.traps.mtval.csrReadData[27] ),
    .S(net867),
    .X(_02733_));
 sky130_fd_sc_hd__a221o_1 _15937_ (.A1(\core.csr.traps.mcause.csrReadData[27] ),
    .A2(net871),
    .B1(net820),
    .B2(_02733_),
    .C1(net863),
    .X(_02734_));
 sky130_fd_sc_hd__o21a_1 _15938_ (.A1(\core.csr.trapReturnVector[27] ),
    .A2(net858),
    .B1(_02734_),
    .X(_02735_));
 sky130_fd_sc_hd__a221o_1 _15939_ (.A1(\core.csr.traps.mtvec.csrReadData[27] ),
    .A2(net904),
    .B1(net899),
    .B2(\core.csr.traps.mscratch.currentValue[27] ),
    .C1(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__o21a_1 _15940_ (.A1(net911),
    .A2(_02736_),
    .B1(_02732_),
    .X(_02737_));
 sky130_fd_sc_hd__a221o_4 _15941_ (.A1(\core.csr.mconfigptr.currentValue[27] ),
    .A2(net854),
    .B1(_02731_),
    .B2(net999),
    .C1(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__a211o_1 _15942_ (.A1(\core.csr.cycleTimer.currentValue[59] ),
    .A2(net875),
    .B1(_02738_),
    .C1(net882),
    .X(_02739_));
 sky130_fd_sc_hd__a22o_4 _15943_ (.A1(net1001),
    .A2(_02729_),
    .B1(_02730_),
    .B2(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__a21o_1 _15944_ (.A1(net1167),
    .A2(_02740_),
    .B1(_02728_),
    .X(_02741_));
 sky130_fd_sc_hd__o21ai_1 _15945_ (.A1(net1210),
    .A2(_02728_),
    .B1(net1164),
    .Y(_02742_));
 sky130_fd_sc_hd__a32o_1 _15946_ (.A1(net1213),
    .A2(_02741_),
    .A3(_02742_),
    .B1(_08339_),
    .B2(net1272),
    .X(_02743_));
 sky130_fd_sc_hd__a2bb2o_1 _15947_ (.A1_N(net1029),
    .A2_N(_02743_),
    .B1(_02727_),
    .B2(net1079),
    .X(_02744_));
 sky130_fd_sc_hd__a22o_1 _15948_ (.A1(net1182),
    .A2(_07792_),
    .B1(_02744_),
    .B2(net1290),
    .X(_02745_));
 sky130_fd_sc_hd__nor2_1 _15949_ (.A(net1277),
    .B(_08339_),
    .Y(_02746_));
 sky130_fd_sc_hd__a21oi_1 _15950_ (.A1(net1277),
    .A2(_02745_),
    .B1(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__a21oi_1 _15951_ (.A1(net1820),
    .A2(net1257),
    .B1(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__nand2_1 _15952_ (.A(net653),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__o211a_1 _15953_ (.A1(\core.pipe1_resultRegister[27] ),
    .A2(net651),
    .B1(_02749_),
    .C1(net1891),
    .X(_00470_));
 sky130_fd_sc_hd__nand2_1 _15954_ (.A(net765),
    .B(net1009),
    .Y(_02750_));
 sky130_fd_sc_hd__nand2_1 _15955_ (.A(_07116_),
    .B(net1012),
    .Y(_02751_));
 sky130_fd_sc_hd__o221a_1 _15956_ (.A1(_07111_),
    .A2(_07379_),
    .B1(_07381_),
    .B2(_07110_),
    .C1(net1327),
    .X(_02752_));
 sky130_fd_sc_hd__o22a_2 _15957_ (.A1(net1310),
    .A2(_01998_),
    .B1(_02003_),
    .B2(net1325),
    .X(_02753_));
 sky130_fd_sc_hd__o211a_1 _15958_ (.A1(_07112_),
    .A2(_07369_),
    .B1(_02752_),
    .C1(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__a31o_1 _15959_ (.A1(_02039_),
    .A2(_02750_),
    .A3(_02751_),
    .B1(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__and2_1 _15960_ (.A(_07107_),
    .B(net1171),
    .X(_02756_));
 sky130_fd_sc_hd__a22o_1 _15961_ (.A1(\core.csr.cycleTimer.currentValue[28] ),
    .A2(net927),
    .B1(net923),
    .B2(\core.csr.cycleTimer.currentValue[60] ),
    .X(_02757_));
 sky130_fd_sc_hd__or2_1 _15962_ (.A(\core.csr.cycleTimer.currentValue[28] ),
    .B(net878),
    .X(_02758_));
 sky130_fd_sc_hd__a22o_4 _15963_ (.A1(\core.csr.instretTimer.currentValue[28] ),
    .A2(net920),
    .B1(net916),
    .B2(\core.csr.instretTimer.currentValue[60] ),
    .X(_02759_));
 sky130_fd_sc_hd__o21ba_1 _15964_ (.A1(\core.csr.traps.mie.currentValue[28] ),
    .A2(net907),
    .B1_N(net818),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _15965_ (.A0(\core.csr.traps.mip.csrReadData[28] ),
    .A1(\core.csr.traps.mtval.csrReadData[28] ),
    .S(net866),
    .X(_02761_));
 sky130_fd_sc_hd__a221o_1 _15966_ (.A1(\core.csr.traps.mcause.csrReadData[28] ),
    .A2(net870),
    .B1(net820),
    .B2(_02761_),
    .C1(net862),
    .X(_02762_));
 sky130_fd_sc_hd__o21a_1 _15967_ (.A1(\core.csr.trapReturnVector[28] ),
    .A2(net858),
    .B1(_02762_),
    .X(_02763_));
 sky130_fd_sc_hd__a221o_1 _15968_ (.A1(\core.csr.traps.mtvec.csrReadData[28] ),
    .A2(net903),
    .B1(net899),
    .B2(\core.csr.traps.mscratch.currentValue[28] ),
    .C1(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__o21a_4 _15969_ (.A1(net911),
    .A2(_02764_),
    .B1(_02760_),
    .X(_02765_));
 sky130_fd_sc_hd__a221o_1 _15970_ (.A1(\core.csr.mconfigptr.currentValue[28] ),
    .A2(net857),
    .B1(_02759_),
    .B2(net1001),
    .C1(_02765_),
    .X(_02766_));
 sky130_fd_sc_hd__a211o_1 _15971_ (.A1(\core.csr.cycleTimer.currentValue[60] ),
    .A2(net874),
    .B1(_02766_),
    .C1(net882),
    .X(_02767_));
 sky130_fd_sc_hd__a22o_4 _15972_ (.A1(net1001),
    .A2(_02757_),
    .B1(_02758_),
    .B2(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__a21o_1 _15973_ (.A1(net1167),
    .A2(_02768_),
    .B1(_02756_),
    .X(_02769_));
 sky130_fd_sc_hd__o21ai_1 _15974_ (.A1(net1210),
    .A2(_02756_),
    .B1(net1164),
    .Y(_02770_));
 sky130_fd_sc_hd__a32o_1 _15975_ (.A1(net1213),
    .A2(_02769_),
    .A3(_02770_),
    .B1(net765),
    .B2(net1272),
    .X(_02771_));
 sky130_fd_sc_hd__o2bb2a_1 _15976_ (.A1_N(net1079),
    .A2_N(_02755_),
    .B1(_02771_),
    .B2(net1029),
    .X(_02772_));
 sky130_fd_sc_hd__o22a_1 _15977_ (.A1(net1186),
    .A2(_07814_),
    .B1(_02772_),
    .B2(net1293),
    .X(_02773_));
 sky130_fd_sc_hd__a22o_1 _15978_ (.A1(net1819),
    .A2(net1257),
    .B1(net765),
    .B2(net1285),
    .X(_02774_));
 sky130_fd_sc_hd__or3b_2 _15979_ (.A(_02773_),
    .B(_02774_),
    .C_N(net651),
    .X(_02775_));
 sky130_fd_sc_hd__o211a_1 _15980_ (.A1(\core.pipe1_resultRegister[28] ),
    .A2(net652),
    .B1(_02775_),
    .C1(net1888),
    .X(_00471_));
 sky130_fd_sc_hd__or2_1 _15981_ (.A(_08093_),
    .B(net1012),
    .X(_02776_));
 sky130_fd_sc_hd__or3_1 _15982_ (.A(_07198_),
    .B(_07199_),
    .C(net1009),
    .X(_02777_));
 sky130_fd_sc_hd__nand2_1 _15983_ (.A(net1313),
    .B(_09456_),
    .Y(_02778_));
 sky130_fd_sc_hd__a221o_1 _15984_ (.A1(_07195_),
    .A2(net1320),
    .B1(net1317),
    .B2(_07194_),
    .C1(net1330),
    .X(_02779_));
 sky130_fd_sc_hd__a21oi_1 _15985_ (.A1(_07196_),
    .A2(net1372),
    .B1(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__o211a_1 _15986_ (.A1(net1323),
    .A2(_09461_),
    .B1(_02778_),
    .C1(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__a31o_1 _15987_ (.A1(_02039_),
    .A2(_02776_),
    .A3(_02777_),
    .B1(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__nand2_1 _15988_ (.A(_07190_),
    .B(net1171),
    .Y(_02783_));
 sky130_fd_sc_hd__a22o_1 _15989_ (.A1(\core.csr.cycleTimer.currentValue[29] ),
    .A2(net928),
    .B1(net924),
    .B2(\core.csr.cycleTimer.currentValue[61] ),
    .X(_02784_));
 sky130_fd_sc_hd__or2_1 _15990_ (.A(\core.csr.cycleTimer.currentValue[29] ),
    .B(net878),
    .X(_02785_));
 sky130_fd_sc_hd__a22o_2 _15991_ (.A1(\core.csr.instretTimer.currentValue[29] ),
    .A2(net920),
    .B1(net916),
    .B2(\core.csr.instretTimer.currentValue[61] ),
    .X(_02786_));
 sky130_fd_sc_hd__o21ba_1 _15992_ (.A1(\core.csr.traps.mie.currentValue[29] ),
    .A2(net908),
    .B1_N(net818),
    .X(_02787_));
 sky130_fd_sc_hd__mux2_1 _15993_ (.A0(\core.csr.traps.mip.csrReadData[29] ),
    .A1(\core.csr.traps.mtval.csrReadData[29] ),
    .S(net867),
    .X(_02788_));
 sky130_fd_sc_hd__a221o_1 _15994_ (.A1(\core.csr.traps.mcause.csrReadData[29] ),
    .A2(net870),
    .B1(net821),
    .B2(_02788_),
    .C1(net862),
    .X(_02789_));
 sky130_fd_sc_hd__o21a_1 _15995_ (.A1(\core.csr.trapReturnVector[29] ),
    .A2(net859),
    .B1(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__a221o_1 _15996_ (.A1(\core.csr.traps.mtvec.csrReadData[29] ),
    .A2(net903),
    .B1(net900),
    .B2(\core.csr.traps.mscratch.currentValue[29] ),
    .C1(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__o21a_4 _15997_ (.A1(net912),
    .A2(_02791_),
    .B1(_02787_),
    .X(_02792_));
 sky130_fd_sc_hd__a221o_1 _15998_ (.A1(\core.csr.mconfigptr.currentValue[29] ),
    .A2(net857),
    .B1(_02786_),
    .B2(net1001),
    .C1(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__a211o_1 _15999_ (.A1(\core.csr.cycleTimer.currentValue[61] ),
    .A2(net874),
    .B1(_02793_),
    .C1(net883),
    .X(_02794_));
 sky130_fd_sc_hd__a22o_4 _16000_ (.A1(net1001),
    .A2(_02784_),
    .B1(_02785_),
    .B2(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__a21boi_1 _16001_ (.A1(net1168),
    .A2(_02795_),
    .B1_N(_02783_),
    .Y(_02796_));
 sky130_fd_sc_hd__a21oi_1 _16002_ (.A1(net1212),
    .A2(_02783_),
    .B1(net1208),
    .Y(_02797_));
 sky130_fd_sc_hd__o32a_1 _16003_ (.A1(net1174),
    .A2(_02796_),
    .A3(_02797_),
    .B1(_08093_),
    .B2(_04480_),
    .X(_02798_));
 sky130_fd_sc_hd__a22o_1 _16004_ (.A1(net1079),
    .A2(_02782_),
    .B1(_02798_),
    .B2(_02337_),
    .X(_02799_));
 sky130_fd_sc_hd__a22o_1 _16005_ (.A1(net1183),
    .A2(_07536_),
    .B1(_02799_),
    .B2(net1290),
    .X(_02800_));
 sky130_fd_sc_hd__o2bb2a_1 _16006_ (.A1_N(\core.pipe0_currentInstruction[29] ),
    .A2_N(net1258),
    .B1(_08093_),
    .B2(net1280),
    .X(_02801_));
 sky130_fd_sc_hd__nand3_1 _16007_ (.A(net653),
    .B(_02800_),
    .C(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__o211a_1 _16008_ (.A1(\core.pipe1_resultRegister[29] ),
    .A2(net653),
    .B1(_02802_),
    .C1(net1906),
    .X(_00472_));
 sky130_fd_sc_hd__and2_1 _16009_ (.A(_07346_),
    .B(net1173),
    .X(_02803_));
 sky130_fd_sc_hd__a22o_1 _16010_ (.A1(\core.csr.cycleTimer.currentValue[30] ),
    .A2(_09273_),
    .B1(_09275_),
    .B2(\core.csr.cycleTimer.currentValue[62] ),
    .X(_02804_));
 sky130_fd_sc_hd__a22o_1 _16011_ (.A1(\core.csr.instretTimer.currentValue[30] ),
    .A2(net920),
    .B1(net916),
    .B2(\core.csr.instretTimer.currentValue[62] ),
    .X(_02805_));
 sky130_fd_sc_hd__a221o_1 _16012_ (.A1(\core.csr.cycleTimer.currentValue[62] ),
    .A2(_09288_),
    .B1(_02805_),
    .B2(net1006),
    .C1(net884),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _16013_ (.A0(\core.csr.traps.mip.csrReadData[30] ),
    .A1(\core.csr.traps.mtval.csrReadData[30] ),
    .S(net866),
    .X(_02807_));
 sky130_fd_sc_hd__a221o_1 _16014_ (.A1(\core.csr.traps.mcause.csrReadData[30] ),
    .A2(net870),
    .B1(net820),
    .B2(_02807_),
    .C1(net862),
    .X(_02808_));
 sky130_fd_sc_hd__o21a_1 _16015_ (.A1(\core.csr.trapReturnVector[30] ),
    .A2(net858),
    .B1(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _16016_ (.A0(_02809_),
    .A1(\core.csr.traps.mscratch.currentValue[30] ),
    .S(net899),
    .X(_02810_));
 sky130_fd_sc_hd__a211o_1 _16017_ (.A1(\core.csr.traps.mtvec.csrReadData[30] ),
    .A2(net903),
    .B1(_02810_),
    .C1(net911),
    .X(_02811_));
 sky130_fd_sc_hd__o21a_4 _16018_ (.A1(\core.csr.traps.mie.currentValue[30] ),
    .A2(net907),
    .B1(_02811_),
    .X(_02812_));
 sky130_fd_sc_hd__o22a_1 _16019_ (.A1(\core.csr.mconfigptr.currentValue[30] ),
    .A2(_09356_),
    .B1(_02200_),
    .B2(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__o22a_1 _16020_ (.A1(\core.csr.cycleTimer.currentValue[30] ),
    .A2(_09280_),
    .B1(_02806_),
    .B2(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__a21o_4 _16021_ (.A1(net1006),
    .A2(_02804_),
    .B1(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__a21o_1 _16022_ (.A1(net1168),
    .A2(_02815_),
    .B1(_02803_),
    .X(_02816_));
 sky130_fd_sc_hd__o21ai_1 _16023_ (.A1(net1210),
    .A2(_02803_),
    .B1(net1164),
    .Y(_02817_));
 sky130_fd_sc_hd__a32o_1 _16024_ (.A1(net1213),
    .A2(_02816_),
    .A3(_02817_),
    .B1(_08089_),
    .B2(net1273),
    .X(_02818_));
 sky130_fd_sc_hd__nor2_1 _16025_ (.A(net1323),
    .B(_09409_),
    .Y(_02819_));
 sky130_fd_sc_hd__mux2_1 _16026_ (.A0(net1316),
    .A1(net1321),
    .S(_07349_),
    .X(_02820_));
 sky130_fd_sc_hd__o22a_1 _16027_ (.A1(_07317_),
    .A2(_07347_),
    .B1(net1318),
    .B2(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__and3_1 _16028_ (.A(_07363_),
    .B(_07365_),
    .C(net1013),
    .X(_02822_));
 sky130_fd_sc_hd__a211o_1 _16029_ (.A1(_08089_),
    .A2(net1009),
    .B1(net1207),
    .C1(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__a2111o_1 _16030_ (.A1(net1313),
    .A2(_09405_),
    .B1(_02819_),
    .C1(_02821_),
    .D1(net1330),
    .X(_02824_));
 sky130_fd_sc_hd__a21o_1 _16031_ (.A1(_02823_),
    .A2(_02824_),
    .B1(net1081),
    .X(_02825_));
 sky130_fd_sc_hd__o21a_1 _16032_ (.A1(net1030),
    .A2(_02818_),
    .B1(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__o2bb2a_1 _16033_ (.A1_N(net1183),
    .A2_N(_07529_),
    .B1(_02826_),
    .B2(net1297),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _16034_ (.A0(_08089_),
    .A1(_02827_),
    .S(net1280),
    .X(_02828_));
 sky130_fd_sc_hd__a21bo_1 _16035_ (.A1(net1817),
    .A2(net1258),
    .B1_N(net653),
    .X(_02829_));
 sky130_fd_sc_hd__o221a_1 _16036_ (.A1(\core.pipe1_resultRegister[30] ),
    .A2(net654),
    .B1(_02828_),
    .B2(_02829_),
    .C1(net1907),
    .X(_00473_));
 sky130_fd_sc_hd__nor2_1 _16037_ (.A(_07273_),
    .B(_09234_),
    .Y(_02830_));
 sky130_fd_sc_hd__a22o_1 _16038_ (.A1(\core.csr.cycleTimer.currentValue[31] ),
    .A2(_09273_),
    .B1(_09275_),
    .B2(\core.csr.cycleTimer.currentValue[63] ),
    .X(_02831_));
 sky130_fd_sc_hd__or2_1 _16039_ (.A(\core.csr.cycleTimer.currentValue[31] ),
    .B(_09280_),
    .X(_02832_));
 sky130_fd_sc_hd__mux2_1 _16040_ (.A0(\core.csr.traps.mip.csrReadData[31] ),
    .A1(\core.csr.traps.mtval.csrReadData[31] ),
    .S(net866),
    .X(_02833_));
 sky130_fd_sc_hd__a22o_2 _16041_ (.A1(\core.csr.instretTimer.currentValue[31] ),
    .A2(net919),
    .B1(net915),
    .B2(\core.csr.instretTimer.currentValue[63] ),
    .X(_02834_));
 sky130_fd_sc_hd__o21ba_1 _16042_ (.A1(\core.csr.traps.mie.currentValue[31] ),
    .A2(net908),
    .B1_N(net819),
    .X(_02835_));
 sky130_fd_sc_hd__a221o_1 _16043_ (.A1(\core.csr.traps.mcause.csrReadData[31] ),
    .A2(net870),
    .B1(net820),
    .B2(_02833_),
    .C1(net862),
    .X(_02836_));
 sky130_fd_sc_hd__o21a_1 _16044_ (.A1(\core.csr.trapReturnVector[31] ),
    .A2(net858),
    .B1(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__a221o_1 _16045_ (.A1(\core.csr.traps.mtvec.csrReadData[31] ),
    .A2(net903),
    .B1(net899),
    .B2(\core.csr.traps.mscratch.currentValue[31] ),
    .C1(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__o21a_4 _16046_ (.A1(net912),
    .A2(_02838_),
    .B1(_02835_),
    .X(_02839_));
 sky130_fd_sc_hd__a221o_1 _16047_ (.A1(\core.csr.mconfigptr.currentValue[31] ),
    .A2(net856),
    .B1(_02834_),
    .B2(net1006),
    .C1(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__a211o_1 _16048_ (.A1(\core.csr.cycleTimer.currentValue[63] ),
    .A2(_09288_),
    .B1(_02840_),
    .C1(net884),
    .X(_02841_));
 sky130_fd_sc_hd__a22o_4 _16049_ (.A1(net1006),
    .A2(_02831_),
    .B1(_02832_),
    .B2(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__a21o_1 _16050_ (.A1(net1168),
    .A2(_02842_),
    .B1(_02830_),
    .X(_02843_));
 sky130_fd_sc_hd__o21ai_1 _16051_ (.A1(net1210),
    .A2(_02830_),
    .B1(net1164),
    .Y(_02844_));
 sky130_fd_sc_hd__a32o_1 _16052_ (.A1(net1214),
    .A2(_02843_),
    .A3(_02844_),
    .B1(_08091_),
    .B2(net1273),
    .X(_02845_));
 sky130_fd_sc_hd__nor2_1 _16053_ (.A(net1323),
    .B(_09230_),
    .Y(_02846_));
 sky130_fd_sc_hd__nor2_1 _16054_ (.A(_07360_),
    .B(_07369_),
    .Y(_02847_));
 sky130_fd_sc_hd__o21a_1 _16055_ (.A1(_07362_),
    .A2(_07364_),
    .B1(net1013),
    .X(_02848_));
 sky130_fd_sc_hd__a211o_1 _16056_ (.A1(_08091_),
    .A2(net1009),
    .B1(net1207),
    .C1(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__a21bo_1 _16057_ (.A1(_07275_),
    .A2(net1318),
    .B1_N(_07243_),
    .X(_02850_));
 sky130_fd_sc_hd__a21o_1 _16058_ (.A1(_07275_),
    .A2(net1321),
    .B1(_07380_),
    .X(_02851_));
 sky130_fd_sc_hd__a221o_1 _16059_ (.A1(net1313),
    .A2(_09216_),
    .B1(_02850_),
    .B2(_02851_),
    .C1(_02847_),
    .X(_02852_));
 sky130_fd_sc_hd__o31a_1 _16060_ (.A1(net1328),
    .A2(_02846_),
    .A3(_02852_),
    .B1(_02849_),
    .X(_02853_));
 sky130_fd_sc_hd__o22a_2 _16061_ (.A1(net1030),
    .A2(_02845_),
    .B1(_02853_),
    .B2(net1082),
    .X(_02854_));
 sky130_fd_sc_hd__o2bb2a_1 _16062_ (.A1_N(net1182),
    .A2_N(_07826_),
    .B1(_02854_),
    .B2(net1293),
    .X(_02855_));
 sky130_fd_sc_hd__a22o_1 _16063_ (.A1(net1815),
    .A2(net1258),
    .B1(_08091_),
    .B2(net1285),
    .X(_02856_));
 sky130_fd_sc_hd__or3b_1 _16064_ (.A(_02855_),
    .B(_02856_),
    .C_N(net651),
    .X(_02857_));
 sky130_fd_sc_hd__o211a_1 _16065_ (.A1(\core.pipe1_resultRegister[31] ),
    .A2(net651),
    .B1(_02857_),
    .C1(net1891),
    .X(_00474_));
 sky130_fd_sc_hd__nor2_2 _16066_ (.A(_04467_),
    .B(_08097_),
    .Y(_02858_));
 sky130_fd_sc_hd__and4bb_4 _16067_ (.A_N(net1765),
    .B_N(_08639_),
    .C(_08642_),
    .D(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__nand3_4 _16068_ (.A(_08642_),
    .B(net664),
    .C(_02858_),
    .Y(_02860_));
 sky130_fd_sc_hd__o21a_1 _16069_ (.A1(\core.pipe1_loadResult[0] ),
    .A2(net646),
    .B1(net1923),
    .X(_02861_));
 sky130_fd_sc_hd__o21a_1 _16070_ (.A1(_06152_),
    .A2(net586),
    .B1(_02861_),
    .X(_00475_));
 sky130_fd_sc_hd__nand2_1 _16071_ (.A(_06055_),
    .B(net646),
    .Y(_02862_));
 sky130_fd_sc_hd__o211a_1 _16072_ (.A1(\core.pipe1_loadResult[1] ),
    .A2(net646),
    .B1(_02862_),
    .C1(net1923),
    .X(_00476_));
 sky130_fd_sc_hd__nand2_1 _16073_ (.A(_05973_),
    .B(net646),
    .Y(_02863_));
 sky130_fd_sc_hd__o211a_1 _16074_ (.A1(\core.pipe1_loadResult[2] ),
    .A2(net646),
    .B1(_02863_),
    .C1(net1927),
    .X(_00477_));
 sky130_fd_sc_hd__nand2_1 _16075_ (.A(_05888_),
    .B(net647),
    .Y(_02864_));
 sky130_fd_sc_hd__o211a_1 _16076_ (.A1(\core.pipe1_loadResult[3] ),
    .A2(net647),
    .B1(_02864_),
    .C1(net1942),
    .X(_00478_));
 sky130_fd_sc_hd__nand2_1 _16077_ (.A(_05804_),
    .B(net650),
    .Y(_02865_));
 sky130_fd_sc_hd__o211a_1 _16078_ (.A1(\core.pipe1_loadResult[4] ),
    .A2(net650),
    .B1(_02865_),
    .C1(net1942),
    .X(_00479_));
 sky130_fd_sc_hd__nand2_1 _16079_ (.A(_05723_),
    .B(net647),
    .Y(_02866_));
 sky130_fd_sc_hd__o211a_1 _16080_ (.A1(\core.pipe1_loadResult[5] ),
    .A2(net647),
    .B1(_02866_),
    .C1(net1942),
    .X(_00480_));
 sky130_fd_sc_hd__nand2_1 _16081_ (.A(_05638_),
    .B(net646),
    .Y(_02867_));
 sky130_fd_sc_hd__o211a_1 _16082_ (.A1(\core.pipe1_loadResult[6] ),
    .A2(net646),
    .B1(_02867_),
    .C1(net1942),
    .X(_00481_));
 sky130_fd_sc_hd__o21a_1 _16083_ (.A1(\core.pipe1_loadResult[7] ),
    .A2(net647),
    .B1(net1940),
    .X(_02868_));
 sky130_fd_sc_hd__o21a_1 _16084_ (.A1(_04570_),
    .A2(net585),
    .B1(_02868_),
    .X(_00482_));
 sky130_fd_sc_hd__o21a_1 _16085_ (.A1(\core.pipe1_loadResult[8] ),
    .A2(_02859_),
    .B1(net1925),
    .X(_02869_));
 sky130_fd_sc_hd__o21a_1 _16086_ (.A1(_06145_),
    .A2(net586),
    .B1(_02869_),
    .X(_00483_));
 sky130_fd_sc_hd__o21a_1 _16087_ (.A1(\core.pipe1_loadResult[9] ),
    .A2(net646),
    .B1(net1923),
    .X(_02870_));
 sky130_fd_sc_hd__o21a_1 _16088_ (.A1(_05459_),
    .A2(net586),
    .B1(_02870_),
    .X(_00484_));
 sky130_fd_sc_hd__o21a_1 _16089_ (.A1(\core.pipe1_loadResult[10] ),
    .A2(net646),
    .B1(net1925),
    .X(_02871_));
 sky130_fd_sc_hd__o21a_1 _16090_ (.A1(_05372_),
    .A2(net586),
    .B1(_02871_),
    .X(_00485_));
 sky130_fd_sc_hd__o21a_1 _16091_ (.A1(\core.pipe1_loadResult[11] ),
    .A2(net647),
    .B1(net1940),
    .X(_02872_));
 sky130_fd_sc_hd__o21a_1 _16092_ (.A1(_05284_),
    .A2(net585),
    .B1(_02872_),
    .X(_00486_));
 sky130_fd_sc_hd__o21a_1 _16093_ (.A1(\core.pipe1_loadResult[12] ),
    .A2(net646),
    .B1(net1940),
    .X(_02873_));
 sky130_fd_sc_hd__o21a_1 _16094_ (.A1(_04939_),
    .A2(net586),
    .B1(_02873_),
    .X(_00487_));
 sky130_fd_sc_hd__o21a_1 _16095_ (.A1(\core.pipe1_loadResult[13] ),
    .A2(net647),
    .B1(net1940),
    .X(_02874_));
 sky130_fd_sc_hd__o21a_1 _16096_ (.A1(_05029_),
    .A2(net585),
    .B1(_02874_),
    .X(_00488_));
 sky130_fd_sc_hd__o21a_1 _16097_ (.A1(\core.pipe1_loadResult[14] ),
    .A2(net650),
    .B1(net1942),
    .X(_02875_));
 sky130_fd_sc_hd__o21a_1 _16098_ (.A1(_05195_),
    .A2(net585),
    .B1(_02875_),
    .X(_00489_));
 sky130_fd_sc_hd__a21bo_1 _16099_ (.A1(_04577_),
    .A2(_04578_),
    .B1_N(net647),
    .X(_02876_));
 sky130_fd_sc_hd__o211a_1 _16100_ (.A1(\core.pipe1_loadResult[15] ),
    .A2(net647),
    .B1(_02876_),
    .C1(net1940),
    .X(_00490_));
 sky130_fd_sc_hd__o21a_1 _16101_ (.A1(\core.pipe1_loadResult[16] ),
    .A2(net648),
    .B1(net1940),
    .X(_02877_));
 sky130_fd_sc_hd__o21a_1 _16102_ (.A1(_06155_),
    .A2(net585),
    .B1(_02877_),
    .X(_00491_));
 sky130_fd_sc_hd__o21a_1 _16103_ (.A1(\core.pipe1_loadResult[17] ),
    .A2(net648),
    .B1(net1940),
    .X(_02878_));
 sky130_fd_sc_hd__o21a_1 _16104_ (.A1(_05464_),
    .A2(net584),
    .B1(_02878_),
    .X(_00492_));
 sky130_fd_sc_hd__o21a_1 _16105_ (.A1(\core.pipe1_loadResult[18] ),
    .A2(_02859_),
    .B1(net1925),
    .X(_02879_));
 sky130_fd_sc_hd__o21a_1 _16106_ (.A1(_05376_),
    .A2(net586),
    .B1(_02879_),
    .X(_00493_));
 sky130_fd_sc_hd__o21a_1 _16107_ (.A1(\core.pipe1_loadResult[19] ),
    .A2(net647),
    .B1(net1940),
    .X(_02880_));
 sky130_fd_sc_hd__o21a_1 _16108_ (.A1(_05288_),
    .A2(net585),
    .B1(_02880_),
    .X(_00494_));
 sky130_fd_sc_hd__o21a_1 _16109_ (.A1(\core.pipe1_loadResult[20] ),
    .A2(net648),
    .B1(net1939),
    .X(_02881_));
 sky130_fd_sc_hd__o21a_1 _16110_ (.A1(_04857_),
    .A2(net584),
    .B1(_02881_),
    .X(_00495_));
 sky130_fd_sc_hd__o21a_1 _16111_ (.A1(\core.pipe1_loadResult[21] ),
    .A2(net648),
    .B1(net1941),
    .X(_02882_));
 sky130_fd_sc_hd__o21a_1 _16112_ (.A1(_04780_),
    .A2(net584),
    .B1(_02882_),
    .X(_00496_));
 sky130_fd_sc_hd__o21a_1 _16113_ (.A1(\core.pipe1_loadResult[22] ),
    .A2(net649),
    .B1(net1944),
    .X(_02883_));
 sky130_fd_sc_hd__o21a_1 _16114_ (.A1(_04700_),
    .A2(net585),
    .B1(_02883_),
    .X(_00497_));
 sky130_fd_sc_hd__a21bo_1 _16115_ (.A1(_04585_),
    .A2(_04586_),
    .B1_N(net649),
    .X(_02884_));
 sky130_fd_sc_hd__o211a_1 _16116_ (.A1(\core.pipe1_loadResult[23] ),
    .A2(net648),
    .B1(_02884_),
    .C1(net1944),
    .X(_00498_));
 sky130_fd_sc_hd__o21a_1 _16117_ (.A1(\core.pipe1_loadResult[24] ),
    .A2(net648),
    .B1(net1939),
    .X(_02885_));
 sky130_fd_sc_hd__o21a_1 _16118_ (.A1(_06141_),
    .A2(net584),
    .B1(_02885_),
    .X(_00499_));
 sky130_fd_sc_hd__o21a_1 _16119_ (.A1(\core.pipe1_loadResult[25] ),
    .A2(net648),
    .B1(net1939),
    .X(_02886_));
 sky130_fd_sc_hd__o21a_1 _16120_ (.A1(_05469_),
    .A2(net584),
    .B1(_02886_),
    .X(_00500_));
 sky130_fd_sc_hd__o21a_1 _16121_ (.A1(\core.pipe1_loadResult[26] ),
    .A2(net648),
    .B1(net1941),
    .X(_02887_));
 sky130_fd_sc_hd__o21a_1 _16122_ (.A1(_05381_),
    .A2(net584),
    .B1(_02887_),
    .X(_00501_));
 sky130_fd_sc_hd__o21a_1 _16123_ (.A1(\core.pipe1_loadResult[27] ),
    .A2(net648),
    .B1(net1939),
    .X(_02888_));
 sky130_fd_sc_hd__o21a_1 _16124_ (.A1(_05293_),
    .A2(net584),
    .B1(_02888_),
    .X(_00502_));
 sky130_fd_sc_hd__o21a_1 _16125_ (.A1(\core.pipe1_loadResult[28] ),
    .A2(net649),
    .B1(net1944),
    .X(_02889_));
 sky130_fd_sc_hd__o21a_1 _16126_ (.A1(_04952_),
    .A2(net585),
    .B1(_02889_),
    .X(_00503_));
 sky130_fd_sc_hd__o21a_1 _16127_ (.A1(\core.pipe1_loadResult[29] ),
    .A2(net648),
    .B1(net1939),
    .X(_02890_));
 sky130_fd_sc_hd__o21a_1 _16128_ (.A1(_05035_),
    .A2(net584),
    .B1(_02890_),
    .X(_00504_));
 sky130_fd_sc_hd__o21a_1 _16129_ (.A1(\core.pipe1_loadResult[30] ),
    .A2(net649),
    .B1(net1944),
    .X(_02891_));
 sky130_fd_sc_hd__o21a_1 _16130_ (.A1(_05201_),
    .A2(net584),
    .B1(_02891_),
    .X(_00505_));
 sky130_fd_sc_hd__o21a_1 _16131_ (.A1(\core.pipe1_loadResult[31] ),
    .A2(net649),
    .B1(net1941),
    .X(_02892_));
 sky130_fd_sc_hd__o21a_1 _16132_ (.A1(_04563_),
    .A2(net584),
    .B1(_02892_),
    .X(_00506_));
 sky130_fd_sc_hd__and3_2 _16133_ (.A(_08639_),
    .B(net697),
    .C(net1215),
    .X(_02893_));
 sky130_fd_sc_hd__nand2_1 _16134_ (.A(_09349_),
    .B(net643),
    .Y(_02894_));
 sky130_fd_sc_hd__o211a_1 _16135_ (.A1(\core.pipe1_csrData[0] ),
    .A2(net643),
    .B1(_02894_),
    .C1(net1924),
    .X(_00507_));
 sky130_fd_sc_hd__nand2_1 _16136_ (.A(_09432_),
    .B(net643),
    .Y(_02895_));
 sky130_fd_sc_hd__o211a_1 _16137_ (.A1(\core.pipe1_csrData[1] ),
    .A2(net643),
    .B1(_02895_),
    .C1(net1924),
    .X(_00508_));
 sky130_fd_sc_hd__nand2_1 _16138_ (.A(_01969_),
    .B(net641),
    .Y(_02896_));
 sky130_fd_sc_hd__o211a_1 _16139_ (.A1(\core.pipe1_csrData[2] ),
    .A2(net641),
    .B1(_02896_),
    .C1(net1924),
    .X(_00509_));
 sky130_fd_sc_hd__nand2_1 _16140_ (.A(_02024_),
    .B(net644),
    .Y(_02897_));
 sky130_fd_sc_hd__o211a_1 _16141_ (.A1(\core.pipe1_csrData[3] ),
    .A2(net644),
    .B1(_02897_),
    .C1(net1927),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _16142_ (.A0(\core.pipe1_csrData[4] ),
    .A1(_02063_),
    .S(net643),
    .X(_02898_));
 sky130_fd_sc_hd__and2_1 _16143_ (.A(net1925),
    .B(_02898_),
    .X(_00511_));
 sky130_fd_sc_hd__nand2_1 _16144_ (.A(_02100_),
    .B(net643),
    .Y(_02899_));
 sky130_fd_sc_hd__o211a_1 _16145_ (.A1(\core.pipe1_csrData[5] ),
    .A2(net644),
    .B1(_02899_),
    .C1(net1927),
    .X(_00512_));
 sky130_fd_sc_hd__nand2_1 _16146_ (.A(_02139_),
    .B(net644),
    .Y(_02900_));
 sky130_fd_sc_hd__o211a_1 _16147_ (.A1(\core.pipe1_csrData[6] ),
    .A2(net644),
    .B1(_02900_),
    .C1(net1927),
    .X(_00513_));
 sky130_fd_sc_hd__nand2_1 _16148_ (.A(_02162_),
    .B(net643),
    .Y(_02901_));
 sky130_fd_sc_hd__o211a_1 _16149_ (.A1(\core.pipe1_csrData[7] ),
    .A2(net643),
    .B1(_02901_),
    .C1(net1926),
    .X(_00514_));
 sky130_fd_sc_hd__nand2_1 _16150_ (.A(_02212_),
    .B(net642),
    .Y(_02902_));
 sky130_fd_sc_hd__o211a_1 _16151_ (.A1(\core.pipe1_csrData[8] ),
    .A2(net642),
    .B1(_02902_),
    .C1(net1924),
    .X(_00515_));
 sky130_fd_sc_hd__nand2_1 _16152_ (.A(_02240_),
    .B(net642),
    .Y(_02903_));
 sky130_fd_sc_hd__o211a_1 _16153_ (.A1(\core.pipe1_csrData[9] ),
    .A2(net642),
    .B1(_02903_),
    .C1(net1920),
    .X(_00516_));
 sky130_fd_sc_hd__nand2_1 _16154_ (.A(_02269_),
    .B(net642),
    .Y(_02904_));
 sky130_fd_sc_hd__o211a_1 _16155_ (.A1(\core.pipe1_csrData[10] ),
    .A2(net642),
    .B1(_02904_),
    .C1(net1920),
    .X(_00517_));
 sky130_fd_sc_hd__nand2_1 _16156_ (.A(_02299_),
    .B(net641),
    .Y(_02905_));
 sky130_fd_sc_hd__o211a_1 _16157_ (.A1(\core.pipe1_csrData[11] ),
    .A2(net641),
    .B1(_02905_),
    .C1(net1925),
    .X(_00518_));
 sky130_fd_sc_hd__nand2_1 _16158_ (.A(_02329_),
    .B(net642),
    .Y(_02906_));
 sky130_fd_sc_hd__o211a_1 _16159_ (.A1(\core.pipe1_csrData[12] ),
    .A2(net642),
    .B1(_02906_),
    .C1(net1920),
    .X(_00519_));
 sky130_fd_sc_hd__nand2_1 _16160_ (.A(_02352_),
    .B(net641),
    .Y(_02907_));
 sky130_fd_sc_hd__o211a_1 _16161_ (.A1(\core.pipe1_csrData[13] ),
    .A2(net641),
    .B1(_02907_),
    .C1(net1924),
    .X(_00520_));
 sky130_fd_sc_hd__nand2_1 _16162_ (.A(_02384_),
    .B(net641),
    .Y(_02908_));
 sky130_fd_sc_hd__o211a_1 _16163_ (.A1(\core.pipe1_csrData[14] ),
    .A2(net641),
    .B1(_02908_),
    .C1(net1924),
    .X(_00521_));
 sky130_fd_sc_hd__nand2_1 _16164_ (.A(_02415_),
    .B(net641),
    .Y(_02909_));
 sky130_fd_sc_hd__o211a_1 _16165_ (.A1(\core.pipe1_csrData[15] ),
    .A2(net641),
    .B1(_02909_),
    .C1(net1924),
    .X(_00522_));
 sky130_fd_sc_hd__nand2_1 _16166_ (.A(_02451_),
    .B(net640),
    .Y(_02910_));
 sky130_fd_sc_hd__o211a_1 _16167_ (.A1(\core.pipe1_csrData[16] ),
    .A2(net645),
    .B1(_02910_),
    .C1(net1908),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _16168_ (.A0(\core.pipe1_csrData[17] ),
    .A1(_02478_),
    .S(net645),
    .X(_02911_));
 sky130_fd_sc_hd__and2_1 _16169_ (.A(net1906),
    .B(_02911_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _16170_ (.A0(\core.pipe1_csrData[18] ),
    .A1(_02504_),
    .S(net645),
    .X(_02912_));
 sky130_fd_sc_hd__and2_1 _16171_ (.A(net1907),
    .B(_02912_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _16172_ (.A0(\core.pipe1_csrData[19] ),
    .A1(_02530_),
    .S(net640),
    .X(_02913_));
 sky130_fd_sc_hd__and2_1 _16173_ (.A(net1891),
    .B(_02913_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _16174_ (.A0(\core.pipe1_csrData[20] ),
    .A1(_02557_),
    .S(net640),
    .X(_02914_));
 sky130_fd_sc_hd__and2_1 _16175_ (.A(net1891),
    .B(_02914_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _16176_ (.A0(\core.pipe1_csrData[21] ),
    .A1(_02583_),
    .S(net640),
    .X(_02915_));
 sky130_fd_sc_hd__and2_1 _16177_ (.A(net1888),
    .B(_02915_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _16178_ (.A0(\core.pipe1_csrData[22] ),
    .A1(_02609_),
    .S(net642),
    .X(_02916_));
 sky130_fd_sc_hd__and2_1 _16179_ (.A(net1921),
    .B(_02916_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _16180_ (.A0(\core.pipe1_csrData[23] ),
    .A1(_02635_),
    .S(net640),
    .X(_02917_));
 sky130_fd_sc_hd__and2_1 _16181_ (.A(net1890),
    .B(_02917_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _16182_ (.A0(\core.pipe1_csrData[24] ),
    .A1(_02661_),
    .S(net640),
    .X(_02918_));
 sky130_fd_sc_hd__and2_1 _16183_ (.A(net1890),
    .B(_02918_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _16184_ (.A0(\core.pipe1_csrData[25] ),
    .A1(_02681_),
    .S(net640),
    .X(_02919_));
 sky130_fd_sc_hd__and2_1 _16185_ (.A(net1892),
    .B(_02919_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _16186_ (.A0(\core.pipe1_csrData[26] ),
    .A1(_02714_),
    .S(net640),
    .X(_02920_));
 sky130_fd_sc_hd__and2_1 _16187_ (.A(net1891),
    .B(_02920_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _16188_ (.A0(\core.pipe1_csrData[27] ),
    .A1(_02740_),
    .S(net640),
    .X(_02921_));
 sky130_fd_sc_hd__and2_1 _16189_ (.A(net1906),
    .B(_02921_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _16190_ (.A0(\core.pipe1_csrData[28] ),
    .A1(_02768_),
    .S(net640),
    .X(_02922_));
 sky130_fd_sc_hd__and2_1 _16191_ (.A(net1888),
    .B(_02922_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _16192_ (.A0(\core.pipe1_csrData[29] ),
    .A1(_02795_),
    .S(net643),
    .X(_02923_));
 sky130_fd_sc_hd__and2_1 _16193_ (.A(net1928),
    .B(_02923_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _16194_ (.A0(\core.pipe1_csrData[30] ),
    .A1(_02815_),
    .S(net644),
    .X(_02924_));
 sky130_fd_sc_hd__and2_1 _16195_ (.A(net1927),
    .B(_02924_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _16196_ (.A0(\core.pipe1_csrData[31] ),
    .A1(_02842_),
    .S(net643),
    .X(_02925_));
 sky130_fd_sc_hd__and2_1 _16197_ (.A(net1926),
    .B(_02925_),
    .X(_00538_));
 sky130_fd_sc_hd__nor2_1 _16198_ (.A(_04512_),
    .B(_09094_),
    .Y(_02926_));
 sky130_fd_sc_hd__and3_4 _16199_ (.A(net680),
    .B(net1075),
    .C(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__mux2_1 _16200_ (.A0(\core.registers[16][0] ),
    .A1(net1037),
    .S(net582),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _16201_ (.A0(\core.registers[16][1] ),
    .A1(net1040),
    .S(net582),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _16202_ (.A0(\core.registers[16][2] ),
    .A1(net1044),
    .S(net583),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _16203_ (.A0(\core.registers[16][3] ),
    .A1(net1048),
    .S(net582),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _16204_ (.A0(\core.registers[16][4] ),
    .A1(net1053),
    .S(net582),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _16205_ (.A0(\core.registers[16][5] ),
    .A1(net1057),
    .S(net583),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _16206_ (.A0(\core.registers[16][6] ),
    .A1(net1061),
    .S(net583),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _16207_ (.A0(\core.registers[16][7] ),
    .A1(net1133),
    .S(net583),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _16208_ (.A0(\core.registers[16][8] ),
    .A1(net959),
    .S(net583),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _16209_ (.A0(\core.registers[16][9] ),
    .A1(net964),
    .S(net581),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _16210_ (.A0(\core.registers[16][10] ),
    .A1(net969),
    .S(net582),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _16211_ (.A0(\core.registers[16][11] ),
    .A1(net972),
    .S(net581),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _16212_ (.A0(\core.registers[16][12] ),
    .A1(net989),
    .S(net582),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _16213_ (.A0(\core.registers[16][13] ),
    .A1(net986),
    .S(net583),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _16214_ (.A0(\core.registers[16][14] ),
    .A1(net975),
    .S(net582),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _16215_ (.A0(\core.registers[16][15] ),
    .A1(net981),
    .S(net582),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _16216_ (.A0(\core.registers[16][16] ),
    .A1(net1124),
    .S(net580),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _16217_ (.A0(\core.registers[16][17] ),
    .A1(net1128),
    .S(net580),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _16218_ (.A0(\core.registers[16][18] ),
    .A1(net1118),
    .S(net580),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _16219_ (.A0(\core.registers[16][19] ),
    .A1(net1120),
    .S(net580),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _16220_ (.A0(\core.registers[16][20] ),
    .A1(net1138),
    .S(net580),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _16221_ (.A0(\core.registers[16][21] ),
    .A1(net1143),
    .S(net580),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _16222_ (.A0(\core.registers[16][22] ),
    .A1(net1147),
    .S(net581),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _16223_ (.A0(\core.registers[16][23] ),
    .A1(net1151),
    .S(net580),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _16224_ (.A0(\core.registers[16][24] ),
    .A1(net1115),
    .S(net580),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _16225_ (.A0(\core.registers[16][25] ),
    .A1(net1109),
    .S(net580),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _16226_ (.A0(\core.registers[16][26] ),
    .A1(net1102),
    .S(net581),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _16227_ (.A0(\core.registers[16][27] ),
    .A1(net1106),
    .S(net581),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _16228_ (.A0(\core.registers[16][28] ),
    .A1(net1096),
    .S(net580),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _16229_ (.A0(\core.registers[16][29] ),
    .A1(net1092),
    .S(net582),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _16230_ (.A0(\core.registers[16][30] ),
    .A1(net1085),
    .S(net583),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _16231_ (.A0(\core.registers[16][31] ),
    .A1(net1089),
    .S(net582),
    .X(_00570_));
 sky130_fd_sc_hd__nor2_2 _16232_ (.A(net1970),
    .B(_08354_),
    .Y(_00611_));
 sky130_fd_sc_hd__and2b_1 _16233_ (.A_N(_08349_),
    .B(_08505_),
    .X(_02928_));
 sky130_fd_sc_hd__o21a_2 _16234_ (.A1(net725),
    .A2(_02928_),
    .B1(_00611_),
    .X(_00571_));
 sky130_fd_sc_hd__and2b_1 _16235_ (.A_N(_08349_),
    .B(_08506_),
    .X(_02929_));
 sky130_fd_sc_hd__o21a_4 _16236_ (.A1(net725),
    .A2(_02929_),
    .B1(_00611_),
    .X(_00572_));
 sky130_fd_sc_hd__and2b_1 _16237_ (.A_N(_08349_),
    .B(_08509_),
    .X(_02930_));
 sky130_fd_sc_hd__o21a_2 _16238_ (.A1(net725),
    .A2(_02930_),
    .B1(_00611_),
    .X(_00573_));
 sky130_fd_sc_hd__and2b_1 _16239_ (.A_N(_08349_),
    .B(_08510_),
    .X(_02931_));
 sky130_fd_sc_hd__o21a_2 _16240_ (.A1(net725),
    .A2(_02931_),
    .B1(_00611_),
    .X(_00574_));
 sky130_fd_sc_hd__nor2_1 _16241_ (.A(net1970),
    .B(_08153_),
    .Y(_00575_));
 sky130_fd_sc_hd__nor2_1 _16242_ (.A(net1990),
    .B(_08345_),
    .Y(_00576_));
 sky130_fd_sc_hd__or3_2 _16243_ (.A(\core.csr.currentInstruction[11] ),
    .B(_04424_),
    .C(_04514_),
    .X(_02932_));
 sky130_fd_sc_hd__nor2_1 _16244_ (.A(_04512_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__and3_2 _16245_ (.A(net675),
    .B(net1072),
    .C(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__mux2_1 _16246_ (.A0(\core.registers[12][0] ),
    .A1(net1035),
    .S(net578),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _16247_ (.A0(\core.registers[12][1] ),
    .A1(net1041),
    .S(net577),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _16248_ (.A0(\core.registers[12][2] ),
    .A1(net1043),
    .S(net577),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _16249_ (.A0(\core.registers[12][3] ),
    .A1(net1050),
    .S(net577),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _16250_ (.A0(\core.registers[12][4] ),
    .A1(net1055),
    .S(net577),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _16251_ (.A0(\core.registers[12][5] ),
    .A1(net1059),
    .S(net577),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _16252_ (.A0(\core.registers[12][6] ),
    .A1(net1064),
    .S(net577),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _16253_ (.A0(\core.registers[12][7] ),
    .A1(net1134),
    .S(net578),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _16254_ (.A0(\core.registers[12][8] ),
    .A1(net958),
    .S(net577),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _16255_ (.A0(\core.registers[12][9] ),
    .A1(net964),
    .S(net579),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _16256_ (.A0(\core.registers[12][10] ),
    .A1(net967),
    .S(net578),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _16257_ (.A0(\core.registers[12][11] ),
    .A1(net970),
    .S(net578),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _16258_ (.A0(\core.registers[12][12] ),
    .A1(net987),
    .S(net578),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _16259_ (.A0(\core.registers[12][13] ),
    .A1(net984),
    .S(net578),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _16260_ (.A0(\core.registers[12][14] ),
    .A1(net976),
    .S(net578),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _16261_ (.A0(\core.registers[12][15] ),
    .A1(net980),
    .S(net577),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _16262_ (.A0(\core.registers[12][16] ),
    .A1(net1124),
    .S(net576),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _16263_ (.A0(\core.registers[12][17] ),
    .A1(net1128),
    .S(net576),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _16264_ (.A0(\core.registers[12][18] ),
    .A1(net1116),
    .S(net579),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _16265_ (.A0(\core.registers[12][19] ),
    .A1(net1120),
    .S(net576),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _16266_ (.A0(\core.registers[12][20] ),
    .A1(net1136),
    .S(net576),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _16267_ (.A0(\core.registers[12][21] ),
    .A1(net1140),
    .S(net576),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _16268_ (.A0(\core.registers[12][22] ),
    .A1(net1146),
    .S(net579),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _16269_ (.A0(\core.registers[12][23] ),
    .A1(net1150),
    .S(net576),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _16270_ (.A0(\core.registers[12][24] ),
    .A1(net1112),
    .S(net576),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _16271_ (.A0(\core.registers[12][25] ),
    .A1(net1110),
    .S(net576),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _16272_ (.A0(\core.registers[12][26] ),
    .A1(net1101),
    .S(net579),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _16273_ (.A0(\core.registers[12][27] ),
    .A1(net1105),
    .S(net576),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _16274_ (.A0(\core.registers[12][28] ),
    .A1(net1096),
    .S(net576),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _16275_ (.A0(\core.registers[12][29] ),
    .A1(net1095),
    .S(net578),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _16276_ (.A0(\core.registers[12][30] ),
    .A1(net1086),
    .S(net577),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _16277_ (.A0(\core.registers[12][31] ),
    .A1(net1088),
    .S(net577),
    .X(_00609_));
 sky130_fd_sc_hd__nor2_1 _16278_ (.A(net284),
    .B(net375),
    .Y(_00610_));
 sky130_fd_sc_hd__nor3_4 _16279_ (.A(net1989),
    .B(net713),
    .C(_08375_),
    .Y(_00617_));
 sky130_fd_sc_hd__and3_1 _16280_ (.A(\wbSRAMInterface.currentByteSelect[0] ),
    .B(_07837_),
    .C(_00617_),
    .X(_00612_));
 sky130_fd_sc_hd__and3_1 _16281_ (.A(\wbSRAMInterface.currentByteSelect[1] ),
    .B(_07837_),
    .C(_00617_),
    .X(_00613_));
 sky130_fd_sc_hd__and3_1 _16282_ (.A(\wbSRAMInterface.currentByteSelect[2] ),
    .B(_07837_),
    .C(_00617_),
    .X(_00614_));
 sky130_fd_sc_hd__and3_1 _16283_ (.A(\wbSRAMInterface.currentByteSelect[3] ),
    .B(_07837_),
    .C(_00617_),
    .X(_00615_));
 sky130_fd_sc_hd__and3_1 _16284_ (.A(\wbSRAMInterface.currentAddress[11] ),
    .B(net2008),
    .C(_00617_),
    .X(_00616_));
 sky130_fd_sc_hd__nor2_1 _16285_ (.A(net1991),
    .B(\core.csr.cycleTimer.currentValue[0] ),
    .Y(_00618_));
 sky130_fd_sc_hd__a21oi_1 _16286_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(\core.csr.cycleTimer.currentValue[1] ),
    .B1(net1991),
    .Y(_02935_));
 sky130_fd_sc_hd__o21a_1 _16287_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(\core.csr.cycleTimer.currentValue[1] ),
    .B1(_02935_),
    .X(_00619_));
 sky130_fd_sc_hd__a21oi_1 _16288_ (.A1(\core.csr.cycleTimer.currentValue[0] ),
    .A2(\core.csr.cycleTimer.currentValue[1] ),
    .B1(\core.csr.cycleTimer.currentValue[2] ),
    .Y(_02936_));
 sky130_fd_sc_hd__and3_2 _16289_ (.A(\core.csr.cycleTimer.currentValue[0] ),
    .B(\core.csr.cycleTimer.currentValue[1] ),
    .C(\core.csr.cycleTimer.currentValue[2] ),
    .X(_02937_));
 sky130_fd_sc_hd__nor3_1 _16290_ (.A(net1991),
    .B(_02936_),
    .C(_02937_),
    .Y(_00620_));
 sky130_fd_sc_hd__and2_1 _16291_ (.A(\core.csr.cycleTimer.currentValue[3] ),
    .B(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__o21ai_1 _16292_ (.A1(\core.csr.cycleTimer.currentValue[3] ),
    .A2(_02937_),
    .B1(net1952),
    .Y(_02939_));
 sky130_fd_sc_hd__nor2_1 _16293_ (.A(_02938_),
    .B(_02939_),
    .Y(_00621_));
 sky130_fd_sc_hd__and3_2 _16294_ (.A(\core.csr.cycleTimer.currentValue[3] ),
    .B(\core.csr.cycleTimer.currentValue[4] ),
    .C(_02937_),
    .X(_02940_));
 sky130_fd_sc_hd__o21ai_1 _16295_ (.A1(\core.csr.cycleTimer.currentValue[4] ),
    .A2(_02938_),
    .B1(net1952),
    .Y(_02941_));
 sky130_fd_sc_hd__nor2_1 _16296_ (.A(_02940_),
    .B(_02941_),
    .Y(_00622_));
 sky130_fd_sc_hd__and2_1 _16297_ (.A(\core.csr.cycleTimer.currentValue[5] ),
    .B(_02940_),
    .X(_02942_));
 sky130_fd_sc_hd__nor2_1 _16298_ (.A(net1992),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__o21a_1 _16299_ (.A1(\core.csr.cycleTimer.currentValue[5] ),
    .A2(_02940_),
    .B1(_02943_),
    .X(_00623_));
 sky130_fd_sc_hd__and3_2 _16300_ (.A(\core.csr.cycleTimer.currentValue[5] ),
    .B(\core.csr.cycleTimer.currentValue[6] ),
    .C(_02940_),
    .X(_02944_));
 sky130_fd_sc_hd__o21ai_1 _16301_ (.A1(\core.csr.cycleTimer.currentValue[6] ),
    .A2(_02942_),
    .B1(net1958),
    .Y(_02945_));
 sky130_fd_sc_hd__nor2_1 _16302_ (.A(_02944_),
    .B(_02945_),
    .Y(_00624_));
 sky130_fd_sc_hd__a21oi_1 _16303_ (.A1(\core.csr.cycleTimer.currentValue[7] ),
    .A2(_02944_),
    .B1(net1991),
    .Y(_02946_));
 sky130_fd_sc_hd__o21a_1 _16304_ (.A1(\core.csr.cycleTimer.currentValue[7] ),
    .A2(_02944_),
    .B1(_02946_),
    .X(_00625_));
 sky130_fd_sc_hd__a21oi_1 _16305_ (.A1(\core.csr.cycleTimer.currentValue[7] ),
    .A2(_02944_),
    .B1(\core.csr.cycleTimer.currentValue[8] ),
    .Y(_02947_));
 sky130_fd_sc_hd__and3_1 _16306_ (.A(\core.csr.cycleTimer.currentValue[7] ),
    .B(\core.csr.cycleTimer.currentValue[8] ),
    .C(_02944_),
    .X(_02948_));
 sky130_fd_sc_hd__nor3_1 _16307_ (.A(net1991),
    .B(_02947_),
    .C(_02948_),
    .Y(_00626_));
 sky130_fd_sc_hd__and2_2 _16308_ (.A(\core.csr.cycleTimer.currentValue[9] ),
    .B(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__o21ai_1 _16309_ (.A1(\core.csr.cycleTimer.currentValue[9] ),
    .A2(_02948_),
    .B1(net1958),
    .Y(_02950_));
 sky130_fd_sc_hd__nor2_1 _16310_ (.A(_02949_),
    .B(_02950_),
    .Y(_00627_));
 sky130_fd_sc_hd__a21oi_1 _16311_ (.A1(\core.csr.cycleTimer.currentValue[10] ),
    .A2(_02949_),
    .B1(net1998),
    .Y(_02951_));
 sky130_fd_sc_hd__o21a_1 _16312_ (.A1(\core.csr.cycleTimer.currentValue[10] ),
    .A2(_02949_),
    .B1(_02951_),
    .X(_00628_));
 sky130_fd_sc_hd__a21oi_1 _16313_ (.A1(\core.csr.cycleTimer.currentValue[10] ),
    .A2(_02949_),
    .B1(\core.csr.cycleTimer.currentValue[11] ),
    .Y(_02952_));
 sky130_fd_sc_hd__and3_1 _16314_ (.A(\core.csr.cycleTimer.currentValue[10] ),
    .B(\core.csr.cycleTimer.currentValue[11] ),
    .C(_02949_),
    .X(_02953_));
 sky130_fd_sc_hd__nor3_1 _16315_ (.A(net1998),
    .B(_02952_),
    .C(_02953_),
    .Y(_00629_));
 sky130_fd_sc_hd__and2_2 _16316_ (.A(\core.csr.cycleTimer.currentValue[12] ),
    .B(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__o21ai_1 _16317_ (.A1(\core.csr.cycleTimer.currentValue[12] ),
    .A2(_02953_),
    .B1(net1958),
    .Y(_02955_));
 sky130_fd_sc_hd__nor2_1 _16318_ (.A(_02954_),
    .B(_02955_),
    .Y(_00630_));
 sky130_fd_sc_hd__a21oi_1 _16319_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(_02954_),
    .B1(net1998),
    .Y(_02956_));
 sky130_fd_sc_hd__o21a_1 _16320_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(_02954_),
    .B1(_02956_),
    .X(_00631_));
 sky130_fd_sc_hd__a21oi_1 _16321_ (.A1(\core.csr.cycleTimer.currentValue[13] ),
    .A2(_02954_),
    .B1(\core.csr.cycleTimer.currentValue[14] ),
    .Y(_02957_));
 sky130_fd_sc_hd__and3_1 _16322_ (.A(\core.csr.cycleTimer.currentValue[13] ),
    .B(\core.csr.cycleTimer.currentValue[14] ),
    .C(_02954_),
    .X(_02958_));
 sky130_fd_sc_hd__nor3_1 _16323_ (.A(net1998),
    .B(_02957_),
    .C(_02958_),
    .Y(_00632_));
 sky130_fd_sc_hd__and2_4 _16324_ (.A(\core.csr.cycleTimer.currentValue[15] ),
    .B(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__o21ai_1 _16325_ (.A1(\core.csr.cycleTimer.currentValue[15] ),
    .A2(_02958_),
    .B1(net1955),
    .Y(_02960_));
 sky130_fd_sc_hd__nor2_1 _16326_ (.A(_02959_),
    .B(_02960_),
    .Y(_00633_));
 sky130_fd_sc_hd__a21oi_1 _16327_ (.A1(\core.csr.cycleTimer.currentValue[16] ),
    .A2(_02959_),
    .B1(net1985),
    .Y(_02961_));
 sky130_fd_sc_hd__o21a_1 _16328_ (.A1(\core.csr.cycleTimer.currentValue[16] ),
    .A2(_02959_),
    .B1(_02961_),
    .X(_00634_));
 sky130_fd_sc_hd__a21oi_1 _16329_ (.A1(\core.csr.cycleTimer.currentValue[16] ),
    .A2(_02959_),
    .B1(\core.csr.cycleTimer.currentValue[17] ),
    .Y(_02962_));
 sky130_fd_sc_hd__and3_2 _16330_ (.A(\core.csr.cycleTimer.currentValue[16] ),
    .B(\core.csr.cycleTimer.currentValue[17] ),
    .C(_02959_),
    .X(_02963_));
 sky130_fd_sc_hd__nor3_1 _16331_ (.A(net1981),
    .B(_02962_),
    .C(_02963_),
    .Y(_00635_));
 sky130_fd_sc_hd__and2_2 _16332_ (.A(\core.csr.cycleTimer.currentValue[18] ),
    .B(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__o21ai_1 _16333_ (.A1(\core.csr.cycleTimer.currentValue[18] ),
    .A2(_02963_),
    .B1(net1916),
    .Y(_02965_));
 sky130_fd_sc_hd__nor2_1 _16334_ (.A(_02964_),
    .B(_02965_),
    .Y(_00636_));
 sky130_fd_sc_hd__a21oi_1 _16335_ (.A1(\core.csr.cycleTimer.currentValue[19] ),
    .A2(_02964_),
    .B1(net1976),
    .Y(_02966_));
 sky130_fd_sc_hd__o21a_1 _16336_ (.A1(\core.csr.cycleTimer.currentValue[19] ),
    .A2(_02964_),
    .B1(_02966_),
    .X(_00637_));
 sky130_fd_sc_hd__a21oi_1 _16337_ (.A1(\core.csr.cycleTimer.currentValue[19] ),
    .A2(_02964_),
    .B1(\core.csr.cycleTimer.currentValue[20] ),
    .Y(_02967_));
 sky130_fd_sc_hd__and3_1 _16338_ (.A(\core.csr.cycleTimer.currentValue[19] ),
    .B(\core.csr.cycleTimer.currentValue[20] ),
    .C(_02964_),
    .X(_02968_));
 sky130_fd_sc_hd__nor3_1 _16339_ (.A(net1976),
    .B(_02967_),
    .C(_02968_),
    .Y(_00638_));
 sky130_fd_sc_hd__and2_2 _16340_ (.A(\core.csr.cycleTimer.currentValue[21] ),
    .B(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__o21ai_1 _16341_ (.A1(\core.csr.cycleTimer.currentValue[21] ),
    .A2(_02968_),
    .B1(net1916),
    .Y(_02970_));
 sky130_fd_sc_hd__nor2_1 _16342_ (.A(_02969_),
    .B(_02970_),
    .Y(_00639_));
 sky130_fd_sc_hd__a21oi_1 _16343_ (.A1(\core.csr.cycleTimer.currentValue[22] ),
    .A2(_02969_),
    .B1(net1976),
    .Y(_02971_));
 sky130_fd_sc_hd__o21a_1 _16344_ (.A1(\core.csr.cycleTimer.currentValue[22] ),
    .A2(_02969_),
    .B1(_02971_),
    .X(_00640_));
 sky130_fd_sc_hd__a21oi_1 _16345_ (.A1(\core.csr.cycleTimer.currentValue[22] ),
    .A2(_02969_),
    .B1(\core.csr.cycleTimer.currentValue[23] ),
    .Y(_02972_));
 sky130_fd_sc_hd__and3_1 _16346_ (.A(\core.csr.cycleTimer.currentValue[22] ),
    .B(\core.csr.cycleTimer.currentValue[23] ),
    .C(_02969_),
    .X(_02973_));
 sky130_fd_sc_hd__nor3_1 _16347_ (.A(net1976),
    .B(_02972_),
    .C(_02973_),
    .Y(_00641_));
 sky130_fd_sc_hd__and2_2 _16348_ (.A(\core.csr.cycleTimer.currentValue[24] ),
    .B(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__o21ai_1 _16349_ (.A1(\core.csr.cycleTimer.currentValue[24] ),
    .A2(_02973_),
    .B1(net1916),
    .Y(_02975_));
 sky130_fd_sc_hd__nor2_1 _16350_ (.A(_02974_),
    .B(_02975_),
    .Y(_00642_));
 sky130_fd_sc_hd__a21oi_1 _16351_ (.A1(\core.csr.cycleTimer.currentValue[25] ),
    .A2(_02974_),
    .B1(net1977),
    .Y(_02976_));
 sky130_fd_sc_hd__o21a_1 _16352_ (.A1(\core.csr.cycleTimer.currentValue[25] ),
    .A2(_02974_),
    .B1(_02976_),
    .X(_00643_));
 sky130_fd_sc_hd__a21oi_1 _16353_ (.A1(\core.csr.cycleTimer.currentValue[25] ),
    .A2(_02974_),
    .B1(\core.csr.cycleTimer.currentValue[26] ),
    .Y(_02977_));
 sky130_fd_sc_hd__and3_1 _16354_ (.A(\core.csr.cycleTimer.currentValue[25] ),
    .B(\core.csr.cycleTimer.currentValue[26] ),
    .C(_02974_),
    .X(_02978_));
 sky130_fd_sc_hd__nor3_1 _16355_ (.A(net1977),
    .B(_02977_),
    .C(_02978_),
    .Y(_00644_));
 sky130_fd_sc_hd__and2_2 _16356_ (.A(\core.csr.cycleTimer.currentValue[27] ),
    .B(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__o21ai_1 _16357_ (.A1(\core.csr.cycleTimer.currentValue[27] ),
    .A2(_02978_),
    .B1(net1917),
    .Y(_02980_));
 sky130_fd_sc_hd__nor2_1 _16358_ (.A(_02979_),
    .B(_02980_),
    .Y(_00645_));
 sky130_fd_sc_hd__a21oi_1 _16359_ (.A1(\core.csr.cycleTimer.currentValue[28] ),
    .A2(_02979_),
    .B1(net1977),
    .Y(_02981_));
 sky130_fd_sc_hd__o21a_1 _16360_ (.A1(\core.csr.cycleTimer.currentValue[28] ),
    .A2(_02979_),
    .B1(_02981_),
    .X(_00646_));
 sky130_fd_sc_hd__a21oi_1 _16361_ (.A1(\core.csr.cycleTimer.currentValue[28] ),
    .A2(_02979_),
    .B1(\core.csr.cycleTimer.currentValue[29] ),
    .Y(_02982_));
 sky130_fd_sc_hd__and3_4 _16362_ (.A(\core.csr.cycleTimer.currentValue[28] ),
    .B(\core.csr.cycleTimer.currentValue[29] ),
    .C(_02979_),
    .X(_02983_));
 sky130_fd_sc_hd__nor3_1 _16363_ (.A(net1981),
    .B(_02982_),
    .C(_02983_),
    .Y(_00647_));
 sky130_fd_sc_hd__and2_2 _16364_ (.A(\core.csr.cycleTimer.currentValue[30] ),
    .B(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__o21ai_1 _16365_ (.A1(\core.csr.cycleTimer.currentValue[30] ),
    .A2(_02983_),
    .B1(net1937),
    .Y(_02985_));
 sky130_fd_sc_hd__nor2_1 _16366_ (.A(_02984_),
    .B(_02985_),
    .Y(_00648_));
 sky130_fd_sc_hd__a21oi_1 _16367_ (.A1(\core.csr.cycleTimer.currentValue[31] ),
    .A2(_02984_),
    .B1(net1995),
    .Y(_02986_));
 sky130_fd_sc_hd__o21a_1 _16368_ (.A1(\core.csr.cycleTimer.currentValue[31] ),
    .A2(_02984_),
    .B1(_02986_),
    .X(_00649_));
 sky130_fd_sc_hd__a21oi_1 _16369_ (.A1(\core.csr.cycleTimer.currentValue[31] ),
    .A2(_02984_),
    .B1(\core.csr.cycleTimer.currentValue[32] ),
    .Y(_02987_));
 sky130_fd_sc_hd__and3_2 _16370_ (.A(\core.csr.cycleTimer.currentValue[32] ),
    .B(\core.csr.cycleTimer.currentValue[31] ),
    .C(_02984_),
    .X(_02988_));
 sky130_fd_sc_hd__nor3_1 _16371_ (.A(net1995),
    .B(_02987_),
    .C(_02988_),
    .Y(_00650_));
 sky130_fd_sc_hd__and2_2 _16372_ (.A(\core.csr.cycleTimer.currentValue[33] ),
    .B(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__o21ai_1 _16373_ (.A1(\core.csr.cycleTimer.currentValue[33] ),
    .A2(_02988_),
    .B1(net1945),
    .Y(_02990_));
 sky130_fd_sc_hd__nor2_1 _16374_ (.A(_02989_),
    .B(_02990_),
    .Y(_00651_));
 sky130_fd_sc_hd__a21oi_1 _16375_ (.A1(\core.csr.cycleTimer.currentValue[34] ),
    .A2(_02989_),
    .B1(net1991),
    .Y(_02991_));
 sky130_fd_sc_hd__o21a_1 _16376_ (.A1(\core.csr.cycleTimer.currentValue[34] ),
    .A2(_02989_),
    .B1(_02991_),
    .X(_00652_));
 sky130_fd_sc_hd__a21oi_1 _16377_ (.A1(\core.csr.cycleTimer.currentValue[34] ),
    .A2(_02989_),
    .B1(\core.csr.cycleTimer.currentValue[35] ),
    .Y(_02992_));
 sky130_fd_sc_hd__and3_1 _16378_ (.A(\core.csr.cycleTimer.currentValue[34] ),
    .B(\core.csr.cycleTimer.currentValue[35] ),
    .C(_02989_),
    .X(_02993_));
 sky130_fd_sc_hd__nor3_1 _16379_ (.A(net1991),
    .B(_02992_),
    .C(_02993_),
    .Y(_00653_));
 sky130_fd_sc_hd__and2_2 _16380_ (.A(\core.csr.cycleTimer.currentValue[36] ),
    .B(_02993_),
    .X(_02994_));
 sky130_fd_sc_hd__o21ai_1 _16381_ (.A1(\core.csr.cycleTimer.currentValue[36] ),
    .A2(_02993_),
    .B1(net1952),
    .Y(_02995_));
 sky130_fd_sc_hd__nor2_1 _16382_ (.A(_02994_),
    .B(_02995_),
    .Y(_00654_));
 sky130_fd_sc_hd__a21oi_1 _16383_ (.A1(\core.csr.cycleTimer.currentValue[37] ),
    .A2(_02994_),
    .B1(net1993),
    .Y(_02996_));
 sky130_fd_sc_hd__o21a_1 _16384_ (.A1(\core.csr.cycleTimer.currentValue[37] ),
    .A2(_02994_),
    .B1(_02996_),
    .X(_00655_));
 sky130_fd_sc_hd__a21oi_1 _16385_ (.A1(\core.csr.cycleTimer.currentValue[37] ),
    .A2(_02994_),
    .B1(\core.csr.cycleTimer.currentValue[38] ),
    .Y(_02997_));
 sky130_fd_sc_hd__and3_1 _16386_ (.A(\core.csr.cycleTimer.currentValue[37] ),
    .B(\core.csr.cycleTimer.currentValue[38] ),
    .C(_02994_),
    .X(_02998_));
 sky130_fd_sc_hd__nor3_1 _16387_ (.A(net1992),
    .B(_02997_),
    .C(_02998_),
    .Y(_00656_));
 sky130_fd_sc_hd__and2_2 _16388_ (.A(\core.csr.cycleTimer.currentValue[39] ),
    .B(_02998_),
    .X(_02999_));
 sky130_fd_sc_hd__nor2_1 _16389_ (.A(net1992),
    .B(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__o21a_1 _16390_ (.A1(\core.csr.cycleTimer.currentValue[39] ),
    .A2(_02998_),
    .B1(_03000_),
    .X(_00657_));
 sky130_fd_sc_hd__a21oi_1 _16391_ (.A1(\core.csr.cycleTimer.currentValue[40] ),
    .A2(_02999_),
    .B1(net1992),
    .Y(_03001_));
 sky130_fd_sc_hd__o21a_1 _16392_ (.A1(\core.csr.cycleTimer.currentValue[40] ),
    .A2(_02999_),
    .B1(_03001_),
    .X(_00658_));
 sky130_fd_sc_hd__a21oi_1 _16393_ (.A1(\core.csr.cycleTimer.currentValue[40] ),
    .A2(_02999_),
    .B1(\core.csr.cycleTimer.currentValue[41] ),
    .Y(_03002_));
 sky130_fd_sc_hd__and3_1 _16394_ (.A(\core.csr.cycleTimer.currentValue[40] ),
    .B(\core.csr.cycleTimer.currentValue[41] ),
    .C(_02999_),
    .X(_03003_));
 sky130_fd_sc_hd__nor3_1 _16395_ (.A(net1992),
    .B(_03002_),
    .C(_03003_),
    .Y(_00659_));
 sky130_fd_sc_hd__and2_2 _16396_ (.A(\core.csr.cycleTimer.currentValue[42] ),
    .B(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__nor2_1 _16397_ (.A(net1997),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__o21a_1 _16398_ (.A1(\core.csr.cycleTimer.currentValue[42] ),
    .A2(_03003_),
    .B1(_03005_),
    .X(_00660_));
 sky130_fd_sc_hd__a21oi_1 _16399_ (.A1(\core.csr.cycleTimer.currentValue[43] ),
    .A2(_03004_),
    .B1(net1998),
    .Y(_03006_));
 sky130_fd_sc_hd__o21a_1 _16400_ (.A1(\core.csr.cycleTimer.currentValue[43] ),
    .A2(_03004_),
    .B1(_03006_),
    .X(_00661_));
 sky130_fd_sc_hd__a21oi_1 _16401_ (.A1(\core.csr.cycleTimer.currentValue[43] ),
    .A2(_03004_),
    .B1(\core.csr.cycleTimer.currentValue[44] ),
    .Y(_03007_));
 sky130_fd_sc_hd__and3_1 _16402_ (.A(\core.csr.cycleTimer.currentValue[43] ),
    .B(\core.csr.cycleTimer.currentValue[44] ),
    .C(_03004_),
    .X(_03008_));
 sky130_fd_sc_hd__nor3_1 _16403_ (.A(net1998),
    .B(_03007_),
    .C(_03008_),
    .Y(_00662_));
 sky130_fd_sc_hd__and2_2 _16404_ (.A(\core.csr.cycleTimer.currentValue[45] ),
    .B(_03008_),
    .X(_03009_));
 sky130_fd_sc_hd__nor2_1 _16405_ (.A(net1998),
    .B(_03009_),
    .Y(_03010_));
 sky130_fd_sc_hd__o21a_1 _16406_ (.A1(\core.csr.cycleTimer.currentValue[45] ),
    .A2(_03008_),
    .B1(_03010_),
    .X(_00663_));
 sky130_fd_sc_hd__a21oi_1 _16407_ (.A1(\core.csr.cycleTimer.currentValue[46] ),
    .A2(_03009_),
    .B1(net1999),
    .Y(_03011_));
 sky130_fd_sc_hd__o21a_1 _16408_ (.A1(\core.csr.cycleTimer.currentValue[46] ),
    .A2(_03009_),
    .B1(_03011_),
    .X(_00664_));
 sky130_fd_sc_hd__a21oi_1 _16409_ (.A1(\core.csr.cycleTimer.currentValue[46] ),
    .A2(_03009_),
    .B1(\core.csr.cycleTimer.currentValue[47] ),
    .Y(_03012_));
 sky130_fd_sc_hd__and3_4 _16410_ (.A(\core.csr.cycleTimer.currentValue[46] ),
    .B(\core.csr.cycleTimer.currentValue[47] ),
    .C(_03009_),
    .X(_03013_));
 sky130_fd_sc_hd__nor3_1 _16411_ (.A(net1999),
    .B(_03012_),
    .C(_03013_),
    .Y(_00665_));
 sky130_fd_sc_hd__and2_2 _16412_ (.A(\core.csr.cycleTimer.currentValue[48] ),
    .B(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__nor2_1 _16413_ (.A(net1985),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__o21a_1 _16414_ (.A1(\core.csr.cycleTimer.currentValue[48] ),
    .A2(_03013_),
    .B1(_03015_),
    .X(_00666_));
 sky130_fd_sc_hd__a21oi_1 _16415_ (.A1(\core.csr.cycleTimer.currentValue[49] ),
    .A2(_03014_),
    .B1(net1981),
    .Y(_03016_));
 sky130_fd_sc_hd__o21a_1 _16416_ (.A1(\core.csr.cycleTimer.currentValue[49] ),
    .A2(_03014_),
    .B1(_03016_),
    .X(_00667_));
 sky130_fd_sc_hd__a21oi_1 _16417_ (.A1(\core.csr.cycleTimer.currentValue[49] ),
    .A2(_03014_),
    .B1(\core.csr.cycleTimer.currentValue[50] ),
    .Y(_03017_));
 sky130_fd_sc_hd__and3_4 _16418_ (.A(\core.csr.cycleTimer.currentValue[49] ),
    .B(\core.csr.cycleTimer.currentValue[50] ),
    .C(_03014_),
    .X(_03018_));
 sky130_fd_sc_hd__nor3_1 _16419_ (.A(net1981),
    .B(_03017_),
    .C(_03018_),
    .Y(_00668_));
 sky130_fd_sc_hd__and2_2 _16420_ (.A(\core.csr.cycleTimer.currentValue[51] ),
    .B(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__nor2_1 _16421_ (.A(net1972),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__o21a_1 _16422_ (.A1(\core.csr.cycleTimer.currentValue[51] ),
    .A2(_03018_),
    .B1(_03020_),
    .X(_00669_));
 sky130_fd_sc_hd__a21oi_1 _16423_ (.A1(\core.csr.cycleTimer.currentValue[52] ),
    .A2(_03019_),
    .B1(net1972),
    .Y(_03021_));
 sky130_fd_sc_hd__o21a_1 _16424_ (.A1(\core.csr.cycleTimer.currentValue[52] ),
    .A2(_03019_),
    .B1(_03021_),
    .X(_00670_));
 sky130_fd_sc_hd__a21oi_1 _16425_ (.A1(\core.csr.cycleTimer.currentValue[52] ),
    .A2(_03019_),
    .B1(\core.csr.cycleTimer.currentValue[53] ),
    .Y(_03022_));
 sky130_fd_sc_hd__and3_1 _16426_ (.A(\core.csr.cycleTimer.currentValue[52] ),
    .B(\core.csr.cycleTimer.currentValue[53] ),
    .C(_03019_),
    .X(_03023_));
 sky130_fd_sc_hd__nor3_1 _16427_ (.A(net1973),
    .B(_03022_),
    .C(_03023_),
    .Y(_00671_));
 sky130_fd_sc_hd__and2_2 _16428_ (.A(\core.csr.cycleTimer.currentValue[54] ),
    .B(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__nor2_1 _16429_ (.A(net1973),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__o21a_1 _16430_ (.A1(\core.csr.cycleTimer.currentValue[54] ),
    .A2(_03023_),
    .B1(_03025_),
    .X(_00672_));
 sky130_fd_sc_hd__a21oi_1 _16431_ (.A1(\core.csr.cycleTimer.currentValue[55] ),
    .A2(_03024_),
    .B1(net1976),
    .Y(_03026_));
 sky130_fd_sc_hd__o21a_1 _16432_ (.A1(\core.csr.cycleTimer.currentValue[55] ),
    .A2(_03024_),
    .B1(_03026_),
    .X(_00673_));
 sky130_fd_sc_hd__a21oi_1 _16433_ (.A1(\core.csr.cycleTimer.currentValue[55] ),
    .A2(_03024_),
    .B1(\core.csr.cycleTimer.currentValue[56] ),
    .Y(_03027_));
 sky130_fd_sc_hd__and3_1 _16434_ (.A(\core.csr.cycleTimer.currentValue[55] ),
    .B(\core.csr.cycleTimer.currentValue[56] ),
    .C(_03024_),
    .X(_03028_));
 sky130_fd_sc_hd__nor3_1 _16435_ (.A(net1976),
    .B(_03027_),
    .C(_03028_),
    .Y(_00674_));
 sky130_fd_sc_hd__nor2_1 _16436_ (.A(\core.csr.cycleTimer.currentValue[57] ),
    .B(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__and2_2 _16437_ (.A(\core.csr.cycleTimer.currentValue[57] ),
    .B(_03028_),
    .X(_03030_));
 sky130_fd_sc_hd__nor3_1 _16438_ (.A(net1976),
    .B(_03029_),
    .C(_03030_),
    .Y(_00675_));
 sky130_fd_sc_hd__a21oi_1 _16439_ (.A1(\core.csr.cycleTimer.currentValue[58] ),
    .A2(_03030_),
    .B1(net1977),
    .Y(_03031_));
 sky130_fd_sc_hd__o21a_1 _16440_ (.A1(\core.csr.cycleTimer.currentValue[58] ),
    .A2(_03030_),
    .B1(_03031_),
    .X(_00676_));
 sky130_fd_sc_hd__a21oi_1 _16441_ (.A1(\core.csr.cycleTimer.currentValue[58] ),
    .A2(_03030_),
    .B1(\core.csr.cycleTimer.currentValue[59] ),
    .Y(_03032_));
 sky130_fd_sc_hd__and3_1 _16442_ (.A(\core.csr.cycleTimer.currentValue[58] ),
    .B(\core.csr.cycleTimer.currentValue[59] ),
    .C(_03030_),
    .X(_03033_));
 sky130_fd_sc_hd__nor3_1 _16443_ (.A(net1977),
    .B(_03032_),
    .C(_03033_),
    .Y(_00677_));
 sky130_fd_sc_hd__and2_4 _16444_ (.A(\core.csr.cycleTimer.currentValue[60] ),
    .B(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__nor2_1 _16445_ (.A(net1977),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__o21a_1 _16446_ (.A1(\core.csr.cycleTimer.currentValue[60] ),
    .A2(_03033_),
    .B1(_03035_),
    .X(_00678_));
 sky130_fd_sc_hd__a21oi_1 _16447_ (.A1(\core.csr.cycleTimer.currentValue[61] ),
    .A2(_03034_),
    .B1(net1982),
    .Y(_03036_));
 sky130_fd_sc_hd__o21a_1 _16448_ (.A1(\core.csr.cycleTimer.currentValue[61] ),
    .A2(_03034_),
    .B1(_03036_),
    .X(_00679_));
 sky130_fd_sc_hd__a21oi_1 _16449_ (.A1(\core.csr.cycleTimer.currentValue[61] ),
    .A2(_03034_),
    .B1(\core.csr.cycleTimer.currentValue[62] ),
    .Y(_03037_));
 sky130_fd_sc_hd__and3_1 _16450_ (.A(\core.csr.cycleTimer.currentValue[61] ),
    .B(\core.csr.cycleTimer.currentValue[62] ),
    .C(_03034_),
    .X(_03038_));
 sky130_fd_sc_hd__nor3_1 _16451_ (.A(net1985),
    .B(_03037_),
    .C(_03038_),
    .Y(_00680_));
 sky130_fd_sc_hd__a21oi_1 _16452_ (.A1(\core.csr.cycleTimer.currentValue[63] ),
    .A2(_03038_),
    .B1(net1985),
    .Y(_03039_));
 sky130_fd_sc_hd__o21a_1 _16453_ (.A1(\core.csr.cycleTimer.currentValue[63] ),
    .A2(_03038_),
    .B1(_03039_),
    .X(_00681_));
 sky130_fd_sc_hd__nand2_4 _16454_ (.A(_04510_),
    .B(_04511_),
    .Y(_03040_));
 sky130_fd_sc_hd__nor2_1 _16455_ (.A(_09105_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__and3_4 _16456_ (.A(net680),
    .B(net1075),
    .C(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__mux2_1 _16457_ (.A0(\core.registers[25][0] ),
    .A1(net1036),
    .S(net575),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _16458_ (.A0(\core.registers[25][1] ),
    .A1(net1041),
    .S(net574),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _16459_ (.A0(\core.registers[25][2] ),
    .A1(net1043),
    .S(net574),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _16460_ (.A0(\core.registers[25][3] ),
    .A1(net1051),
    .S(net575),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _16461_ (.A0(\core.registers[25][4] ),
    .A1(net1055),
    .S(net575),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _16462_ (.A0(\core.registers[25][5] ),
    .A1(net1058),
    .S(net575),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _16463_ (.A0(\core.registers[25][6] ),
    .A1(net1061),
    .S(net574),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _16464_ (.A0(\core.registers[25][7] ),
    .A1(net1132),
    .S(net574),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _16465_ (.A0(\core.registers[25][8] ),
    .A1(net957),
    .S(net574),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _16466_ (.A0(\core.registers[25][9] ),
    .A1(net962),
    .S(net573),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _16467_ (.A0(\core.registers[25][10] ),
    .A1(net966),
    .S(net575),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _16468_ (.A0(\core.registers[25][11] ),
    .A1(net971),
    .S(net575),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _16469_ (.A0(\core.registers[25][12] ),
    .A1(net987),
    .S(net573),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _16470_ (.A0(\core.registers[25][13] ),
    .A1(net983),
    .S(net574),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _16471_ (.A0(\core.registers[25][14] ),
    .A1(net976),
    .S(net575),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _16472_ (.A0(\core.registers[25][15] ),
    .A1(net979),
    .S(net574),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _16473_ (.A0(\core.registers[25][16] ),
    .A1(net1127),
    .S(net572),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _16474_ (.A0(\core.registers[25][17] ),
    .A1(net1131),
    .S(net572),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _16475_ (.A0(\core.registers[25][18] ),
    .A1(net1117),
    .S(net573),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _16476_ (.A0(\core.registers[25][19] ),
    .A1(net1121),
    .S(net572),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _16477_ (.A0(\core.registers[25][20] ),
    .A1(net1137),
    .S(net572),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _16478_ (.A0(\core.registers[25][21] ),
    .A1(net1140),
    .S(net572),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _16479_ (.A0(\core.registers[25][22] ),
    .A1(net1145),
    .S(net573),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _16480_ (.A0(\core.registers[25][23] ),
    .A1(net1149),
    .S(net572),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _16481_ (.A0(\core.registers[25][24] ),
    .A1(net1112),
    .S(net572),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _16482_ (.A0(\core.registers[25][25] ),
    .A1(net1108),
    .S(net572),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _16483_ (.A0(\core.registers[25][26] ),
    .A1(net1100),
    .S(net573),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _16484_ (.A0(\core.registers[25][27] ),
    .A1(net1104),
    .S(net572),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _16485_ (.A0(\core.registers[25][28] ),
    .A1(net1098),
    .S(net572),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _16486_ (.A0(\core.registers[25][29] ),
    .A1(net1094),
    .S(net574),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _16487_ (.A0(\core.registers[25][30] ),
    .A1(net1084),
    .S(net574),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _16488_ (.A0(\core.registers[25][31] ),
    .A1(net1088),
    .S(net574),
    .X(_00713_));
 sky130_fd_sc_hd__nor2_1 _16489_ (.A(_09094_),
    .B(_09097_),
    .Y(_03043_));
 sky130_fd_sc_hd__and3_4 _16490_ (.A(net679),
    .B(net1075),
    .C(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__mux2_1 _16491_ (.A0(\core.registers[18][0] ),
    .A1(net1037),
    .S(net570),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _16492_ (.A0(\core.registers[18][1] ),
    .A1(net1040),
    .S(net570),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _16493_ (.A0(\core.registers[18][2] ),
    .A1(net1044),
    .S(net570),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _16494_ (.A0(\core.registers[18][3] ),
    .A1(net1048),
    .S(net570),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _16495_ (.A0(\core.registers[18][4] ),
    .A1(net1053),
    .S(net570),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _16496_ (.A0(\core.registers[18][5] ),
    .A1(net1057),
    .S(net571),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _16497_ (.A0(\core.registers[18][6] ),
    .A1(net1062),
    .S(net571),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _16498_ (.A0(\core.registers[18][7] ),
    .A1(net1133),
    .S(net571),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _16499_ (.A0(\core.registers[18][8] ),
    .A1(net960),
    .S(net571),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _16500_ (.A0(\core.registers[18][9] ),
    .A1(net963),
    .S(net569),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _16501_ (.A0(\core.registers[18][10] ),
    .A1(net968),
    .S(net570),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _16502_ (.A0(\core.registers[18][11] ),
    .A1(net972),
    .S(net569),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _16503_ (.A0(\core.registers[18][12] ),
    .A1(net989),
    .S(net569),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _16504_ (.A0(\core.registers[18][13] ),
    .A1(net986),
    .S(net571),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _16505_ (.A0(\core.registers[18][14] ),
    .A1(net974),
    .S(net570),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _16506_ (.A0(\core.registers[18][15] ),
    .A1(net981),
    .S(net570),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _16507_ (.A0(\core.registers[18][16] ),
    .A1(net1124),
    .S(net568),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _16508_ (.A0(\core.registers[18][17] ),
    .A1(net1130),
    .S(net568),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _16509_ (.A0(\core.registers[18][18] ),
    .A1(net1117),
    .S(net569),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _16510_ (.A0(\core.registers[18][19] ),
    .A1(net1123),
    .S(net568),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _16511_ (.A0(\core.registers[18][20] ),
    .A1(net1138),
    .S(net568),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _16512_ (.A0(\core.registers[18][21] ),
    .A1(net1142),
    .S(net568),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _16513_ (.A0(\core.registers[18][22] ),
    .A1(net1147),
    .S(net569),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _16514_ (.A0(\core.registers[18][23] ),
    .A1(net1151),
    .S(net568),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _16515_ (.A0(\core.registers[18][24] ),
    .A1(net1115),
    .S(net568),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _16516_ (.A0(\core.registers[18][25] ),
    .A1(net1108),
    .S(net568),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _16517_ (.A0(\core.registers[18][26] ),
    .A1(net1102),
    .S(net569),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _16518_ (.A0(\core.registers[18][27] ),
    .A1(net1106),
    .S(net568),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _16519_ (.A0(\core.registers[18][28] ),
    .A1(net1096),
    .S(net568),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _16520_ (.A0(\core.registers[18][29] ),
    .A1(net1092),
    .S(net570),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _16521_ (.A0(\core.registers[18][30] ),
    .A1(net1085),
    .S(net571),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _16522_ (.A0(\core.registers[18][31] ),
    .A1(net1089),
    .S(net570),
    .X(_00745_));
 sky130_fd_sc_hd__nand2_1 _16523_ (.A(\coreWBInterface.state[1] ),
    .B(\coreWBInterface.state[0] ),
    .Y(_03045_));
 sky130_fd_sc_hd__a21oi_1 _16524_ (.A1(_08101_),
    .A2(_03045_),
    .B1(\coreWBInterface.stb ),
    .Y(_03046_));
 sky130_fd_sc_hd__a21o_1 _16525_ (.A1(net42),
    .A2(_07505_),
    .B1(net1968),
    .X(_03047_));
 sky130_fd_sc_hd__a211oi_1 _16526_ (.A1(_07505_),
    .A2(_03045_),
    .B1(_03046_),
    .C1(net1358),
    .Y(_00746_));
 sky130_fd_sc_hd__nand2_1 _16527_ (.A(net9),
    .B(_08101_),
    .Y(_03048_));
 sky130_fd_sc_hd__a21oi_4 _16528_ (.A1(\coreWBInterface.state[1] ),
    .A2(_03048_),
    .B1(\coreWBInterface.state[0] ),
    .Y(_03049_));
 sky130_fd_sc_hd__nand4b_4 _16529_ (.A_N(\coreWBInterface.state[0] ),
    .B(net9),
    .C(_08101_),
    .D(\coreWBInterface.state[1] ),
    .Y(_03050_));
 sky130_fd_sc_hd__o22a_1 _16530_ (.A1(\coreWBInterface.readDataBuffered[0] ),
    .A2(net705),
    .B1(net716),
    .B2(net10),
    .X(_03051_));
 sky130_fd_sc_hd__or2_1 _16531_ (.A(net1356),
    .B(_03051_),
    .X(_00747_));
 sky130_fd_sc_hd__o22a_1 _16532_ (.A1(\coreWBInterface.readDataBuffered[1] ),
    .A2(net706),
    .B1(net717),
    .B2(net21),
    .X(_03052_));
 sky130_fd_sc_hd__or2_1 _16533_ (.A(net1357),
    .B(_03052_),
    .X(_00748_));
 sky130_fd_sc_hd__o22a_1 _16534_ (.A1(\coreWBInterface.readDataBuffered[2] ),
    .A2(net705),
    .B1(net716),
    .B2(net32),
    .X(_03053_));
 sky130_fd_sc_hd__or2_1 _16535_ (.A(net1356),
    .B(_03053_),
    .X(_00749_));
 sky130_fd_sc_hd__o22a_1 _16536_ (.A1(\coreWBInterface.readDataBuffered[3] ),
    .A2(net705),
    .B1(net716),
    .B2(net35),
    .X(_03054_));
 sky130_fd_sc_hd__or2_1 _16537_ (.A(net1356),
    .B(_03054_),
    .X(_00750_));
 sky130_fd_sc_hd__o22a_1 _16538_ (.A1(\coreWBInterface.readDataBuffered[4] ),
    .A2(net703),
    .B1(net714),
    .B2(net36),
    .X(_03055_));
 sky130_fd_sc_hd__or2_1 _16539_ (.A(net1355),
    .B(_03055_),
    .X(_00751_));
 sky130_fd_sc_hd__o22a_1 _16540_ (.A1(\coreWBInterface.readDataBuffered[5] ),
    .A2(net705),
    .B1(net716),
    .B2(net37),
    .X(_03056_));
 sky130_fd_sc_hd__or2_1 _16541_ (.A(net1357),
    .B(_03056_),
    .X(_00752_));
 sky130_fd_sc_hd__o22a_1 _16542_ (.A1(\coreWBInterface.readDataBuffered[6] ),
    .A2(net704),
    .B1(net715),
    .B2(net38),
    .X(_03057_));
 sky130_fd_sc_hd__or2_1 _16543_ (.A(net1356),
    .B(_03057_),
    .X(_00753_));
 sky130_fd_sc_hd__o22a_1 _16544_ (.A1(\coreWBInterface.readDataBuffered[7] ),
    .A2(net705),
    .B1(net716),
    .B2(net39),
    .X(_03058_));
 sky130_fd_sc_hd__or2_1 _16545_ (.A(net1356),
    .B(_03058_),
    .X(_00754_));
 sky130_fd_sc_hd__o22a_1 _16546_ (.A1(\coreWBInterface.readDataBuffered[8] ),
    .A2(net706),
    .B1(net717),
    .B2(net40),
    .X(_03059_));
 sky130_fd_sc_hd__or2_1 _16547_ (.A(net1357),
    .B(_03059_),
    .X(_00755_));
 sky130_fd_sc_hd__o22a_1 _16548_ (.A1(\coreWBInterface.readDataBuffered[9] ),
    .A2(net706),
    .B1(net717),
    .B2(net41),
    .X(_03060_));
 sky130_fd_sc_hd__or2_1 _16549_ (.A(net1358),
    .B(_03060_),
    .X(_00756_));
 sky130_fd_sc_hd__o22a_1 _16550_ (.A1(\coreWBInterface.readDataBuffered[10] ),
    .A2(net705),
    .B1(net716),
    .B2(net11),
    .X(_03061_));
 sky130_fd_sc_hd__or2_1 _16551_ (.A(net1357),
    .B(_03061_),
    .X(_00757_));
 sky130_fd_sc_hd__o22a_1 _16552_ (.A1(\coreWBInterface.readDataBuffered[11] ),
    .A2(net704),
    .B1(net715),
    .B2(net12),
    .X(_03062_));
 sky130_fd_sc_hd__or2_1 _16553_ (.A(net1355),
    .B(_03062_),
    .X(_00758_));
 sky130_fd_sc_hd__o22a_1 _16554_ (.A1(\coreWBInterface.readDataBuffered[12] ),
    .A2(net705),
    .B1(net716),
    .B2(net13),
    .X(_03063_));
 sky130_fd_sc_hd__or2_1 _16555_ (.A(net1356),
    .B(_03063_),
    .X(_00759_));
 sky130_fd_sc_hd__o22a_1 _16556_ (.A1(\coreWBInterface.readDataBuffered[13] ),
    .A2(net704),
    .B1(net715),
    .B2(net14),
    .X(_03064_));
 sky130_fd_sc_hd__or2_1 _16557_ (.A(net1356),
    .B(_03064_),
    .X(_00760_));
 sky130_fd_sc_hd__o22a_1 _16558_ (.A1(\coreWBInterface.readDataBuffered[14] ),
    .A2(net704),
    .B1(net715),
    .B2(net15),
    .X(_03065_));
 sky130_fd_sc_hd__or2_1 _16559_ (.A(net1355),
    .B(_03065_),
    .X(_00761_));
 sky130_fd_sc_hd__o22a_1 _16560_ (.A1(\coreWBInterface.readDataBuffered[15] ),
    .A2(net704),
    .B1(net715),
    .B2(net16),
    .X(_03066_));
 sky130_fd_sc_hd__or2_1 _16561_ (.A(net1355),
    .B(_03066_),
    .X(_00762_));
 sky130_fd_sc_hd__o22a_1 _16562_ (.A1(\coreWBInterface.readDataBuffered[16] ),
    .A2(net703),
    .B1(net714),
    .B2(net17),
    .X(_03067_));
 sky130_fd_sc_hd__or2_1 _16563_ (.A(net1354),
    .B(_03067_),
    .X(_00763_));
 sky130_fd_sc_hd__o22a_1 _16564_ (.A1(\coreWBInterface.readDataBuffered[17] ),
    .A2(net704),
    .B1(net715),
    .B2(net18),
    .X(_03068_));
 sky130_fd_sc_hd__or2_1 _16565_ (.A(net1355),
    .B(_03068_),
    .X(_00764_));
 sky130_fd_sc_hd__o22a_1 _16566_ (.A1(\coreWBInterface.readDataBuffered[18] ),
    .A2(net706),
    .B1(net717),
    .B2(net19),
    .X(_03069_));
 sky130_fd_sc_hd__or2_1 _16567_ (.A(net1358),
    .B(_03069_),
    .X(_00765_));
 sky130_fd_sc_hd__o22a_1 _16568_ (.A1(\coreWBInterface.readDataBuffered[19] ),
    .A2(net704),
    .B1(net715),
    .B2(net20),
    .X(_03070_));
 sky130_fd_sc_hd__or2_1 _16569_ (.A(net1355),
    .B(_03070_),
    .X(_00766_));
 sky130_fd_sc_hd__o22a_1 _16570_ (.A1(\coreWBInterface.readDataBuffered[20] ),
    .A2(net703),
    .B1(net714),
    .B2(net22),
    .X(_03071_));
 sky130_fd_sc_hd__or2_1 _16571_ (.A(net1355),
    .B(_03071_),
    .X(_00767_));
 sky130_fd_sc_hd__o22a_1 _16572_ (.A1(\coreWBInterface.readDataBuffered[21] ),
    .A2(net704),
    .B1(net715),
    .B2(net23),
    .X(_03072_));
 sky130_fd_sc_hd__or2_1 _16573_ (.A(net1354),
    .B(_03072_),
    .X(_00768_));
 sky130_fd_sc_hd__o22a_1 _16574_ (.A1(\coreWBInterface.readDataBuffered[22] ),
    .A2(net705),
    .B1(net716),
    .B2(net24),
    .X(_03073_));
 sky130_fd_sc_hd__or2_1 _16575_ (.A(net1355),
    .B(_03073_),
    .X(_00769_));
 sky130_fd_sc_hd__o22a_1 _16576_ (.A1(\coreWBInterface.readDataBuffered[23] ),
    .A2(net704),
    .B1(net715),
    .B2(net25),
    .X(_03074_));
 sky130_fd_sc_hd__or2_1 _16577_ (.A(net1354),
    .B(_03074_),
    .X(_00770_));
 sky130_fd_sc_hd__o22a_1 _16578_ (.A1(\coreWBInterface.readDataBuffered[24] ),
    .A2(net705),
    .B1(net716),
    .B2(net26),
    .X(_03075_));
 sky130_fd_sc_hd__or2_1 _16579_ (.A(net1354),
    .B(_03075_),
    .X(_00771_));
 sky130_fd_sc_hd__o22a_1 _16580_ (.A1(\coreWBInterface.readDataBuffered[25] ),
    .A2(net703),
    .B1(net714),
    .B2(net27),
    .X(_03076_));
 sky130_fd_sc_hd__or2_1 _16581_ (.A(net1354),
    .B(_03076_),
    .X(_00772_));
 sky130_fd_sc_hd__o22a_1 _16582_ (.A1(\coreWBInterface.readDataBuffered[26] ),
    .A2(net703),
    .B1(net714),
    .B2(net28),
    .X(_03077_));
 sky130_fd_sc_hd__or2_1 _16583_ (.A(net1354),
    .B(_03077_),
    .X(_00773_));
 sky130_fd_sc_hd__o22a_1 _16584_ (.A1(\coreWBInterface.readDataBuffered[27] ),
    .A2(net703),
    .B1(net714),
    .B2(net29),
    .X(_03078_));
 sky130_fd_sc_hd__or2_1 _16585_ (.A(net1354),
    .B(_03078_),
    .X(_00774_));
 sky130_fd_sc_hd__o22a_1 _16586_ (.A1(\coreWBInterface.readDataBuffered[28] ),
    .A2(net703),
    .B1(net714),
    .B2(net30),
    .X(_03079_));
 sky130_fd_sc_hd__or2_1 _16587_ (.A(net1354),
    .B(_03079_),
    .X(_00775_));
 sky130_fd_sc_hd__o22a_1 _16588_ (.A1(\coreWBInterface.readDataBuffered[29] ),
    .A2(net703),
    .B1(net714),
    .B2(net31),
    .X(_03080_));
 sky130_fd_sc_hd__or2_1 _16589_ (.A(net1354),
    .B(_03080_),
    .X(_00776_));
 sky130_fd_sc_hd__o22a_1 _16590_ (.A1(\coreWBInterface.readDataBuffered[30] ),
    .A2(net703),
    .B1(net714),
    .B2(net33),
    .X(_03081_));
 sky130_fd_sc_hd__or2_1 _16591_ (.A(net1354),
    .B(_03081_),
    .X(_00777_));
 sky130_fd_sc_hd__o22a_1 _16592_ (.A1(\coreWBInterface.readDataBuffered[31] ),
    .A2(net703),
    .B1(net714),
    .B2(net34),
    .X(_03082_));
 sky130_fd_sc_hd__or2_1 _16593_ (.A(net1355),
    .B(_03082_),
    .X(_00778_));
 sky130_fd_sc_hd__and3_1 _16594_ (.A(_07505_),
    .B(_08101_),
    .C(_03045_),
    .X(_03083_));
 sky130_fd_sc_hd__inv_2 _16595_ (.A(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__o21a_1 _16596_ (.A1(_07505_),
    .A2(_08101_),
    .B1(_03084_),
    .X(_03085_));
 sky130_fd_sc_hd__o22a_1 _16597_ (.A1(_07505_),
    .A2(_08101_),
    .B1(_03084_),
    .B2(net9),
    .X(_03086_));
 sky130_fd_sc_hd__or3_2 _16598_ (.A(_07505_),
    .B(_08351_),
    .C(_08381_),
    .X(_03087_));
 sky130_fd_sc_hd__a21oi_1 _16599_ (.A1(_03085_),
    .A2(_03087_),
    .B1(net1358),
    .Y(_03088_));
 sky130_fd_sc_hd__o21a_1 _16600_ (.A1(\coreWBInterface.state[0] ),
    .A2(_03086_),
    .B1(_03088_),
    .X(_00779_));
 sky130_fd_sc_hd__a21o_1 _16601_ (.A1(_08352_),
    .A2(net718),
    .B1(_07505_),
    .X(_03089_));
 sky130_fd_sc_hd__a21oi_1 _16602_ (.A1(_03085_),
    .A2(_03089_),
    .B1(net1358),
    .Y(_03090_));
 sky130_fd_sc_hd__o21a_1 _16603_ (.A1(\coreWBInterface.state[1] ),
    .A2(_03086_),
    .B1(_03090_),
    .X(_00780_));
 sky130_fd_sc_hd__nor2_1 _16604_ (.A(_04512_),
    .B(_09105_),
    .Y(_03091_));
 sky130_fd_sc_hd__and3_4 _16605_ (.A(net680),
    .B(net1075),
    .C(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__mux2_1 _16606_ (.A0(\core.registers[24][0] ),
    .A1(net1036),
    .S(net567),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _16607_ (.A0(\core.registers[24][1] ),
    .A1(net1041),
    .S(net566),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _16608_ (.A0(\core.registers[24][2] ),
    .A1(net1046),
    .S(net566),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _16609_ (.A0(\core.registers[24][3] ),
    .A1(net1051),
    .S(net567),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _16610_ (.A0(\core.registers[24][4] ),
    .A1(net1055),
    .S(net567),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _16611_ (.A0(\core.registers[24][5] ),
    .A1(net1058),
    .S(net567),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _16612_ (.A0(\core.registers[24][6] ),
    .A1(net1061),
    .S(net566),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _16613_ (.A0(\core.registers[24][7] ),
    .A1(net1132),
    .S(net566),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _16614_ (.A0(\core.registers[24][8] ),
    .A1(net957),
    .S(net566),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _16615_ (.A0(\core.registers[24][9] ),
    .A1(net962),
    .S(net565),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _16616_ (.A0(\core.registers[24][10] ),
    .A1(net966),
    .S(net567),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _16617_ (.A0(\core.registers[24][11] ),
    .A1(net971),
    .S(net567),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _16618_ (.A0(\core.registers[24][12] ),
    .A1(net987),
    .S(net565),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _16619_ (.A0(\core.registers[24][13] ),
    .A1(net984),
    .S(net566),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _16620_ (.A0(\core.registers[24][14] ),
    .A1(net976),
    .S(net567),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _16621_ (.A0(\core.registers[24][15] ),
    .A1(net979),
    .S(net566),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _16622_ (.A0(\core.registers[24][16] ),
    .A1(net1127),
    .S(net564),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _16623_ (.A0(\core.registers[24][17] ),
    .A1(net1131),
    .S(net564),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _16624_ (.A0(\core.registers[24][18] ),
    .A1(net1117),
    .S(net565),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _16625_ (.A0(\core.registers[24][19] ),
    .A1(net1121),
    .S(net564),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _16626_ (.A0(\core.registers[24][20] ),
    .A1(net1137),
    .S(net564),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _16627_ (.A0(\core.registers[24][21] ),
    .A1(net1140),
    .S(net564),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _16628_ (.A0(\core.registers[24][22] ),
    .A1(net1145),
    .S(net565),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _16629_ (.A0(\core.registers[24][23] ),
    .A1(net1149),
    .S(net564),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _16630_ (.A0(\core.registers[24][24] ),
    .A1(net1112),
    .S(net564),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _16631_ (.A0(\core.registers[24][25] ),
    .A1(net1108),
    .S(net564),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _16632_ (.A0(\core.registers[24][26] ),
    .A1(net1100),
    .S(net565),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _16633_ (.A0(\core.registers[24][27] ),
    .A1(net1104),
    .S(net564),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _16634_ (.A0(\core.registers[24][28] ),
    .A1(net1098),
    .S(net564),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _16635_ (.A0(\core.registers[24][29] ),
    .A1(net1094),
    .S(net566),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _16636_ (.A0(\core.registers[24][30] ),
    .A1(net1084),
    .S(net566),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _16637_ (.A0(\core.registers[24][31] ),
    .A1(net1089),
    .S(net566),
    .X(_00812_));
 sky130_fd_sc_hd__nor2_1 _16638_ (.A(_09086_),
    .B(_09093_),
    .Y(_03093_));
 sky130_fd_sc_hd__and3_4 _16639_ (.A(net676),
    .B(net1072),
    .C(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__mux2_1 _16640_ (.A0(\core.registers[23][0] ),
    .A1(net1037),
    .S(net562),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _16641_ (.A0(\core.registers[23][1] ),
    .A1(net1040),
    .S(net562),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _16642_ (.A0(\core.registers[23][2] ),
    .A1(net1044),
    .S(net563),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _16643_ (.A0(\core.registers[23][3] ),
    .A1(net1048),
    .S(net562),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _16644_ (.A0(\core.registers[23][4] ),
    .A1(net1054),
    .S(net562),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _16645_ (.A0(\core.registers[23][5] ),
    .A1(net1060),
    .S(net563),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _16646_ (.A0(\core.registers[23][6] ),
    .A1(net1062),
    .S(net563),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _16647_ (.A0(\core.registers[23][7] ),
    .A1(net1132),
    .S(net563),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _16648_ (.A0(\core.registers[23][8] ),
    .A1(net960),
    .S(net563),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _16649_ (.A0(\core.registers[23][9] ),
    .A1(net963),
    .S(net561),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _16650_ (.A0(\core.registers[23][10] ),
    .A1(net968),
    .S(net562),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _16651_ (.A0(\core.registers[23][11] ),
    .A1(net972),
    .S(net561),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _16652_ (.A0(\core.registers[23][12] ),
    .A1(net989),
    .S(net561),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _16653_ (.A0(\core.registers[23][13] ),
    .A1(net986),
    .S(net562),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _16654_ (.A0(\core.registers[23][14] ),
    .A1(net974),
    .S(net562),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _16655_ (.A0(\core.registers[23][15] ),
    .A1(net981),
    .S(net562),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _16656_ (.A0(\core.registers[23][16] ),
    .A1(net1125),
    .S(net560),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _16657_ (.A0(\core.registers[23][17] ),
    .A1(net1129),
    .S(net560),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _16658_ (.A0(\core.registers[23][18] ),
    .A1(net1118),
    .S(net561),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _16659_ (.A0(\core.registers[23][19] ),
    .A1(net1122),
    .S(net560),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _16660_ (.A0(\core.registers[23][20] ),
    .A1(net1138),
    .S(net560),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _16661_ (.A0(\core.registers[23][21] ),
    .A1(net1142),
    .S(net560),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _16662_ (.A0(\core.registers[23][22] ),
    .A1(net1147),
    .S(net561),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _16663_ (.A0(\core.registers[23][23] ),
    .A1(net1151),
    .S(net560),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _16664_ (.A0(\core.registers[23][24] ),
    .A1(net1114),
    .S(net560),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _16665_ (.A0(\core.registers[23][25] ),
    .A1(net1108),
    .S(net560),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _16666_ (.A0(\core.registers[23][26] ),
    .A1(net1102),
    .S(net561),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _16667_ (.A0(\core.registers[23][27] ),
    .A1(net1106),
    .S(net560),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _16668_ (.A0(\core.registers[23][28] ),
    .A1(net1098),
    .S(net560),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _16669_ (.A0(\core.registers[23][29] ),
    .A1(net1092),
    .S(net562),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _16670_ (.A0(\core.registers[23][30] ),
    .A1(net1085),
    .S(net563),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _16671_ (.A0(\core.registers[23][31] ),
    .A1(net1089),
    .S(net562),
    .X(_00844_));
 sky130_fd_sc_hd__nor2_1 _16672_ (.A(_09094_),
    .B(_03040_),
    .Y(_03095_));
 sky130_fd_sc_hd__and3_4 _16673_ (.A(net679),
    .B(net1075),
    .C(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__mux2_1 _16674_ (.A0(\core.registers[17][0] ),
    .A1(net1037),
    .S(net558),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _16675_ (.A0(\core.registers[17][1] ),
    .A1(net1040),
    .S(net558),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _16676_ (.A0(\core.registers[17][2] ),
    .A1(net1044),
    .S(net559),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _16677_ (.A0(\core.registers[17][3] ),
    .A1(net1048),
    .S(net558),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _16678_ (.A0(\core.registers[17][4] ),
    .A1(net1054),
    .S(net558),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _16679_ (.A0(\core.registers[17][5] ),
    .A1(net1057),
    .S(net559),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _16680_ (.A0(\core.registers[17][6] ),
    .A1(net1062),
    .S(net559),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _16681_ (.A0(\core.registers[17][7] ),
    .A1(net1133),
    .S(net559),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _16682_ (.A0(\core.registers[17][8] ),
    .A1(net959),
    .S(net559),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _16683_ (.A0(\core.registers[17][9] ),
    .A1(net964),
    .S(net557),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _16684_ (.A0(\core.registers[17][10] ),
    .A1(net969),
    .S(net558),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _16685_ (.A0(\core.registers[17][11] ),
    .A1(net972),
    .S(net557),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _16686_ (.A0(\core.registers[17][12] ),
    .A1(net989),
    .S(net558),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _16687_ (.A0(\core.registers[17][13] ),
    .A1(net986),
    .S(net559),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _16688_ (.A0(\core.registers[17][14] ),
    .A1(net975),
    .S(net558),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _16689_ (.A0(\core.registers[17][15] ),
    .A1(net981),
    .S(net558),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _16690_ (.A0(\core.registers[17][16] ),
    .A1(net1124),
    .S(net556),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _16691_ (.A0(\core.registers[17][17] ),
    .A1(net1128),
    .S(net556),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _16692_ (.A0(\core.registers[17][18] ),
    .A1(net1116),
    .S(net556),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _16693_ (.A0(\core.registers[17][19] ),
    .A1(net1121),
    .S(net556),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _16694_ (.A0(\core.registers[17][20] ),
    .A1(net1138),
    .S(net556),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _16695_ (.A0(\core.registers[17][21] ),
    .A1(net1142),
    .S(net556),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _16696_ (.A0(\core.registers[17][22] ),
    .A1(net1147),
    .S(net557),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _16697_ (.A0(\core.registers[17][23] ),
    .A1(net1151),
    .S(net556),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _16698_ (.A0(\core.registers[17][24] ),
    .A1(net1115),
    .S(net556),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _16699_ (.A0(\core.registers[17][25] ),
    .A1(net1108),
    .S(net556),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _16700_ (.A0(\core.registers[17][26] ),
    .A1(net1102),
    .S(net557),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _16701_ (.A0(\core.registers[17][27] ),
    .A1(net1106),
    .S(net557),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _16702_ (.A0(\core.registers[17][28] ),
    .A1(net1096),
    .S(net556),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _16703_ (.A0(\core.registers[17][29] ),
    .A1(net1092),
    .S(net558),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _16704_ (.A0(\core.registers[17][30] ),
    .A1(net1085),
    .S(net559),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _16705_ (.A0(\core.registers[17][31] ),
    .A1(net1089),
    .S(net558),
    .X(_00876_));
 sky130_fd_sc_hd__a221o_4 _16706_ (.A1(_07836_),
    .A2(_07841_),
    .B1(net713),
    .B2(net1254),
    .C1(_08377_),
    .X(_03097_));
 sky130_fd_sc_hd__o21ba_4 _16707_ (.A1(\wbSRAMInterface.state[0] ),
    .A2(_03097_),
    .B1_N(_07839_),
    .X(_03098_));
 sky130_fd_sc_hd__nand2_1 _16708_ (.A(net1034),
    .B(_09349_),
    .Y(_03099_));
 sky130_fd_sc_hd__or3_4 _16709_ (.A(_07858_),
    .B(_07871_),
    .C(_09240_),
    .X(_03100_));
 sky130_fd_sc_hd__or2_1 _16710_ (.A(_07871_),
    .B(_08771_),
    .X(_03101_));
 sky130_fd_sc_hd__nor2_1 _16711_ (.A(_07844_),
    .B(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__and2_4 _16712_ (.A(\wbSRAMInterface.currentByteSelect[0] ),
    .B(net1255),
    .X(_03103_));
 sky130_fd_sc_hd__and2_2 _16713_ (.A(_07863_),
    .B(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__or4_2 _16714_ (.A(_07858_),
    .B(_07859_),
    .C(_07862_),
    .D(_03101_),
    .X(_03105_));
 sky130_fd_sc_hd__inv_2 _16715_ (.A(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand2_1 _16716_ (.A(net1256),
    .B(_07866_),
    .Y(_03107_));
 sky130_fd_sc_hd__a21o_2 _16717_ (.A1(_07835_),
    .A2(_03107_),
    .B1(_03105_),
    .X(_03108_));
 sky130_fd_sc_hd__a21bo_4 _16718_ (.A1(_07864_),
    .A2(_03108_),
    .B1_N(_07841_),
    .X(_03109_));
 sky130_fd_sc_hd__or4b_4 _16719_ (.A(_07858_),
    .B(_07869_),
    .C(_09240_),
    .D_N(_07870_),
    .X(_03110_));
 sky130_fd_sc_hd__or4_2 _16720_ (.A(_07845_),
    .B(_07855_),
    .C(_07857_),
    .D(_09240_),
    .X(_03111_));
 sky130_fd_sc_hd__a21o_1 _16721_ (.A1(\core.registers[0][0] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03112_));
 sky130_fd_sc_hd__o221a_1 _16722_ (.A1(\core.fetchProgramCounter[0] ),
    .A2(net997),
    .B1(net993),
    .B2(\core.csr.currentInstruction[0] ),
    .C1(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__a21o_1 _16723_ (.A1(net1791),
    .A2(_03103_),
    .B1(_03108_),
    .X(_03114_));
 sky130_fd_sc_hd__a31o_1 _16724_ (.A1(_03099_),
    .A2(_03103_),
    .A3(_03113_),
    .B1(_07864_),
    .X(_03115_));
 sky130_fd_sc_hd__a21bo_1 _16725_ (.A1(_03114_),
    .A2(_03115_),
    .B1_N(_07841_),
    .X(_03116_));
 sky130_fd_sc_hd__and2_4 _16726_ (.A(\localMemoryInterface.wbReadReady ),
    .B(\localMemoryInterface.lastWBByteSelect[0] ),
    .X(_03117_));
 sky130_fd_sc_hd__nand2_1 _16727_ (.A(net68),
    .B(net1799),
    .Y(_03118_));
 sky130_fd_sc_hd__o211a_4 _16728_ (.A1(_04432_),
    .A2(net1799),
    .B1(_03117_),
    .C1(_03118_),
    .X(_03119_));
 sky130_fd_sc_hd__o2bb2a_2 _16729_ (.A1_N(net1305),
    .A2_N(_03116_),
    .B1(_03119_),
    .B2(net2004),
    .X(_03120_));
 sky130_fd_sc_hd__nor2_1 _16730_ (.A(net634),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__a211o_1 _16731_ (.A1(net410),
    .A2(net634),
    .B1(_03121_),
    .C1(net1982),
    .X(_00877_));
 sky130_fd_sc_hd__nand2_1 _16732_ (.A(net1033),
    .B(_09432_),
    .Y(_03122_));
 sky130_fd_sc_hd__a21o_1 _16733_ (.A1(\core.registers[0][1] ),
    .A2(net1027),
    .B1(net1023),
    .X(_03123_));
 sky130_fd_sc_hd__o221a_1 _16734_ (.A1(\core.fetchProgramCounter[1] ),
    .A2(net998),
    .B1(net994),
    .B2(\core.csr.currentInstruction[1] ),
    .C1(_03123_),
    .X(_03124_));
 sky130_fd_sc_hd__a21o_1 _16735_ (.A1(\coreManagement.control[1] ),
    .A2(_03103_),
    .B1(_03108_),
    .X(_03125_));
 sky130_fd_sc_hd__a31o_1 _16736_ (.A1(_03103_),
    .A2(_03122_),
    .A3(_03124_),
    .B1(_07864_),
    .X(_03126_));
 sky130_fd_sc_hd__a21bo_1 _16737_ (.A1(_03125_),
    .A2(_03126_),
    .B1_N(_07841_),
    .X(_03127_));
 sky130_fd_sc_hd__nand2_1 _16738_ (.A(net1799),
    .B(net69),
    .Y(_03128_));
 sky130_fd_sc_hd__o211a_4 _16739_ (.A1(net1799),
    .A2(_04433_),
    .B1(_03117_),
    .C1(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__o2bb2a_2 _16740_ (.A1_N(net1303),
    .A2_N(_03127_),
    .B1(_03129_),
    .B2(net2004),
    .X(_03130_));
 sky130_fd_sc_hd__nor2_1 _16741_ (.A(net634),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__a211o_1 _16742_ (.A1(net421),
    .A2(net634),
    .B1(_03131_),
    .C1(net1982),
    .X(_00878_));
 sky130_fd_sc_hd__nand2_1 _16743_ (.A(net1033),
    .B(_01969_),
    .Y(_03132_));
 sky130_fd_sc_hd__a21o_1 _16744_ (.A1(\core.registers[0][2] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03133_));
 sky130_fd_sc_hd__o221a_1 _16745_ (.A1(\core.fetchProgramCounter[2] ),
    .A2(net997),
    .B1(net993),
    .B2(\core.csr.currentInstruction[2] ),
    .C1(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__a21o_1 _16746_ (.A1(\core.management_interruptEnable ),
    .A2(_03103_),
    .B1(_03108_),
    .X(_03135_));
 sky130_fd_sc_hd__a31o_1 _16747_ (.A1(_03103_),
    .A2(_03132_),
    .A3(_03134_),
    .B1(_07864_),
    .X(_03136_));
 sky130_fd_sc_hd__a21bo_1 _16748_ (.A1(_03135_),
    .A2(_03136_),
    .B1_N(_07841_),
    .X(_03137_));
 sky130_fd_sc_hd__nand2_1 _16749_ (.A(net1799),
    .B(net70),
    .Y(_03138_));
 sky130_fd_sc_hd__o211a_4 _16750_ (.A1(net1799),
    .A2(_04434_),
    .B1(_03117_),
    .C1(_03138_),
    .X(_03139_));
 sky130_fd_sc_hd__o2bb2a_2 _16751_ (.A1_N(net1303),
    .A2_N(_03137_),
    .B1(_03139_),
    .B2(net2005),
    .X(_03140_));
 sky130_fd_sc_hd__nor2_1 _16752_ (.A(net634),
    .B(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__a211o_1 _16753_ (.A1(net432),
    .A2(net634),
    .B1(_03141_),
    .C1(net1982),
    .X(_00879_));
 sky130_fd_sc_hd__nand2_1 _16754_ (.A(net1033),
    .B(_02024_),
    .Y(_03142_));
 sky130_fd_sc_hd__a21o_1 _16755_ (.A1(\core.registers[0][3] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03143_));
 sky130_fd_sc_hd__o21a_1 _16756_ (.A1(\core.csr.currentInstruction[3] ),
    .A2(net993),
    .B1(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__o2111a_1 _16757_ (.A1(\core.fetchProgramCounter[3] ),
    .A2(net998),
    .B1(_03104_),
    .C1(_03142_),
    .D1(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__o21ai_2 _16758_ (.A1(net898),
    .A2(_03145_),
    .B1(net1304),
    .Y(_03146_));
 sky130_fd_sc_hd__mux2_2 _16759_ (.A0(net76),
    .A1(net71),
    .S(net1799),
    .X(_03147_));
 sky130_fd_sc_hd__clkinv_4 _16760_ (.A(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__a21o_2 _16761_ (.A1(_03117_),
    .A2(_03148_),
    .B1(net2003),
    .X(_03149_));
 sky130_fd_sc_hd__a21oi_4 _16762_ (.A1(_03146_),
    .A2(_03149_),
    .B1(net637),
    .Y(_03150_));
 sky130_fd_sc_hd__a211o_1 _16763_ (.A1(net435),
    .A2(net635),
    .B1(_03150_),
    .C1(net1985),
    .X(_00880_));
 sky130_fd_sc_hd__a21o_1 _16764_ (.A1(\core.registers[0][4] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03151_));
 sky130_fd_sc_hd__o21a_1 _16765_ (.A1(\core.csr.currentInstruction[4] ),
    .A2(net993),
    .B1(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__o211a_1 _16766_ (.A1(\core.fetchProgramCounter[4] ),
    .A2(net997),
    .B1(_03104_),
    .C1(_03152_),
    .X(_03153_));
 sky130_fd_sc_hd__o21a_1 _16767_ (.A1(net1032),
    .A2(_02063_),
    .B1(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__o21ai_2 _16768_ (.A1(net898),
    .A2(_03154_),
    .B1(net1304),
    .Y(_03155_));
 sky130_fd_sc_hd__mux2_2 _16769_ (.A0(net87),
    .A1(net72),
    .S(net1804),
    .X(_03156_));
 sky130_fd_sc_hd__clkinv_4 _16770_ (.A(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__a21o_2 _16771_ (.A1(_03117_),
    .A2(_03157_),
    .B1(net2003),
    .X(_03158_));
 sky130_fd_sc_hd__a21oi_4 _16772_ (.A1(_03155_),
    .A2(_03158_),
    .B1(net637),
    .Y(_03159_));
 sky130_fd_sc_hd__a211o_1 _16773_ (.A1(net436),
    .A2(net635),
    .B1(_03159_),
    .C1(net1985),
    .X(_00881_));
 sky130_fd_sc_hd__nand2_1 _16774_ (.A(net1033),
    .B(_02100_),
    .Y(_03160_));
 sky130_fd_sc_hd__a21o_1 _16775_ (.A1(\core.registers[0][5] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03161_));
 sky130_fd_sc_hd__o21a_1 _16776_ (.A1(\core.csr.currentInstruction[5] ),
    .A2(net993),
    .B1(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__o2111a_1 _16777_ (.A1(\core.fetchProgramCounter[5] ),
    .A2(net997),
    .B1(_03104_),
    .C1(_03160_),
    .D1(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__o21ai_2 _16778_ (.A1(net898),
    .A2(_03163_),
    .B1(net1304),
    .Y(_03164_));
 sky130_fd_sc_hd__mux2_2 _16779_ (.A0(net98),
    .A1(net73),
    .S(net1799),
    .X(_03165_));
 sky130_fd_sc_hd__clkinv_4 _16780_ (.A(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__a21o_2 _16781_ (.A1(_03117_),
    .A2(_03166_),
    .B1(net2003),
    .X(_03167_));
 sky130_fd_sc_hd__a21oi_4 _16782_ (.A1(_03164_),
    .A2(_03167_),
    .B1(net637),
    .Y(_03168_));
 sky130_fd_sc_hd__a211o_1 _16783_ (.A1(net437),
    .A2(net635),
    .B1(_03168_),
    .C1(net1985),
    .X(_00882_));
 sky130_fd_sc_hd__nand2_1 _16784_ (.A(net1033),
    .B(_02139_),
    .Y(_03169_));
 sky130_fd_sc_hd__a21o_1 _16785_ (.A1(\core.registers[0][6] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03170_));
 sky130_fd_sc_hd__o21a_1 _16786_ (.A1(\core.csr.currentInstruction[6] ),
    .A2(net993),
    .B1(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__o2111a_1 _16787_ (.A1(\core.fetchProgramCounter[6] ),
    .A2(net997),
    .B1(_03104_),
    .C1(_03169_),
    .D1(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__o21ai_2 _16788_ (.A1(_03109_),
    .A2(_03172_),
    .B1(net1304),
    .Y(_03173_));
 sky130_fd_sc_hd__mux2_2 _16789_ (.A0(net103),
    .A1(net74),
    .S(net1799),
    .X(_03174_));
 sky130_fd_sc_hd__clkinv_4 _16790_ (.A(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__a21o_2 _16791_ (.A1(_03117_),
    .A2(_03175_),
    .B1(net2003),
    .X(_03176_));
 sky130_fd_sc_hd__a21oi_4 _16792_ (.A1(_03173_),
    .A2(_03176_),
    .B1(net637),
    .Y(_03177_));
 sky130_fd_sc_hd__a211o_1 _16793_ (.A1(net438),
    .A2(net635),
    .B1(_03177_),
    .C1(net1985),
    .X(_00883_));
 sky130_fd_sc_hd__nand2_1 _16794_ (.A(net1033),
    .B(_02162_),
    .Y(_03178_));
 sky130_fd_sc_hd__a21o_1 _16795_ (.A1(\core.registers[0][7] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03179_));
 sky130_fd_sc_hd__o21a_1 _16796_ (.A1(\core.csr.currentInstruction[7] ),
    .A2(net993),
    .B1(_03179_),
    .X(_03180_));
 sky130_fd_sc_hd__o2111a_1 _16797_ (.A1(\core.fetchProgramCounter[7] ),
    .A2(net998),
    .B1(_03104_),
    .C1(_03178_),
    .D1(_03180_),
    .X(_03181_));
 sky130_fd_sc_hd__o21ai_2 _16798_ (.A1(_03109_),
    .A2(_03181_),
    .B1(net1305),
    .Y(_03182_));
 sky130_fd_sc_hd__mux2_2 _16799_ (.A0(net104),
    .A1(net75),
    .S(net1799),
    .X(_03183_));
 sky130_fd_sc_hd__clkinv_4 _16800_ (.A(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__a21o_2 _16801_ (.A1(_03117_),
    .A2(_03184_),
    .B1(net2003),
    .X(_03185_));
 sky130_fd_sc_hd__a21oi_4 _16802_ (.A1(_03182_),
    .A2(_03185_),
    .B1(net637),
    .Y(_03186_));
 sky130_fd_sc_hd__a211o_1 _16803_ (.A1(net439),
    .A2(net636),
    .B1(_03186_),
    .C1(net1986),
    .X(_00884_));
 sky130_fd_sc_hd__nand2_1 _16804_ (.A(net1033),
    .B(_02212_),
    .Y(_03187_));
 sky130_fd_sc_hd__and3_4 _16805_ (.A(\wbSRAMInterface.currentByteSelect[1] ),
    .B(net1255),
    .C(_07863_),
    .X(_03188_));
 sky130_fd_sc_hd__a21o_2 _16806_ (.A1(\core.registers[0][8] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03189_));
 sky130_fd_sc_hd__o221a_1 _16807_ (.A1(\core.fetchProgramCounter[8] ),
    .A2(net997),
    .B1(net994),
    .B2(\core.csr.currentInstruction[8] ),
    .C1(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__a31o_1 _16808_ (.A1(_03187_),
    .A2(_03188_),
    .A3(_03190_),
    .B1(net898),
    .X(_03191_));
 sky130_fd_sc_hd__and2_4 _16809_ (.A(\localMemoryInterface.wbReadReady ),
    .B(\localMemoryInterface.lastWBByteSelect[1] ),
    .X(_03192_));
 sky130_fd_sc_hd__nand2_1 _16810_ (.A(net1800),
    .B(net77),
    .Y(_03193_));
 sky130_fd_sc_hd__o211a_4 _16811_ (.A1(net1800),
    .A2(_04435_),
    .B1(_03192_),
    .C1(_03193_),
    .X(_03194_));
 sky130_fd_sc_hd__o2bb2a_2 _16812_ (.A1_N(net1304),
    .A2_N(_03191_),
    .B1(_03194_),
    .B2(net2006),
    .X(_03195_));
 sky130_fd_sc_hd__nor2_1 _16813_ (.A(net635),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__a211o_1 _16814_ (.A1(net440),
    .A2(net636),
    .B1(_03196_),
    .C1(net1986),
    .X(_00885_));
 sky130_fd_sc_hd__nand2_1 _16815_ (.A(net1034),
    .B(_02240_),
    .Y(_03197_));
 sky130_fd_sc_hd__a21o_1 _16816_ (.A1(\core.registers[0][9] ),
    .A2(net1028),
    .B1(net1024),
    .X(_03198_));
 sky130_fd_sc_hd__o221a_1 _16817_ (.A1(\core.fetchProgramCounter[9] ),
    .A2(net996),
    .B1(net992),
    .B2(\core.csr.currentInstruction[9] ),
    .C1(_03198_),
    .X(_03199_));
 sky130_fd_sc_hd__a31o_1 _16818_ (.A1(_03188_),
    .A2(_03197_),
    .A3(_03199_),
    .B1(net896),
    .X(_03200_));
 sky130_fd_sc_hd__nand2_1 _16819_ (.A(net1800),
    .B(net78),
    .Y(_03201_));
 sky130_fd_sc_hd__o211a_4 _16820_ (.A1(net1800),
    .A2(_04436_),
    .B1(_03192_),
    .C1(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__o2bb2a_2 _16821_ (.A1_N(net1302),
    .A2_N(_03200_),
    .B1(_03202_),
    .B2(net2003),
    .X(_03203_));
 sky130_fd_sc_hd__nor2_1 _16822_ (.A(net634),
    .B(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__a211o_1 _16823_ (.A1(net441),
    .A2(_03098_),
    .B1(_03204_),
    .C1(net1981),
    .X(_00886_));
 sky130_fd_sc_hd__nand2_1 _16824_ (.A(net1034),
    .B(_02269_),
    .Y(_03205_));
 sky130_fd_sc_hd__a21o_1 _16825_ (.A1(\core.registers[0][10] ),
    .A2(net1027),
    .B1(net1023),
    .X(_03206_));
 sky130_fd_sc_hd__o221a_1 _16826_ (.A1(\core.fetchProgramCounter[10] ),
    .A2(net998),
    .B1(net994),
    .B2(\core.csr.currentInstruction[10] ),
    .C1(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__a31o_1 _16827_ (.A1(_03188_),
    .A2(_03205_),
    .A3(_03207_),
    .B1(net896),
    .X(_03208_));
 sky130_fd_sc_hd__nand2_1 _16828_ (.A(net1800),
    .B(net79),
    .Y(_03209_));
 sky130_fd_sc_hd__o211a_4 _16829_ (.A1(net1800),
    .A2(_04437_),
    .B1(_03192_),
    .C1(_03209_),
    .X(_03210_));
 sky130_fd_sc_hd__o2bb2a_4 _16830_ (.A1_N(net1302),
    .A2_N(_03208_),
    .B1(_03210_),
    .B2(net2003),
    .X(_03211_));
 sky130_fd_sc_hd__nor2_1 _16831_ (.A(net635),
    .B(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__a211o_1 _16832_ (.A1(net411),
    .A2(net635),
    .B1(_03212_),
    .C1(net1986),
    .X(_00887_));
 sky130_fd_sc_hd__nand2_1 _16833_ (.A(net1034),
    .B(_02299_),
    .Y(_03213_));
 sky130_fd_sc_hd__a21o_1 _16834_ (.A1(\core.registers[0][11] ),
    .A2(net1027),
    .B1(net1023),
    .X(_03214_));
 sky130_fd_sc_hd__o221a_1 _16835_ (.A1(\core.fetchProgramCounter[11] ),
    .A2(net996),
    .B1(net992),
    .B2(\core.csr.currentInstruction[11] ),
    .C1(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__a31o_1 _16836_ (.A1(_03188_),
    .A2(_03213_),
    .A3(_03215_),
    .B1(net896),
    .X(_03216_));
 sky130_fd_sc_hd__nand2_1 _16837_ (.A(net1800),
    .B(net80),
    .Y(_03217_));
 sky130_fd_sc_hd__o211a_4 _16838_ (.A1(net1800),
    .A2(_04438_),
    .B1(_03192_),
    .C1(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__o2bb2a_4 _16839_ (.A1_N(net1302),
    .A2_N(_03216_),
    .B1(_03218_),
    .B2(net2003),
    .X(_03219_));
 sky130_fd_sc_hd__nor2_1 _16840_ (.A(net639),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__a211o_1 _16841_ (.A1(net412),
    .A2(net639),
    .B1(_03220_),
    .C1(net1986),
    .X(_00888_));
 sky130_fd_sc_hd__nand2_1 _16842_ (.A(net1034),
    .B(_02329_),
    .Y(_03221_));
 sky130_fd_sc_hd__a21o_1 _16843_ (.A1(\core.registers[0][12] ),
    .A2(net1027),
    .B1(net1023),
    .X(_03222_));
 sky130_fd_sc_hd__o221a_1 _16844_ (.A1(\core.fetchProgramCounter[12] ),
    .A2(net998),
    .B1(net992),
    .B2(\core.csr.currentInstruction[12] ),
    .C1(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__a31o_1 _16845_ (.A1(_03188_),
    .A2(_03221_),
    .A3(_03223_),
    .B1(net896),
    .X(_03224_));
 sky130_fd_sc_hd__nand2_1 _16846_ (.A(net1800),
    .B(net81),
    .Y(_03225_));
 sky130_fd_sc_hd__o211a_4 _16847_ (.A1(net1800),
    .A2(_04439_),
    .B1(_03192_),
    .C1(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__o2bb2a_4 _16848_ (.A1_N(net1302),
    .A2_N(_03224_),
    .B1(_03226_),
    .B2(net2003),
    .X(_03227_));
 sky130_fd_sc_hd__nor2_1 _16849_ (.A(net635),
    .B(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__a211o_1 _16850_ (.A1(net413),
    .A2(net635),
    .B1(_03228_),
    .C1(net1986),
    .X(_00889_));
 sky130_fd_sc_hd__nand2_1 _16851_ (.A(net1033),
    .B(_02352_),
    .Y(_03229_));
 sky130_fd_sc_hd__a21o_1 _16852_ (.A1(\core.registers[0][13] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03230_));
 sky130_fd_sc_hd__o221a_1 _16853_ (.A1(\core.fetchProgramCounter[13] ),
    .A2(net997),
    .B1(net993),
    .B2(\core.csr.currentInstruction[13] ),
    .C1(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__a31o_1 _16854_ (.A1(_03188_),
    .A2(_03229_),
    .A3(_03231_),
    .B1(net898),
    .X(_03232_));
 sky130_fd_sc_hd__nand2_1 _16855_ (.A(net1801),
    .B(net82),
    .Y(_03233_));
 sky130_fd_sc_hd__o211a_4 _16856_ (.A1(net1801),
    .A2(_04440_),
    .B1(_03192_),
    .C1(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__o2bb2a_2 _16857_ (.A1_N(net1304),
    .A2_N(_03232_),
    .B1(_03234_),
    .B2(net2006),
    .X(_03235_));
 sky130_fd_sc_hd__nor2_1 _16858_ (.A(net636),
    .B(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__a211o_1 _16859_ (.A1(net414),
    .A2(net636),
    .B1(_03236_),
    .C1(net1986),
    .X(_00890_));
 sky130_fd_sc_hd__nand2_1 _16860_ (.A(net1034),
    .B(_02384_),
    .Y(_03237_));
 sky130_fd_sc_hd__a21o_1 _16861_ (.A1(\core.registers[0][14] ),
    .A2(net1027),
    .B1(net1023),
    .X(_03238_));
 sky130_fd_sc_hd__o221a_1 _16862_ (.A1(\core.fetchProgramCounter[14] ),
    .A2(net998),
    .B1(net994),
    .B2(\core.csr.currentInstruction[14] ),
    .C1(_03238_),
    .X(_03239_));
 sky130_fd_sc_hd__a31o_1 _16863_ (.A1(_03188_),
    .A2(_03237_),
    .A3(_03239_),
    .B1(net897),
    .X(_03240_));
 sky130_fd_sc_hd__nand2_1 _16864_ (.A(net1801),
    .B(net83),
    .Y(_03241_));
 sky130_fd_sc_hd__o211a_4 _16865_ (.A1(net1801),
    .A2(_04441_),
    .B1(_03192_),
    .C1(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__o2bb2a_4 _16866_ (.A1_N(net1303),
    .A2_N(_03240_),
    .B1(_03242_),
    .B2(net2005),
    .X(_03243_));
 sky130_fd_sc_hd__nor2_1 _16867_ (.A(net636),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__a211o_1 _16868_ (.A1(net415),
    .A2(net636),
    .B1(_03244_),
    .C1(net1986),
    .X(_00891_));
 sky130_fd_sc_hd__nand2_1 _16869_ (.A(net1033),
    .B(_02415_),
    .Y(_03245_));
 sky130_fd_sc_hd__a21o_1 _16870_ (.A1(\core.registers[0][15] ),
    .A2(net1026),
    .B1(net1022),
    .X(_03246_));
 sky130_fd_sc_hd__o221a_1 _16871_ (.A1(\core.fetchProgramCounter[15] ),
    .A2(net997),
    .B1(net993),
    .B2(\core.csr.currentInstruction[15] ),
    .C1(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__a31o_1 _16872_ (.A1(_03188_),
    .A2(_03245_),
    .A3(_03247_),
    .B1(net898),
    .X(_03248_));
 sky130_fd_sc_hd__nand2_1 _16873_ (.A(net1801),
    .B(net84),
    .Y(_03249_));
 sky130_fd_sc_hd__o211a_4 _16874_ (.A1(net1801),
    .A2(_04442_),
    .B1(_03192_),
    .C1(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__o2bb2a_4 _16875_ (.A1_N(net1304),
    .A2_N(_03248_),
    .B1(_03250_),
    .B2(net2006),
    .X(_03251_));
 sky130_fd_sc_hd__nor2_1 _16876_ (.A(net639),
    .B(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__a211o_1 _16877_ (.A1(net416),
    .A2(net639),
    .B1(_03252_),
    .C1(net1995),
    .X(_00892_));
 sky130_fd_sc_hd__nand2_1 _16878_ (.A(net1034),
    .B(_02451_),
    .Y(_03253_));
 sky130_fd_sc_hd__and3_4 _16879_ (.A(\wbSRAMInterface.currentByteSelect[2] ),
    .B(net1255),
    .C(_07863_),
    .X(_03254_));
 sky130_fd_sc_hd__a21o_2 _16880_ (.A1(\core.registers[0][16] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03255_));
 sky130_fd_sc_hd__o221a_2 _16881_ (.A1(\core.fetchProgramCounter[16] ),
    .A2(net996),
    .B1(net992),
    .B2(\core.csr.currentInstruction[16] ),
    .C1(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__a31o_1 _16882_ (.A1(_03253_),
    .A2(_03254_),
    .A3(_03256_),
    .B1(net896),
    .X(_03257_));
 sky130_fd_sc_hd__nand2_8 _16883_ (.A(\localMemoryInterface.wbReadReady ),
    .B(\localMemoryInterface.lastWBByteSelect[2] ),
    .Y(_03258_));
 sky130_fd_sc_hd__mux2_8 _16884_ (.A0(net50),
    .A1(net85),
    .S(net1801),
    .X(_03259_));
 sky130_fd_sc_hd__nor2_1 _16885_ (.A(_03258_),
    .B(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__o2bb2a_4 _16886_ (.A1_N(net1302),
    .A2_N(_03257_),
    .B1(_03260_),
    .B2(net2003),
    .X(_03261_));
 sky130_fd_sc_hd__nor2_1 _16887_ (.A(net636),
    .B(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__a211o_1 _16888_ (.A1(net417),
    .A2(net636),
    .B1(_03262_),
    .C1(net1986),
    .X(_00893_));
 sky130_fd_sc_hd__a21o_2 _16889_ (.A1(\core.registers[0][17] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03263_));
 sky130_fd_sc_hd__o221a_1 _16890_ (.A1(\core.fetchProgramCounter[17] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[17] ),
    .C1(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__o211a_2 _16891_ (.A1(net1031),
    .A2(_02478_),
    .B1(_03254_),
    .C1(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__o21ai_2 _16892_ (.A1(net896),
    .A2(_03265_),
    .B1(net1302),
    .Y(_03266_));
 sky130_fd_sc_hd__mux2_8 _16893_ (.A0(net51),
    .A1(net86),
    .S(net1802),
    .X(_03267_));
 sky130_fd_sc_hd__o21bai_4 _16894_ (.A1(_03258_),
    .A2(_03267_),
    .B1_N(net2005),
    .Y(_03268_));
 sky130_fd_sc_hd__a21oi_4 _16895_ (.A1(_03266_),
    .A2(_03268_),
    .B1(net633),
    .Y(_03269_));
 sky130_fd_sc_hd__a211o_1 _16896_ (.A1(net418),
    .A2(net635),
    .B1(_03269_),
    .C1(net1986),
    .X(_00894_));
 sky130_fd_sc_hd__a21o_1 _16897_ (.A1(\core.registers[0][18] ),
    .A2(net1028),
    .B1(net1024),
    .X(_03270_));
 sky130_fd_sc_hd__o221a_1 _16898_ (.A1(\core.fetchProgramCounter[18] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[18] ),
    .C1(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__o211a_2 _16899_ (.A1(net1031),
    .A2(_02504_),
    .B1(_03254_),
    .C1(_03271_),
    .X(_03272_));
 sky130_fd_sc_hd__o21ai_2 _16900_ (.A1(net896),
    .A2(_03272_),
    .B1(net1302),
    .Y(_03273_));
 sky130_fd_sc_hd__mux2_8 _16901_ (.A0(net52),
    .A1(net88),
    .S(net1802),
    .X(_03274_));
 sky130_fd_sc_hd__o21bai_4 _16902_ (.A1(_03258_),
    .A2(_03274_),
    .B1_N(net2005),
    .Y(_03275_));
 sky130_fd_sc_hd__a21oi_4 _16903_ (.A1(_03273_),
    .A2(_03275_),
    .B1(net633),
    .Y(_03276_));
 sky130_fd_sc_hd__a211o_1 _16904_ (.A1(net419),
    .A2(net639),
    .B1(_03276_),
    .C1(net1995),
    .X(_00895_));
 sky130_fd_sc_hd__a21o_1 _16905_ (.A1(\core.registers[0][19] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03277_));
 sky130_fd_sc_hd__o221a_1 _16906_ (.A1(\core.fetchProgramCounter[19] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[19] ),
    .C1(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__o211a_2 _16907_ (.A1(net1031),
    .A2(_02530_),
    .B1(_03254_),
    .C1(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__o21ai_2 _16908_ (.A1(net896),
    .A2(_03279_),
    .B1(net1302),
    .Y(_03280_));
 sky130_fd_sc_hd__mux2_8 _16909_ (.A0(net53),
    .A1(net89),
    .S(net1802),
    .X(_03281_));
 sky130_fd_sc_hd__o21bai_4 _16910_ (.A1(_03258_),
    .A2(_03281_),
    .B1_N(net2004),
    .Y(_03282_));
 sky130_fd_sc_hd__a21oi_4 _16911_ (.A1(_03280_),
    .A2(_03282_),
    .B1(net633),
    .Y(_03283_));
 sky130_fd_sc_hd__a211o_1 _16912_ (.A1(net420),
    .A2(net639),
    .B1(_03283_),
    .C1(net1987),
    .X(_00896_));
 sky130_fd_sc_hd__a21o_2 _16913_ (.A1(\core.registers[0][20] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03284_));
 sky130_fd_sc_hd__o221a_1 _16914_ (.A1(\core.fetchProgramCounter[20] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[20] ),
    .C1(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__o211a_2 _16915_ (.A1(net1031),
    .A2(_02557_),
    .B1(_03254_),
    .C1(_03285_),
    .X(_03286_));
 sky130_fd_sc_hd__o21ai_2 _16916_ (.A1(net896),
    .A2(_03286_),
    .B1(net1302),
    .Y(_03287_));
 sky130_fd_sc_hd__mux2_8 _16917_ (.A0(net55),
    .A1(net90),
    .S(net1802),
    .X(_03288_));
 sky130_fd_sc_hd__o21bai_4 _16918_ (.A1(_03258_),
    .A2(_03288_),
    .B1_N(net2004),
    .Y(_03289_));
 sky130_fd_sc_hd__a21oi_4 _16919_ (.A1(_03287_),
    .A2(_03289_),
    .B1(net633),
    .Y(_03290_));
 sky130_fd_sc_hd__a211o_1 _16920_ (.A1(net422),
    .A2(net639),
    .B1(_03290_),
    .C1(net1996),
    .X(_00897_));
 sky130_fd_sc_hd__a21o_2 _16921_ (.A1(\core.registers[0][21] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03291_));
 sky130_fd_sc_hd__o221a_1 _16922_ (.A1(\core.fetchProgramCounter[21] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[21] ),
    .C1(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__o211a_2 _16923_ (.A1(net1031),
    .A2(_02583_),
    .B1(_03254_),
    .C1(_03292_),
    .X(_03293_));
 sky130_fd_sc_hd__o21ai_2 _16924_ (.A1(net897),
    .A2(_03293_),
    .B1(net1303),
    .Y(_03294_));
 sky130_fd_sc_hd__mux2_8 _16925_ (.A0(net56),
    .A1(net91),
    .S(net1802),
    .X(_03295_));
 sky130_fd_sc_hd__o21bai_4 _16926_ (.A1(_03258_),
    .A2(_03295_),
    .B1_N(net2004),
    .Y(_03296_));
 sky130_fd_sc_hd__a21oi_4 _16927_ (.A1(_03294_),
    .A2(_03296_),
    .B1(net633),
    .Y(_03297_));
 sky130_fd_sc_hd__a211o_1 _16928_ (.A1(net423),
    .A2(net638),
    .B1(_03297_),
    .C1(net1999),
    .X(_00898_));
 sky130_fd_sc_hd__a21o_1 _16929_ (.A1(\core.registers[0][22] ),
    .A2(net1028),
    .B1(net1024),
    .X(_03298_));
 sky130_fd_sc_hd__o221a_2 _16930_ (.A1(\core.fetchProgramCounter[22] ),
    .A2(net996),
    .B1(net992),
    .B2(\core.csr.currentInstruction[22] ),
    .C1(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__o211a_1 _16931_ (.A1(net1032),
    .A2(_02609_),
    .B1(_03254_),
    .C1(_03299_),
    .X(_03300_));
 sky130_fd_sc_hd__o21ai_2 _16932_ (.A1(net896),
    .A2(_03300_),
    .B1(net1302),
    .Y(_03301_));
 sky130_fd_sc_hd__mux2_8 _16933_ (.A0(net57),
    .A1(net92),
    .S(net1802),
    .X(_03302_));
 sky130_fd_sc_hd__o21bai_4 _16934_ (.A1(_03258_),
    .A2(_03302_),
    .B1_N(net2004),
    .Y(_03303_));
 sky130_fd_sc_hd__a21oi_4 _16935_ (.A1(_03301_),
    .A2(_03303_),
    .B1(net634),
    .Y(_03304_));
 sky130_fd_sc_hd__a211o_1 _16936_ (.A1(net424),
    .A2(net638),
    .B1(_03304_),
    .C1(net1999),
    .X(_00899_));
 sky130_fd_sc_hd__a21o_1 _16937_ (.A1(\core.registers[0][23] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03305_));
 sky130_fd_sc_hd__o221a_1 _16938_ (.A1(\core.fetchProgramCounter[23] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[23] ),
    .C1(_03305_),
    .X(_03306_));
 sky130_fd_sc_hd__o211a_2 _16939_ (.A1(net1031),
    .A2(_02635_),
    .B1(_03254_),
    .C1(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__o21ai_2 _16940_ (.A1(net897),
    .A2(_03307_),
    .B1(net1305),
    .Y(_03308_));
 sky130_fd_sc_hd__mux2_8 _16941_ (.A0(net58),
    .A1(net93),
    .S(net1802),
    .X(_03309_));
 sky130_fd_sc_hd__o21bai_4 _16942_ (.A1(_03258_),
    .A2(_03309_),
    .B1_N(net2004),
    .Y(_03310_));
 sky130_fd_sc_hd__a21oi_4 _16943_ (.A1(_03308_),
    .A2(_03310_),
    .B1(net634),
    .Y(_03311_));
 sky130_fd_sc_hd__a211o_1 _16944_ (.A1(net425),
    .A2(net639),
    .B1(_03311_),
    .C1(net2000),
    .X(_00900_));
 sky130_fd_sc_hd__and3_4 _16945_ (.A(\wbSRAMInterface.currentByteSelect[3] ),
    .B(net1255),
    .C(_07863_),
    .X(_03312_));
 sky130_fd_sc_hd__a21o_1 _16946_ (.A1(\core.registers[0][24] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03313_));
 sky130_fd_sc_hd__o221a_1 _16947_ (.A1(\core.fetchProgramCounter[24] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[24] ),
    .C1(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__o211a_2 _16948_ (.A1(net1031),
    .A2(_02661_),
    .B1(_03312_),
    .C1(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__o21ai_2 _16949_ (.A1(net897),
    .A2(_03315_),
    .B1(net1303),
    .Y(_03316_));
 sky130_fd_sc_hd__nand2_8 _16950_ (.A(\localMemoryInterface.wbReadReady ),
    .B(\localMemoryInterface.lastWBByteSelect[3] ),
    .Y(_03317_));
 sky130_fd_sc_hd__mux2_8 _16951_ (.A0(net59),
    .A1(net94),
    .S(net1802),
    .X(_03318_));
 sky130_fd_sc_hd__o21bai_4 _16952_ (.A1(_03317_),
    .A2(_03318_),
    .B1_N(net2004),
    .Y(_03319_));
 sky130_fd_sc_hd__a21oi_4 _16953_ (.A1(_03316_),
    .A2(_03319_),
    .B1(net633),
    .Y(_03320_));
 sky130_fd_sc_hd__a211o_1 _16954_ (.A1(net426),
    .A2(net638),
    .B1(_03320_),
    .C1(net2000),
    .X(_00901_));
 sky130_fd_sc_hd__a21o_1 _16955_ (.A1(\core.registers[0][25] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03321_));
 sky130_fd_sc_hd__o221a_2 _16956_ (.A1(\core.fetchProgramCounter[25] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[25] ),
    .C1(_03321_),
    .X(_03322_));
 sky130_fd_sc_hd__o211a_2 _16957_ (.A1(net1031),
    .A2(_02681_),
    .B1(_03312_),
    .C1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__o21ai_2 _16958_ (.A1(net897),
    .A2(_03323_),
    .B1(net1303),
    .Y(_03324_));
 sky130_fd_sc_hd__mux2_8 _16959_ (.A0(net60),
    .A1(net95),
    .S(net1803),
    .X(_03325_));
 sky130_fd_sc_hd__o21bai_4 _16960_ (.A1(_03317_),
    .A2(_03325_),
    .B1_N(net2004),
    .Y(_03326_));
 sky130_fd_sc_hd__a21oi_4 _16961_ (.A1(_03324_),
    .A2(_03326_),
    .B1(net633),
    .Y(_03327_));
 sky130_fd_sc_hd__a211o_1 _16962_ (.A1(net427),
    .A2(net638),
    .B1(_03327_),
    .C1(net2000),
    .X(_00902_));
 sky130_fd_sc_hd__a21o_1 _16963_ (.A1(\core.registers[0][26] ),
    .A2(net1028),
    .B1(net1024),
    .X(_03328_));
 sky130_fd_sc_hd__o221a_1 _16964_ (.A1(\core.fetchProgramCounter[26] ),
    .A2(net996),
    .B1(net992),
    .B2(\core.csr.currentInstruction[26] ),
    .C1(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__o211a_2 _16965_ (.A1(net1032),
    .A2(_02714_),
    .B1(_03312_),
    .C1(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__o21ai_2 _16966_ (.A1(net897),
    .A2(_03330_),
    .B1(net1303),
    .Y(_03331_));
 sky130_fd_sc_hd__mux2_8 _16967_ (.A0(net61),
    .A1(net96),
    .S(net1802),
    .X(_03332_));
 sky130_fd_sc_hd__o21bai_4 _16968_ (.A1(_03317_),
    .A2(_03332_),
    .B1_N(net2006),
    .Y(_03333_));
 sky130_fd_sc_hd__a21oi_4 _16969_ (.A1(_03331_),
    .A2(_03333_),
    .B1(net633),
    .Y(_03334_));
 sky130_fd_sc_hd__a211o_1 _16970_ (.A1(net428),
    .A2(net638),
    .B1(_03334_),
    .C1(net2000),
    .X(_00903_));
 sky130_fd_sc_hd__a21o_1 _16971_ (.A1(\core.registers[0][27] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03335_));
 sky130_fd_sc_hd__o221a_2 _16972_ (.A1(\core.fetchProgramCounter[27] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[27] ),
    .C1(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__o211a_2 _16973_ (.A1(net1031),
    .A2(_02740_),
    .B1(_03312_),
    .C1(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__o21ai_2 _16974_ (.A1(net897),
    .A2(_03337_),
    .B1(net1303),
    .Y(_03338_));
 sky130_fd_sc_hd__mux2_8 _16975_ (.A0(net62),
    .A1(net97),
    .S(net1802),
    .X(_03339_));
 sky130_fd_sc_hd__o21bai_4 _16976_ (.A1(_03317_),
    .A2(_03339_),
    .B1_N(net2004),
    .Y(_03340_));
 sky130_fd_sc_hd__a21oi_4 _16977_ (.A1(_03338_),
    .A2(_03340_),
    .B1(net633),
    .Y(_03341_));
 sky130_fd_sc_hd__a211o_1 _16978_ (.A1(net429),
    .A2(net638),
    .B1(_03341_),
    .C1(net2000),
    .X(_00904_));
 sky130_fd_sc_hd__a21o_2 _16979_ (.A1(\core.registers[0][28] ),
    .A2(net1025),
    .B1(net1021),
    .X(_03342_));
 sky130_fd_sc_hd__o221a_1 _16980_ (.A1(\core.fetchProgramCounter[28] ),
    .A2(net995),
    .B1(net991),
    .B2(\core.csr.currentInstruction[28] ),
    .C1(_03342_),
    .X(_03343_));
 sky130_fd_sc_hd__o211a_2 _16981_ (.A1(net1031),
    .A2(_02768_),
    .B1(_03312_),
    .C1(_03343_),
    .X(_03344_));
 sky130_fd_sc_hd__o21ai_2 _16982_ (.A1(net898),
    .A2(_03344_),
    .B1(net1303),
    .Y(_03345_));
 sky130_fd_sc_hd__mux2_8 _16983_ (.A0(net63),
    .A1(net99),
    .S(net1803),
    .X(_03346_));
 sky130_fd_sc_hd__o21bai_4 _16984_ (.A1(_03317_),
    .A2(_03346_),
    .B1_N(net2006),
    .Y(_03347_));
 sky130_fd_sc_hd__a21oi_4 _16985_ (.A1(_03345_),
    .A2(_03347_),
    .B1(net633),
    .Y(_03348_));
 sky130_fd_sc_hd__a211o_1 _16986_ (.A1(net430),
    .A2(net638),
    .B1(_03348_),
    .C1(net2001),
    .X(_00905_));
 sky130_fd_sc_hd__o221a_1 _16987_ (.A1(\core.fetchProgramCounter[29] ),
    .A2(net997),
    .B1(net994),
    .B2(\core.csr.currentInstruction[29] ),
    .C1(_03312_),
    .X(_03349_));
 sky130_fd_sc_hd__a21o_1 _16988_ (.A1(\core.registers[0][29] ),
    .A2(net1027),
    .B1(net1023),
    .X(_03350_));
 sky130_fd_sc_hd__o211a_1 _16989_ (.A1(net1032),
    .A2(_02795_),
    .B1(_03349_),
    .C1(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__o21ai_2 _16990_ (.A1(net898),
    .A2(_03351_),
    .B1(net1304),
    .Y(_03352_));
 sky130_fd_sc_hd__mux2_8 _16991_ (.A0(net64),
    .A1(net100),
    .S(net1803),
    .X(_03353_));
 sky130_fd_sc_hd__o21bai_4 _16992_ (.A1(_03317_),
    .A2(_03353_),
    .B1_N(net2006),
    .Y(_03354_));
 sky130_fd_sc_hd__a21oi_4 _16993_ (.A1(_03352_),
    .A2(_03354_),
    .B1(net637),
    .Y(_03355_));
 sky130_fd_sc_hd__a211o_1 _16994_ (.A1(net431),
    .A2(net638),
    .B1(_03355_),
    .C1(net2001),
    .X(_00906_));
 sky130_fd_sc_hd__a21o_1 _16995_ (.A1(\core.registers[0][30] ),
    .A2(net1027),
    .B1(net1023),
    .X(_03356_));
 sky130_fd_sc_hd__o221a_1 _16996_ (.A1(\core.fetchProgramCounter[30] ),
    .A2(net997),
    .B1(net993),
    .B2(\core.csr.currentInstruction[30] ),
    .C1(_03356_),
    .X(_03357_));
 sky130_fd_sc_hd__o211a_1 _16997_ (.A1(net1032),
    .A2(_02815_),
    .B1(_03312_),
    .C1(_03357_),
    .X(_03358_));
 sky130_fd_sc_hd__o21ai_2 _16998_ (.A1(net898),
    .A2(_03358_),
    .B1(net1304),
    .Y(_03359_));
 sky130_fd_sc_hd__mux2_8 _16999_ (.A0(net66),
    .A1(net101),
    .S(net1803),
    .X(_03360_));
 sky130_fd_sc_hd__o21bai_4 _17000_ (.A1(_03317_),
    .A2(_03360_),
    .B1_N(net2006),
    .Y(_03361_));
 sky130_fd_sc_hd__a21oi_4 _17001_ (.A1(_03359_),
    .A2(_03361_),
    .B1(net637),
    .Y(_03362_));
 sky130_fd_sc_hd__a211o_1 _17002_ (.A1(net433),
    .A2(net638),
    .B1(_03362_),
    .C1(net2001),
    .X(_00907_));
 sky130_fd_sc_hd__or2_4 _17003_ (.A(\core.fetchProgramCounter[31] ),
    .B(net996),
    .X(_03363_));
 sky130_fd_sc_hd__a21o_1 _17004_ (.A1(\core.registers[0][31] ),
    .A2(net1027),
    .B1(net1023),
    .X(_03364_));
 sky130_fd_sc_hd__o211a_1 _17005_ (.A1(\core.csr.currentInstruction[31] ),
    .A2(net994),
    .B1(_03312_),
    .C1(_03364_),
    .X(_03365_));
 sky130_fd_sc_hd__o211a_1 _17006_ (.A1(net1032),
    .A2(_02842_),
    .B1(_03363_),
    .C1(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__a21oi_1 _17007_ (.A1(_07864_),
    .A2(_03108_),
    .B1(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__o21ai_2 _17008_ (.A1(net898),
    .A2(_03366_),
    .B1(net1304),
    .Y(_03368_));
 sky130_fd_sc_hd__mux2_8 _17009_ (.A0(net67),
    .A1(net102),
    .S(net1803),
    .X(_03369_));
 sky130_fd_sc_hd__o21bai_4 _17010_ (.A1(_03317_),
    .A2(_03369_),
    .B1_N(net2006),
    .Y(_03370_));
 sky130_fd_sc_hd__a21oi_4 _17011_ (.A1(_03368_),
    .A2(_03370_),
    .B1(net637),
    .Y(_03371_));
 sky130_fd_sc_hd__a211o_1 _17012_ (.A1(net434),
    .A2(net638),
    .B1(_03371_),
    .C1(net2000),
    .X(_00908_));
 sky130_fd_sc_hd__a211oi_1 _17013_ (.A1(_04400_),
    .A2(_03097_),
    .B1(_07839_),
    .C1(net1981),
    .Y(_00909_));
 sky130_fd_sc_hd__nand2_1 _17014_ (.A(net214),
    .B(net251),
    .Y(_03372_));
 sky130_fd_sc_hd__nor3_1 _17015_ (.A(net1981),
    .B(_07837_),
    .C(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__a41o_1 _17016_ (.A1(net442),
    .A2(net1932),
    .A3(_07837_),
    .A4(_07838_),
    .B1(net1350),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _17017_ (.A0(\wbSRAMInterface.currentAddress[0] ),
    .A1(net190),
    .S(net1350),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _17018_ (.A0(\wbSRAMInterface.currentAddress[1] ),
    .A1(net201),
    .S(net1350),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _17019_ (.A0(\wbSRAMInterface.currentAddress[2] ),
    .A1(net206),
    .S(net1350),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _17020_ (.A0(\wbSRAMInterface.currentAddress[3] ),
    .A1(net207),
    .S(net1350),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _17021_ (.A0(\wbSRAMInterface.currentAddress[4] ),
    .A1(net208),
    .S(net1350),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _17022_ (.A0(\wbSRAMInterface.currentAddress[5] ),
    .A1(net209),
    .S(net1351),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _17023_ (.A0(\wbSRAMInterface.currentAddress[6] ),
    .A1(net210),
    .S(net1351),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _17024_ (.A0(\wbSRAMInterface.currentAddress[7] ),
    .A1(net211),
    .S(net1351),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _17025_ (.A0(\wbSRAMInterface.currentAddress[8] ),
    .A1(net212),
    .S(net1351),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _17026_ (.A0(\wbSRAMInterface.currentAddress[9] ),
    .A1(net213),
    .S(net1351),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _17027_ (.A0(\wbSRAMInterface.currentAddress[10] ),
    .A1(net191),
    .S(net1352),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _17028_ (.A0(\wbSRAMInterface.currentAddress[11] ),
    .A1(net192),
    .S(net1352),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _17029_ (.A0(\wbSRAMInterface.currentAddress[12] ),
    .A1(net193),
    .S(net1352),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _17030_ (.A0(\wbSRAMInterface.currentAddress[13] ),
    .A1(net194),
    .S(net1352),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _17031_ (.A0(\wbSRAMInterface.currentAddress[14] ),
    .A1(net195),
    .S(net1352),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _17032_ (.A0(\wbSRAMInterface.currentAddress[15] ),
    .A1(net196),
    .S(net1352),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _17033_ (.A0(\wbSRAMInterface.currentAddress[16] ),
    .A1(net197),
    .S(net1352),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _17034_ (.A0(\wbSRAMInterface.currentAddress[17] ),
    .A1(net198),
    .S(net1352),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _17035_ (.A0(\wbSRAMInterface.currentAddress[18] ),
    .A1(net199),
    .S(net1353),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _17036_ (.A0(\wbSRAMInterface.currentAddress[19] ),
    .A1(net200),
    .S(net1353),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _17037_ (.A0(\wbSRAMInterface.currentAddress[20] ),
    .A1(net202),
    .S(net1353),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _17038_ (.A0(\wbSRAMInterface.currentAddress[21] ),
    .A1(net203),
    .S(net1353),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _17039_ (.A0(\wbSRAMInterface.currentAddress[22] ),
    .A1(net204),
    .S(net1352),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _17040_ (.A0(\wbSRAMInterface.currentAddress[23] ),
    .A1(net205),
    .S(net1352),
    .X(_00934_));
 sky130_fd_sc_hd__nor2_1 _17041_ (.A(net1990),
    .B(_08100_),
    .Y(_00935_));
 sky130_fd_sc_hd__o21ai_1 _17042_ (.A1(\wbSRAMInterface.state[0] ),
    .A2(_03097_),
    .B1(\wbSRAMInterface.state[1] ),
    .Y(_03374_));
 sky130_fd_sc_hd__a31o_1 _17043_ (.A1(net214),
    .A2(net251),
    .A3(net252),
    .B1(_07837_),
    .X(_03375_));
 sky130_fd_sc_hd__and3_1 _17044_ (.A(net1932),
    .B(_03374_),
    .C(_03375_),
    .X(_00936_));
 sky130_fd_sc_hd__o21ba_1 _17045_ (.A1(net252),
    .A2(_03372_),
    .B1_N(_07837_),
    .X(_03376_));
 sky130_fd_sc_hd__a211o_1 _17046_ (.A1(\wbSRAMInterface.state[1] ),
    .A2(\wbSRAMInterface.state[0] ),
    .B1(net1981),
    .C1(_03376_),
    .X(_03377_));
 sky130_fd_sc_hd__a21oi_1 _17047_ (.A1(\wbSRAMInterface.state[0] ),
    .A2(_03097_),
    .B1(_03377_),
    .Y(_00937_));
 sky130_fd_sc_hd__nor2_1 _17048_ (.A(_09086_),
    .B(_09097_),
    .Y(_03378_));
 sky130_fd_sc_hd__and3_4 _17049_ (.A(net676),
    .B(net1073),
    .C(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__mux2_1 _17050_ (.A0(\core.registers[22][0] ),
    .A1(net1038),
    .S(net554),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _17051_ (.A0(\core.registers[22][1] ),
    .A1(net1040),
    .S(net554),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _17052_ (.A0(\core.registers[22][2] ),
    .A1(net1044),
    .S(net555),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _17053_ (.A0(\core.registers[22][3] ),
    .A1(net1048),
    .S(net554),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _17054_ (.A0(\core.registers[22][4] ),
    .A1(net1054),
    .S(net554),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _17055_ (.A0(\core.registers[22][5] ),
    .A1(net1057),
    .S(net555),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _17056_ (.A0(\core.registers[22][6] ),
    .A1(net1061),
    .S(net555),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _17057_ (.A0(\core.registers[22][7] ),
    .A1(net1132),
    .S(net555),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _17058_ (.A0(\core.registers[22][8] ),
    .A1(net960),
    .S(net555),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _17059_ (.A0(\core.registers[22][9] ),
    .A1(net963),
    .S(net553),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _17060_ (.A0(\core.registers[22][10] ),
    .A1(net968),
    .S(net554),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _17061_ (.A0(\core.registers[22][11] ),
    .A1(net972),
    .S(net553),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _17062_ (.A0(\core.registers[22][12] ),
    .A1(net989),
    .S(net553),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _17063_ (.A0(\core.registers[22][13] ),
    .A1(net986),
    .S(net554),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _17064_ (.A0(\core.registers[22][14] ),
    .A1(net974),
    .S(net554),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _17065_ (.A0(\core.registers[22][15] ),
    .A1(net981),
    .S(net554),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _17066_ (.A0(\core.registers[22][16] ),
    .A1(net1125),
    .S(net552),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _17067_ (.A0(\core.registers[22][17] ),
    .A1(net1129),
    .S(net552),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _17068_ (.A0(\core.registers[22][18] ),
    .A1(net1118),
    .S(net553),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _17069_ (.A0(\core.registers[22][19] ),
    .A1(net1122),
    .S(net552),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _17070_ (.A0(\core.registers[22][20] ),
    .A1(net1138),
    .S(net552),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _17071_ (.A0(\core.registers[22][21] ),
    .A1(net1142),
    .S(net552),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _17072_ (.A0(\core.registers[22][22] ),
    .A1(net1147),
    .S(net553),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _17073_ (.A0(\core.registers[22][23] ),
    .A1(net1151),
    .S(net552),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _17074_ (.A0(\core.registers[22][24] ),
    .A1(net1114),
    .S(net552),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _17075_ (.A0(\core.registers[22][25] ),
    .A1(net1108),
    .S(net552),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _17076_ (.A0(\core.registers[22][26] ),
    .A1(net1102),
    .S(net553),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _17077_ (.A0(\core.registers[22][27] ),
    .A1(net1106),
    .S(net552),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _17078_ (.A0(\core.registers[22][28] ),
    .A1(net1098),
    .S(net552),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _17079_ (.A0(\core.registers[22][29] ),
    .A1(net1092),
    .S(net554),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _17080_ (.A0(\core.registers[22][30] ),
    .A1(net1085),
    .S(net555),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _17081_ (.A0(\core.registers[22][31] ),
    .A1(net1089),
    .S(net554),
    .X(_00969_));
 sky130_fd_sc_hd__nor2_1 _17082_ (.A(_09086_),
    .B(_03040_),
    .Y(_03380_));
 sky130_fd_sc_hd__and3_4 _17083_ (.A(net676),
    .B(net1073),
    .C(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__mux2_1 _17084_ (.A0(\core.registers[21][0] ),
    .A1(net1038),
    .S(net550),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _17085_ (.A0(\core.registers[21][1] ),
    .A1(net1039),
    .S(net550),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _17086_ (.A0(\core.registers[21][2] ),
    .A1(net1044),
    .S(net551),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _17087_ (.A0(\core.registers[21][3] ),
    .A1(net1048),
    .S(net550),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _17088_ (.A0(\core.registers[21][4] ),
    .A1(net1053),
    .S(net550),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _17089_ (.A0(\core.registers[21][5] ),
    .A1(net1057),
    .S(net551),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _17090_ (.A0(\core.registers[21][6] ),
    .A1(net1062),
    .S(net551),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _17091_ (.A0(\core.registers[21][7] ),
    .A1(net1133),
    .S(net551),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _17092_ (.A0(\core.registers[21][8] ),
    .A1(net959),
    .S(net551),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _17093_ (.A0(\core.registers[21][9] ),
    .A1(net962),
    .S(net549),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _17094_ (.A0(\core.registers[21][10] ),
    .A1(net969),
    .S(net550),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _17095_ (.A0(\core.registers[21][11] ),
    .A1(net972),
    .S(net549),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _17096_ (.A0(\core.registers[21][12] ),
    .A1(net989),
    .S(net549),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _17097_ (.A0(\core.registers[21][13] ),
    .A1(net986),
    .S(net550),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _17098_ (.A0(\core.registers[21][14] ),
    .A1(net974),
    .S(net550),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _17099_ (.A0(\core.registers[21][15] ),
    .A1(net981),
    .S(net550),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _17100_ (.A0(\core.registers[21][16] ),
    .A1(net1124),
    .S(net548),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _17101_ (.A0(\core.registers[21][17] ),
    .A1(net1129),
    .S(net548),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _17102_ (.A0(\core.registers[21][18] ),
    .A1(net1116),
    .S(net548),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _17103_ (.A0(\core.registers[21][19] ),
    .A1(net1121),
    .S(net548),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _17104_ (.A0(\core.registers[21][20] ),
    .A1(net1138),
    .S(net548),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _17105_ (.A0(\core.registers[21][21] ),
    .A1(net1142),
    .S(net548),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _17106_ (.A0(\core.registers[21][22] ),
    .A1(net1147),
    .S(net549),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _17107_ (.A0(\core.registers[21][23] ),
    .A1(net1151),
    .S(net548),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _17108_ (.A0(\core.registers[21][24] ),
    .A1(net1115),
    .S(net548),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _17109_ (.A0(\core.registers[21][25] ),
    .A1(net1108),
    .S(net548),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _17110_ (.A0(\core.registers[21][26] ),
    .A1(net1103),
    .S(net549),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _17111_ (.A0(\core.registers[21][27] ),
    .A1(net1106),
    .S(net549),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _17112_ (.A0(\core.registers[21][28] ),
    .A1(net1098),
    .S(net548),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _17113_ (.A0(\core.registers[21][29] ),
    .A1(net1092),
    .S(net550),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _17114_ (.A0(\core.registers[21][30] ),
    .A1(net1085),
    .S(net551),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _17115_ (.A0(\core.registers[21][31] ),
    .A1(net1090),
    .S(net550),
    .X(_01001_));
 sky130_fd_sc_hd__nor2_1 _17116_ (.A(_09093_),
    .B(_02932_),
    .Y(_03382_));
 sky130_fd_sc_hd__and3_4 _17117_ (.A(net675),
    .B(net1072),
    .C(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__mux2_1 _17118_ (.A0(\core.registers[15][0] ),
    .A1(net1035),
    .S(net546),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _17119_ (.A0(\core.registers[15][1] ),
    .A1(net1039),
    .S(net545),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _17120_ (.A0(\core.registers[15][2] ),
    .A1(net1043),
    .S(net546),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _17121_ (.A0(\core.registers[15][3] ),
    .A1(net1051),
    .S(net545),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _17122_ (.A0(\core.registers[15][4] ),
    .A1(net1055),
    .S(net545),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _17123_ (.A0(\core.registers[15][5] ),
    .A1(net1059),
    .S(net546),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _17124_ (.A0(\core.registers[15][6] ),
    .A1(net1064),
    .S(net545),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _17125_ (.A0(\core.registers[15][7] ),
    .A1(net1134),
    .S(net545),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _17126_ (.A0(\core.registers[15][8] ),
    .A1(net958),
    .S(net546),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _17127_ (.A0(\core.registers[15][9] ),
    .A1(net963),
    .S(net544),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _17128_ (.A0(\core.registers[15][10] ),
    .A1(net966),
    .S(net546),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _17129_ (.A0(\core.registers[15][11] ),
    .A1(net971),
    .S(net546),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _17130_ (.A0(\core.registers[15][12] ),
    .A1(net987),
    .S(net546),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _17131_ (.A0(\core.registers[15][13] ),
    .A1(net984),
    .S(net545),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _17132_ (.A0(\core.registers[15][14] ),
    .A1(net976),
    .S(net546),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _17133_ (.A0(\core.registers[15][15] ),
    .A1(net980),
    .S(net545),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _17134_ (.A0(\core.registers[15][16] ),
    .A1(net1124),
    .S(net544),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _17135_ (.A0(\core.registers[15][17] ),
    .A1(net1128),
    .S(net544),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _17136_ (.A0(\core.registers[15][18] ),
    .A1(net1116),
    .S(net547),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _17137_ (.A0(\core.registers[15][19] ),
    .A1(net1120),
    .S(net547),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _17138_ (.A0(\core.registers[15][20] ),
    .A1(net1136),
    .S(net544),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _17139_ (.A0(\core.registers[15][21] ),
    .A1(net1140),
    .S(net544),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _17140_ (.A0(\core.registers[15][22] ),
    .A1(net1146),
    .S(net547),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _17141_ (.A0(\core.registers[15][23] ),
    .A1(net1149),
    .S(net544),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _17142_ (.A0(\core.registers[15][24] ),
    .A1(net1112),
    .S(net544),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _17143_ (.A0(\core.registers[15][25] ),
    .A1(net1110),
    .S(net544),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _17144_ (.A0(\core.registers[15][26] ),
    .A1(net1102),
    .S(net547),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _17145_ (.A0(\core.registers[15][27] ),
    .A1(net1105),
    .S(net544),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _17146_ (.A0(\core.registers[15][28] ),
    .A1(net1096),
    .S(net544),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _17147_ (.A0(\core.registers[15][29] ),
    .A1(net1095),
    .S(net545),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _17148_ (.A0(\core.registers[15][30] ),
    .A1(net1086),
    .S(net545),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _17149_ (.A0(\core.registers[15][31] ),
    .A1(net1088),
    .S(net545),
    .X(_01033_));
 sky130_fd_sc_hd__nor2_1 _17150_ (.A(_09097_),
    .B(_02932_),
    .Y(_03384_));
 sky130_fd_sc_hd__and3_4 _17151_ (.A(net675),
    .B(net1072),
    .C(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__mux2_1 _17152_ (.A0(\core.registers[14][0] ),
    .A1(net1035),
    .S(net542),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _17153_ (.A0(\core.registers[14][1] ),
    .A1(net1039),
    .S(net541),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _17154_ (.A0(\core.registers[14][2] ),
    .A1(net1043),
    .S(net542),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _17155_ (.A0(\core.registers[14][3] ),
    .A1(net1051),
    .S(net541),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _17156_ (.A0(\core.registers[14][4] ),
    .A1(net1055),
    .S(net541),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _17157_ (.A0(\core.registers[14][5] ),
    .A1(net1059),
    .S(net542),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _17158_ (.A0(\core.registers[14][6] ),
    .A1(net1064),
    .S(net541),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _17159_ (.A0(\core.registers[14][7] ),
    .A1(net1134),
    .S(net541),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _17160_ (.A0(\core.registers[14][8] ),
    .A1(net958),
    .S(net542),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _17161_ (.A0(\core.registers[14][9] ),
    .A1(net963),
    .S(net540),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _17162_ (.A0(\core.registers[14][10] ),
    .A1(net966),
    .S(net542),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _17163_ (.A0(\core.registers[14][11] ),
    .A1(net971),
    .S(net542),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _17164_ (.A0(\core.registers[14][12] ),
    .A1(net987),
    .S(net542),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _17165_ (.A0(\core.registers[14][13] ),
    .A1(net984),
    .S(net541),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _17166_ (.A0(\core.registers[14][14] ),
    .A1(net976),
    .S(net542),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _17167_ (.A0(\core.registers[14][15] ),
    .A1(net980),
    .S(net541),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _17168_ (.A0(\core.registers[14][16] ),
    .A1(net1124),
    .S(net540),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _17169_ (.A0(\core.registers[14][17] ),
    .A1(net1128),
    .S(net540),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _17170_ (.A0(\core.registers[14][18] ),
    .A1(net1116),
    .S(net543),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _17171_ (.A0(\core.registers[14][19] ),
    .A1(net1120),
    .S(net543),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _17172_ (.A0(\core.registers[14][20] ),
    .A1(net1136),
    .S(net540),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _17173_ (.A0(\core.registers[14][21] ),
    .A1(net1140),
    .S(net540),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _17174_ (.A0(\core.registers[14][22] ),
    .A1(net1146),
    .S(net543),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _17175_ (.A0(\core.registers[14][23] ),
    .A1(net1149),
    .S(net540),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _17176_ (.A0(\core.registers[14][24] ),
    .A1(net1112),
    .S(net540),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _17177_ (.A0(\core.registers[14][25] ),
    .A1(net1110),
    .S(net540),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _17178_ (.A0(\core.registers[14][26] ),
    .A1(net1102),
    .S(net543),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _17179_ (.A0(\core.registers[14][27] ),
    .A1(net1105),
    .S(net540),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _17180_ (.A0(\core.registers[14][28] ),
    .A1(net1096),
    .S(net540),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _17181_ (.A0(\core.registers[14][29] ),
    .A1(net1095),
    .S(net541),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _17182_ (.A0(\core.registers[14][30] ),
    .A1(net1086),
    .S(net541),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _17183_ (.A0(\core.registers[14][31] ),
    .A1(net1088),
    .S(net541),
    .X(_01065_));
 sky130_fd_sc_hd__nor2_1 _17184_ (.A(_02932_),
    .B(_03040_),
    .Y(_03386_));
 sky130_fd_sc_hd__and3_2 _17185_ (.A(net675),
    .B(net1072),
    .C(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__mux2_1 _17186_ (.A0(\core.registers[13][0] ),
    .A1(net1035),
    .S(net538),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _17187_ (.A0(\core.registers[13][1] ),
    .A1(net1041),
    .S(net537),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _17188_ (.A0(\core.registers[13][2] ),
    .A1(net1043),
    .S(net537),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _17189_ (.A0(\core.registers[13][3] ),
    .A1(net1051),
    .S(net537),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _17190_ (.A0(\core.registers[13][4] ),
    .A1(net1055),
    .S(net537),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _17191_ (.A0(\core.registers[13][5] ),
    .A1(net1059),
    .S(net537),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _17192_ (.A0(\core.registers[13][6] ),
    .A1(net1064),
    .S(net537),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _17193_ (.A0(\core.registers[13][7] ),
    .A1(net1134),
    .S(net538),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _17194_ (.A0(\core.registers[13][8] ),
    .A1(net958),
    .S(net537),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _17195_ (.A0(\core.registers[13][9] ),
    .A1(net964),
    .S(net539),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _17196_ (.A0(\core.registers[13][10] ),
    .A1(net967),
    .S(net538),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _17197_ (.A0(\core.registers[13][11] ),
    .A1(net970),
    .S(net538),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _17198_ (.A0(\core.registers[13][12] ),
    .A1(net988),
    .S(net538),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _17199_ (.A0(\core.registers[13][13] ),
    .A1(net984),
    .S(net538),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _17200_ (.A0(\core.registers[13][14] ),
    .A1(net976),
    .S(net538),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _17201_ (.A0(\core.registers[13][15] ),
    .A1(net980),
    .S(net537),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _17202_ (.A0(\core.registers[13][16] ),
    .A1(net1124),
    .S(net536),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _17203_ (.A0(\core.registers[13][17] ),
    .A1(net1128),
    .S(net536),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _17204_ (.A0(\core.registers[13][18] ),
    .A1(net1116),
    .S(net539),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _17205_ (.A0(\core.registers[13][19] ),
    .A1(net1120),
    .S(net536),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _17206_ (.A0(\core.registers[13][20] ),
    .A1(net1136),
    .S(net536),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _17207_ (.A0(\core.registers[13][21] ),
    .A1(net1140),
    .S(net536),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _17208_ (.A0(\core.registers[13][22] ),
    .A1(net1146),
    .S(net539),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _17209_ (.A0(\core.registers[13][23] ),
    .A1(net1150),
    .S(net536),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _17210_ (.A0(\core.registers[13][24] ),
    .A1(net1112),
    .S(net536),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _17211_ (.A0(\core.registers[13][25] ),
    .A1(net1110),
    .S(net536),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _17212_ (.A0(\core.registers[13][26] ),
    .A1(net1101),
    .S(net539),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _17213_ (.A0(\core.registers[13][27] ),
    .A1(net1105),
    .S(net536),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _17214_ (.A0(\core.registers[13][28] ),
    .A1(net1096),
    .S(net536),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _17215_ (.A0(\core.registers[13][29] ),
    .A1(net1095),
    .S(net538),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _17216_ (.A0(\core.registers[13][30] ),
    .A1(net1086),
    .S(net537),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _17217_ (.A0(\core.registers[13][31] ),
    .A1(net1088),
    .S(net537),
    .X(_01097_));
 sky130_fd_sc_hd__and3_1 _17218_ (.A(_07867_),
    .B(_03103_),
    .C(_03106_),
    .X(_03388_));
 sky130_fd_sc_hd__nand3_2 _17219_ (.A(_07867_),
    .B(_03103_),
    .C(_03106_),
    .Y(_03389_));
 sky130_fd_sc_hd__or2_1 _17220_ (.A(\core.management_interruptEnable ),
    .B(_03388_),
    .X(_03390_));
 sky130_fd_sc_hd__o211a_1 _17221_ (.A1(_08786_),
    .A2(_03389_),
    .B1(_03390_),
    .C1(net1934),
    .X(_01098_));
 sky130_fd_sc_hd__or2_1 _17222_ (.A(\coreManagement.control[1] ),
    .B(_03388_),
    .X(_03391_));
 sky130_fd_sc_hd__o211a_1 _17223_ (.A1(_08779_),
    .A2(_03389_),
    .B1(_03391_),
    .C1(net1934),
    .X(_01099_));
 sky130_fd_sc_hd__or2_1 _17224_ (.A(net1789),
    .B(_03388_),
    .X(_03392_));
 sky130_fd_sc_hd__o211a_1 _17225_ (.A1(_08770_),
    .A2(_03389_),
    .B1(_03392_),
    .C1(net1934),
    .X(_01100_));
 sky130_fd_sc_hd__nor2_8 _17226_ (.A(_04398_),
    .B(_08625_),
    .Y(_03393_));
 sky130_fd_sc_hd__nor2_2 _17227_ (.A(\jtag.state[3] ),
    .B(\jtag.state[2] ),
    .Y(_03394_));
 sky130_fd_sc_hd__or2_1 _17228_ (.A(\jtag.state[3] ),
    .B(\jtag.state[2] ),
    .X(_03395_));
 sky130_fd_sc_hd__and3_4 _17229_ (.A(net1778),
    .B(net1780),
    .C(_03394_),
    .X(_03396_));
 sky130_fd_sc_hd__nand3_4 _17230_ (.A(net1778),
    .B(net1780),
    .C(_03394_),
    .Y(_03397_));
 sky130_fd_sc_hd__or2_4 _17231_ (.A(_08634_),
    .B(_03396_),
    .X(_03398_));
 sky130_fd_sc_hd__and2_2 _17232_ (.A(_03393_),
    .B(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__nand2_1 _17233_ (.A(_03393_),
    .B(_03398_),
    .Y(_03400_));
 sky130_fd_sc_hd__and2_1 _17234_ (.A(_03393_),
    .B(_03396_),
    .X(_03401_));
 sky130_fd_sc_hd__nand2_4 _17235_ (.A(_03393_),
    .B(_03396_),
    .Y(_03402_));
 sky130_fd_sc_hd__nand2_1 _17236_ (.A(net188),
    .B(net1342),
    .Y(_03403_));
 sky130_fd_sc_hd__a221o_1 _17237_ (.A1(net188),
    .A2(net1347),
    .B1(net1198),
    .B2(net447),
    .C1(net1200),
    .X(_03404_));
 sky130_fd_sc_hd__o211a_1 _17238_ (.A1(\jtag.dataIDRegister.data[0] ),
    .A2(net1203),
    .B1(_03404_),
    .C1(net1949),
    .X(_01101_));
 sky130_fd_sc_hd__and3_1 _17239_ (.A(net253),
    .B(net1366),
    .C(net1198),
    .X(_03405_));
 sky130_fd_sc_hd__a21o_1 _17240_ (.A1(\jtag.dataIDRegister.data[0] ),
    .A2(_03402_),
    .B1(net1200),
    .X(_03406_));
 sky130_fd_sc_hd__o221a_1 _17241_ (.A1(\jtag.dataIDRegister.data[1] ),
    .A2(net1203),
    .B1(_03405_),
    .B2(_03406_),
    .C1(net1949),
    .X(_01102_));
 sky130_fd_sc_hd__and3_1 _17242_ (.A(net255),
    .B(net1364),
    .C(net1195),
    .X(_03407_));
 sky130_fd_sc_hd__a21o_1 _17243_ (.A1(\jtag.dataIDRegister.data[1] ),
    .A2(_03402_),
    .B1(net1200),
    .X(_03408_));
 sky130_fd_sc_hd__o221a_1 _17244_ (.A1(\jtag.dataIDRegister.data[2] ),
    .A2(net1203),
    .B1(_03407_),
    .B2(_03408_),
    .C1(net1950),
    .X(_01103_));
 sky130_fd_sc_hd__and3_1 _17245_ (.A(net256),
    .B(net1364),
    .C(net1195),
    .X(_03409_));
 sky130_fd_sc_hd__a21o_1 _17246_ (.A1(\jtag.dataIDRegister.data[2] ),
    .A2(_03402_),
    .B1(net1199),
    .X(_03410_));
 sky130_fd_sc_hd__o221a_1 _17247_ (.A1(\jtag.dataIDRegister.data[3] ),
    .A2(net1203),
    .B1(_03409_),
    .B2(_03410_),
    .C1(net1950),
    .X(_01104_));
 sky130_fd_sc_hd__and3_1 _17248_ (.A(net257),
    .B(net1363),
    .C(net1195),
    .X(_03411_));
 sky130_fd_sc_hd__a21o_1 _17249_ (.A1(\jtag.dataIDRegister.data[3] ),
    .A2(_03402_),
    .B1(net1199),
    .X(_03412_));
 sky130_fd_sc_hd__o221a_1 _17250_ (.A1(\jtag.dataIDRegister.data[4] ),
    .A2(net1203),
    .B1(_03411_),
    .B2(_03412_),
    .C1(net1950),
    .X(_01105_));
 sky130_fd_sc_hd__and3_1 _17251_ (.A(net258),
    .B(net1363),
    .C(net1195),
    .X(_03413_));
 sky130_fd_sc_hd__a21o_1 _17252_ (.A1(\jtag.dataIDRegister.data[4] ),
    .A2(_03402_),
    .B1(net1200),
    .X(_03414_));
 sky130_fd_sc_hd__o221a_1 _17253_ (.A1(\jtag.dataIDRegister.data[5] ),
    .A2(net1203),
    .B1(_03413_),
    .B2(_03414_),
    .C1(net1950),
    .X(_01106_));
 sky130_fd_sc_hd__and3_1 _17254_ (.A(net259),
    .B(net1363),
    .C(net1195),
    .X(_03415_));
 sky130_fd_sc_hd__a21o_1 _17255_ (.A1(\jtag.dataIDRegister.data[5] ),
    .A2(_03402_),
    .B1(net1200),
    .X(_03416_));
 sky130_fd_sc_hd__o221a_1 _17256_ (.A1(\jtag.dataIDRegister.data[6] ),
    .A2(net1203),
    .B1(_03415_),
    .B2(_03416_),
    .C1(net1950),
    .X(_01107_));
 sky130_fd_sc_hd__and3_1 _17257_ (.A(net260),
    .B(net1363),
    .C(net1195),
    .X(_03417_));
 sky130_fd_sc_hd__a21o_1 _17258_ (.A1(\jtag.dataIDRegister.data[6] ),
    .A2(_03402_),
    .B1(net1199),
    .X(_03418_));
 sky130_fd_sc_hd__o221a_1 _17259_ (.A1(\jtag.dataIDRegister.data[7] ),
    .A2(net1203),
    .B1(_03417_),
    .B2(_03418_),
    .C1(net1950),
    .X(_01108_));
 sky130_fd_sc_hd__nand2b_1 _17260_ (.A_N(net261),
    .B(net1363),
    .Y(_03419_));
 sky130_fd_sc_hd__a221o_1 _17261_ (.A1(\jtag.dataIDRegister.data[7] ),
    .A2(net1345),
    .B1(net1195),
    .B2(_03419_),
    .C1(net1199),
    .X(_03420_));
 sky130_fd_sc_hd__o211a_1 _17262_ (.A1(\jtag.dataIDRegister.data[8] ),
    .A2(net1204),
    .B1(_03420_),
    .C1(net1951),
    .X(_01109_));
 sky130_fd_sc_hd__and3_1 _17263_ (.A(net262),
    .B(net1363),
    .C(net1195),
    .X(_03421_));
 sky130_fd_sc_hd__a21o_1 _17264_ (.A1(\jtag.dataIDRegister.data[8] ),
    .A2(net1345),
    .B1(net1199),
    .X(_03422_));
 sky130_fd_sc_hd__o221a_1 _17265_ (.A1(\jtag.dataIDRegister.data[9] ),
    .A2(net1203),
    .B1(_03421_),
    .B2(_03422_),
    .C1(net1950),
    .X(_01110_));
 sky130_fd_sc_hd__and3_1 _17266_ (.A(net263),
    .B(net1363),
    .C(net1195),
    .X(_03423_));
 sky130_fd_sc_hd__a21o_1 _17267_ (.A1(\jtag.dataIDRegister.data[9] ),
    .A2(net1345),
    .B1(net1199),
    .X(_03424_));
 sky130_fd_sc_hd__o221a_1 _17268_ (.A1(\jtag.dataIDRegister.data[10] ),
    .A2(net1203),
    .B1(_03423_),
    .B2(_03424_),
    .C1(net1950),
    .X(_01111_));
 sky130_fd_sc_hd__and3_1 _17269_ (.A(net254),
    .B(net1363),
    .C(net1195),
    .X(_03425_));
 sky130_fd_sc_hd__a211o_1 _17270_ (.A1(\jtag.dataIDRegister.data[10] ),
    .A2(net1345),
    .B1(net1199),
    .C1(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__o211a_1 _17271_ (.A1(\jtag.dataIDRegister.data[11] ),
    .A2(net1204),
    .B1(_03426_),
    .C1(net1950),
    .X(_01112_));
 sky130_fd_sc_hd__and3_1 _17272_ (.A(net264),
    .B(net1363),
    .C(net1196),
    .X(_03427_));
 sky130_fd_sc_hd__a21o_1 _17273_ (.A1(\jtag.dataIDRegister.data[11] ),
    .A2(net1345),
    .B1(net1199),
    .X(_03428_));
 sky130_fd_sc_hd__o221a_1 _17274_ (.A1(\jtag.dataIDRegister.data[12] ),
    .A2(net1204),
    .B1(_03427_),
    .B2(_03428_),
    .C1(net1950),
    .X(_01113_));
 sky130_fd_sc_hd__and3_1 _17275_ (.A(net271),
    .B(net1363),
    .C(net1196),
    .X(_03429_));
 sky130_fd_sc_hd__a211o_1 _17276_ (.A1(\jtag.dataIDRegister.data[12] ),
    .A2(net1345),
    .B1(net1199),
    .C1(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__o211a_1 _17277_ (.A1(\jtag.dataIDRegister.data[13] ),
    .A2(net1204),
    .B1(_03430_),
    .C1(net1951),
    .X(_01114_));
 sky130_fd_sc_hd__nand2b_1 _17278_ (.A_N(net272),
    .B(net1364),
    .Y(_03431_));
 sky130_fd_sc_hd__a221o_1 _17279_ (.A1(\jtag.dataIDRegister.data[13] ),
    .A2(net1345),
    .B1(net1196),
    .B2(_03431_),
    .C1(net1199),
    .X(_03432_));
 sky130_fd_sc_hd__o211a_1 _17280_ (.A1(\jtag.dataIDRegister.data[14] ),
    .A2(net1204),
    .B1(_03432_),
    .C1(net1951),
    .X(_01115_));
 sky130_fd_sc_hd__and3_1 _17281_ (.A(net273),
    .B(net1364),
    .C(net1196),
    .X(_03433_));
 sky130_fd_sc_hd__a21o_1 _17282_ (.A1(\jtag.dataIDRegister.data[14] ),
    .A2(net1345),
    .B1(net1200),
    .X(_03434_));
 sky130_fd_sc_hd__o221a_1 _17283_ (.A1(\jtag.dataIDRegister.data[15] ),
    .A2(net1205),
    .B1(_03433_),
    .B2(_03434_),
    .C1(net1951),
    .X(_01116_));
 sky130_fd_sc_hd__and3_1 _17284_ (.A(net274),
    .B(net1364),
    .C(net1196),
    .X(_03435_));
 sky130_fd_sc_hd__a211o_1 _17285_ (.A1(\jtag.dataIDRegister.data[15] ),
    .A2(net1345),
    .B1(net1200),
    .C1(_03435_),
    .X(_03436_));
 sky130_fd_sc_hd__o211a_1 _17286_ (.A1(\jtag.dataIDRegister.data[16] ),
    .A2(net1205),
    .B1(_03436_),
    .C1(net1951),
    .X(_01117_));
 sky130_fd_sc_hd__and3_1 _17287_ (.A(net275),
    .B(net1364),
    .C(net1196),
    .X(_03437_));
 sky130_fd_sc_hd__a21o_1 _17288_ (.A1(\jtag.dataIDRegister.data[16] ),
    .A2(net1346),
    .B1(net1200),
    .X(_03438_));
 sky130_fd_sc_hd__o221a_1 _17289_ (.A1(\jtag.dataIDRegister.data[17] ),
    .A2(net1205),
    .B1(_03437_),
    .B2(_03438_),
    .C1(net1951),
    .X(_01118_));
 sky130_fd_sc_hd__and3_1 _17290_ (.A(net276),
    .B(net1364),
    .C(net1196),
    .X(_03439_));
 sky130_fd_sc_hd__a21o_1 _17291_ (.A1(\jtag.dataIDRegister.data[17] ),
    .A2(net1346),
    .B1(net1200),
    .X(_03440_));
 sky130_fd_sc_hd__o221a_1 _17292_ (.A1(\jtag.dataIDRegister.data[18] ),
    .A2(net1205),
    .B1(_03439_),
    .B2(_03440_),
    .C1(net1951),
    .X(_01119_));
 sky130_fd_sc_hd__and3_1 _17293_ (.A(net277),
    .B(net1365),
    .C(net1197),
    .X(_03441_));
 sky130_fd_sc_hd__a21o_1 _17294_ (.A1(\jtag.dataIDRegister.data[18] ),
    .A2(net1346),
    .B1(net1201),
    .X(_03442_));
 sky130_fd_sc_hd__o221a_1 _17295_ (.A1(\jtag.dataIDRegister.data[19] ),
    .A2(net1206),
    .B1(_03441_),
    .B2(_03442_),
    .C1(net1957),
    .X(_01120_));
 sky130_fd_sc_hd__and3_1 _17296_ (.A(net278),
    .B(net1365),
    .C(net1197),
    .X(_03443_));
 sky130_fd_sc_hd__a21o_1 _17297_ (.A1(\jtag.dataIDRegister.data[19] ),
    .A2(net1346),
    .B1(net1201),
    .X(_03444_));
 sky130_fd_sc_hd__o221a_1 _17298_ (.A1(\jtag.dataIDRegister.data[20] ),
    .A2(net1206),
    .B1(_03443_),
    .B2(_03444_),
    .C1(net1957),
    .X(_01121_));
 sky130_fd_sc_hd__and3_1 _17299_ (.A(net279),
    .B(net1365),
    .C(net1197),
    .X(_03445_));
 sky130_fd_sc_hd__a21o_1 _17300_ (.A1(\jtag.dataIDRegister.data[20] ),
    .A2(net1346),
    .B1(net1201),
    .X(_03446_));
 sky130_fd_sc_hd__o221a_1 _17301_ (.A1(\jtag.dataIDRegister.data[21] ),
    .A2(net1206),
    .B1(_03445_),
    .B2(_03446_),
    .C1(net1957),
    .X(_01122_));
 sky130_fd_sc_hd__and3_1 _17302_ (.A(net265),
    .B(net1365),
    .C(net1198),
    .X(_03447_));
 sky130_fd_sc_hd__a211o_1 _17303_ (.A1(\jtag.dataIDRegister.data[21] ),
    .A2(net1347),
    .B1(net1202),
    .C1(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__o211a_1 _17304_ (.A1(\jtag.dataIDRegister.data[22] ),
    .A2(net1206),
    .B1(_03448_),
    .C1(net1957),
    .X(_01123_));
 sky130_fd_sc_hd__and3_1 _17305_ (.A(net266),
    .B(net1365),
    .C(net1197),
    .X(_03449_));
 sky130_fd_sc_hd__a21o_1 _17306_ (.A1(\jtag.dataIDRegister.data[22] ),
    .A2(net1347),
    .B1(net1202),
    .X(_03450_));
 sky130_fd_sc_hd__o221a_1 _17307_ (.A1(\jtag.dataIDRegister.data[23] ),
    .A2(net1206),
    .B1(_03449_),
    .B2(_03450_),
    .C1(net1957),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _17308_ (.A0(net1),
    .A1(net267),
    .S(net1365),
    .X(_03451_));
 sky130_fd_sc_hd__a221o_1 _17309_ (.A1(\jtag.dataIDRegister.data[23] ),
    .A2(net1347),
    .B1(net1197),
    .B2(_03451_),
    .C1(net1201),
    .X(_03452_));
 sky130_fd_sc_hd__o211a_1 _17310_ (.A1(\jtag.dataIDRegister.data[24] ),
    .A2(net1206),
    .B1(_03452_),
    .C1(net1959),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _17311_ (.A0(net2),
    .A1(net268),
    .S(net1365),
    .X(_03453_));
 sky130_fd_sc_hd__a221o_1 _17312_ (.A1(\jtag.dataIDRegister.data[24] ),
    .A2(net1347),
    .B1(net1197),
    .B2(_03453_),
    .C1(net1201),
    .X(_03454_));
 sky130_fd_sc_hd__o211a_1 _17313_ (.A1(\jtag.dataIDRegister.data[25] ),
    .A2(net1206),
    .B1(_03454_),
    .C1(net1957),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _17314_ (.A0(net3),
    .A1(net269),
    .S(net1366),
    .X(_03455_));
 sky130_fd_sc_hd__a221o_1 _17315_ (.A1(\jtag.dataIDRegister.data[25] ),
    .A2(net1347),
    .B1(net1197),
    .B2(_03455_),
    .C1(net1201),
    .X(_03456_));
 sky130_fd_sc_hd__o211a_1 _17316_ (.A1(\jtag.dataIDRegister.data[26] ),
    .A2(net1206),
    .B1(_03456_),
    .C1(net1959),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _17317_ (.A0(net4),
    .A1(net270),
    .S(net1366),
    .X(_03457_));
 sky130_fd_sc_hd__a221o_1 _17318_ (.A1(\jtag.dataIDRegister.data[26] ),
    .A2(net1347),
    .B1(net1197),
    .B2(_03457_),
    .C1(net1201),
    .X(_03458_));
 sky130_fd_sc_hd__o211a_1 _17319_ (.A1(\jtag.dataIDRegister.data[27] ),
    .A2(_03399_),
    .B1(_03458_),
    .C1(net1957),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _17320_ (.A0(net5),
    .A1(net280),
    .S(net1366),
    .X(_03459_));
 sky130_fd_sc_hd__a221o_1 _17321_ (.A1(\jtag.dataIDRegister.data[27] ),
    .A2(net1347),
    .B1(net1197),
    .B2(_03459_),
    .C1(net1201),
    .X(_03460_));
 sky130_fd_sc_hd__o211a_1 _17322_ (.A1(\jtag.dataIDRegister.data[28] ),
    .A2(net1206),
    .B1(_03460_),
    .C1(net1959),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _17323_ (.A0(net6),
    .A1(net281),
    .S(net1365),
    .X(_03461_));
 sky130_fd_sc_hd__a221o_1 _17324_ (.A1(\jtag.dataIDRegister.data[28] ),
    .A2(net1348),
    .B1(net1198),
    .B2(_03461_),
    .C1(net1202),
    .X(_03462_));
 sky130_fd_sc_hd__o211a_1 _17325_ (.A1(\jtag.dataIDRegister.data[29] ),
    .A2(_03399_),
    .B1(_03462_),
    .C1(net1957),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _17326_ (.A0(net7),
    .A1(net282),
    .S(net1365),
    .X(_03463_));
 sky130_fd_sc_hd__a221o_1 _17327_ (.A1(\jtag.dataIDRegister.data[29] ),
    .A2(net1346),
    .B1(net1198),
    .B2(_03463_),
    .C1(net1201),
    .X(_03464_));
 sky130_fd_sc_hd__o211a_1 _17328_ (.A1(\jtag.dataIDRegister.data[30] ),
    .A2(net1206),
    .B1(_03464_),
    .C1(net1957),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _17329_ (.A0(net8),
    .A1(net283),
    .S(net1365),
    .X(_03465_));
 sky130_fd_sc_hd__a221o_1 _17330_ (.A1(\jtag.dataIDRegister.data[30] ),
    .A2(net1345),
    .B1(net1197),
    .B2(_03465_),
    .C1(net1201),
    .X(_03466_));
 sky130_fd_sc_hd__o211a_1 _17331_ (.A1(\jtag.dataIDRegister.data[31] ),
    .A2(net1205),
    .B1(_03466_),
    .C1(net1951),
    .X(_01132_));
 sky130_fd_sc_hd__a31o_1 _17332_ (.A1(net1781),
    .A2(_08627_),
    .A3(_08634_),
    .B1(\jtag.dataBypassRegister.data ),
    .X(_03467_));
 sky130_fd_sc_hd__a41o_1 _17333_ (.A1(net1781),
    .A2(_08627_),
    .A3(_03398_),
    .A4(_03403_),
    .B1(net1961),
    .X(_03468_));
 sky130_fd_sc_hd__and2b_1 _17334_ (.A_N(_03468_),
    .B(_03467_),
    .X(_01133_));
 sky130_fd_sc_hd__and3_4 _17335_ (.A(net1781),
    .B(_08630_),
    .C(_03398_),
    .X(_03469_));
 sky130_fd_sc_hd__nand2b_4 _17336_ (.A_N(_09061_),
    .B(_03398_),
    .Y(_03470_));
 sky130_fd_sc_hd__nor2_8 _17337_ (.A(_09061_),
    .B(net1342),
    .Y(_03471_));
 sky130_fd_sc_hd__a221o_1 _17338_ (.A1(net188),
    .A2(net1349),
    .B1(net1244),
    .B2(\jtag.managementReadData[0] ),
    .C1(net1248),
    .X(_03472_));
 sky130_fd_sc_hd__o211a_1 _17339_ (.A1(\jtag.dataBSRRegister.data[0] ),
    .A2(net1253),
    .B1(_03472_),
    .C1(net1932),
    .X(_01134_));
 sky130_fd_sc_hd__a221o_1 _17340_ (.A1(\jtag.dataBSRRegister.data[0] ),
    .A2(net1349),
    .B1(net1245),
    .B2(\jtag.managementReadData[1] ),
    .C1(net1249),
    .X(_03473_));
 sky130_fd_sc_hd__o211a_1 _17341_ (.A1(\jtag.dataBSRRegister.data[1] ),
    .A2(net1253),
    .B1(_03473_),
    .C1(net1933),
    .X(_01135_));
 sky130_fd_sc_hd__a221o_1 _17342_ (.A1(\jtag.dataBSRRegister.data[1] ),
    .A2(net1349),
    .B1(net1244),
    .B2(\jtag.managementReadData[2] ),
    .C1(net1248),
    .X(_03474_));
 sky130_fd_sc_hd__o211a_1 _17343_ (.A1(\jtag.dataBSRRegister.data[2] ),
    .A2(net1252),
    .B1(_03474_),
    .C1(net1933),
    .X(_01136_));
 sky130_fd_sc_hd__a221o_1 _17344_ (.A1(\jtag.dataBSRRegister.data[2] ),
    .A2(net1349),
    .B1(net1245),
    .B2(\jtag.managementReadData[3] ),
    .C1(net1249),
    .X(_03475_));
 sky130_fd_sc_hd__o211a_1 _17345_ (.A1(\jtag.dataBSRRegister.data[3] ),
    .A2(net1252),
    .B1(_03475_),
    .C1(net1936),
    .X(_01137_));
 sky130_fd_sc_hd__a221o_1 _17346_ (.A1(\jtag.dataBSRRegister.data[3] ),
    .A2(net1349),
    .B1(net1245),
    .B2(\jtag.managementReadData[4] ),
    .C1(net1249),
    .X(_03476_));
 sky130_fd_sc_hd__o211a_1 _17347_ (.A1(\jtag.dataBSRRegister.data[4] ),
    .A2(net1252),
    .B1(_03476_),
    .C1(net1935),
    .X(_01138_));
 sky130_fd_sc_hd__a221o_1 _17348_ (.A1(\jtag.dataBSRRegister.data[4] ),
    .A2(net1348),
    .B1(net1244),
    .B2(\jtag.managementReadData[5] ),
    .C1(net1248),
    .X(_03477_));
 sky130_fd_sc_hd__o211a_1 _17349_ (.A1(\jtag.dataBSRRegister.data[5] ),
    .A2(net1252),
    .B1(_03477_),
    .C1(net1953),
    .X(_01139_));
 sky130_fd_sc_hd__a221o_1 _17350_ (.A1(\jtag.dataBSRRegister.data[5] ),
    .A2(net1348),
    .B1(net1244),
    .B2(\jtag.managementReadData[6] ),
    .C1(net1248),
    .X(_03478_));
 sky130_fd_sc_hd__o211a_1 _17351_ (.A1(\jtag.dataBSRRegister.data[6] ),
    .A2(net1252),
    .B1(_03478_),
    .C1(net1953),
    .X(_01140_));
 sky130_fd_sc_hd__a221o_1 _17352_ (.A1(\jtag.dataBSRRegister.data[6] ),
    .A2(net1348),
    .B1(net1244),
    .B2(\jtag.managementReadData[7] ),
    .C1(net1248),
    .X(_03479_));
 sky130_fd_sc_hd__o211a_1 _17353_ (.A1(\jtag.dataBSRRegister.data[7] ),
    .A2(net1252),
    .B1(_03479_),
    .C1(net1953),
    .X(_01141_));
 sky130_fd_sc_hd__a221o_1 _17354_ (.A1(\jtag.dataBSRRegister.data[7] ),
    .A2(net1348),
    .B1(net1244),
    .B2(\jtag.managementReadData[8] ),
    .C1(net1248),
    .X(_03480_));
 sky130_fd_sc_hd__o211a_1 _17355_ (.A1(\jtag.dataBSRRegister.data[8] ),
    .A2(net1252),
    .B1(_03480_),
    .C1(net1953),
    .X(_01142_));
 sky130_fd_sc_hd__a221o_1 _17356_ (.A1(\jtag.dataBSRRegister.data[8] ),
    .A2(net1348),
    .B1(net1244),
    .B2(\jtag.managementReadData[9] ),
    .C1(net1248),
    .X(_03481_));
 sky130_fd_sc_hd__o211a_1 _17357_ (.A1(\jtag.dataBSRRegister.data[9] ),
    .A2(net1253),
    .B1(_03481_),
    .C1(net1954),
    .X(_01143_));
 sky130_fd_sc_hd__a221o_1 _17358_ (.A1(\jtag.dataBSRRegister.data[9] ),
    .A2(net1349),
    .B1(net1244),
    .B2(\jtag.managementReadData[10] ),
    .C1(net1248),
    .X(_03482_));
 sky130_fd_sc_hd__o211a_1 _17359_ (.A1(\jtag.dataBSRRegister.data[10] ),
    .A2(net1252),
    .B1(_03482_),
    .C1(net1936),
    .X(_01144_));
 sky130_fd_sc_hd__a221o_1 _17360_ (.A1(\jtag.dataBSRRegister.data[10] ),
    .A2(net1349),
    .B1(net1244),
    .B2(\jtag.managementReadData[11] ),
    .C1(net1248),
    .X(_03483_));
 sky130_fd_sc_hd__o211a_1 _17361_ (.A1(\jtag.dataBSRRegister.data[11] ),
    .A2(net1252),
    .B1(_03483_),
    .C1(net1936),
    .X(_01145_));
 sky130_fd_sc_hd__a221o_1 _17362_ (.A1(\jtag.dataBSRRegister.data[11] ),
    .A2(net1349),
    .B1(net1244),
    .B2(\jtag.managementReadData[12] ),
    .C1(net1248),
    .X(_03484_));
 sky130_fd_sc_hd__o211a_1 _17363_ (.A1(\jtag.dataBSRRegister.data[12] ),
    .A2(net1252),
    .B1(_03484_),
    .C1(net1937),
    .X(_01146_));
 sky130_fd_sc_hd__a221o_1 _17364_ (.A1(\jtag.dataBSRRegister.data[12] ),
    .A2(net1349),
    .B1(net1245),
    .B2(\jtag.managementReadData[13] ),
    .C1(net1249),
    .X(_03485_));
 sky130_fd_sc_hd__o211a_1 _17365_ (.A1(\jtag.dataBSRRegister.data[13] ),
    .A2(net1253),
    .B1(_03485_),
    .C1(net1933),
    .X(_01147_));
 sky130_fd_sc_hd__a221o_1 _17366_ (.A1(\jtag.dataBSRRegister.data[13] ),
    .A2(net1344),
    .B1(net1245),
    .B2(\jtag.managementReadData[14] ),
    .C1(net1249),
    .X(_03486_));
 sky130_fd_sc_hd__o211a_1 _17367_ (.A1(\jtag.dataBSRRegister.data[14] ),
    .A2(net1253),
    .B1(_03486_),
    .C1(net1917),
    .X(_01148_));
 sky130_fd_sc_hd__a221o_1 _17368_ (.A1(\jtag.dataBSRRegister.data[14] ),
    .A2(net1344),
    .B1(net1245),
    .B2(\jtag.managementReadData[15] ),
    .C1(net1249),
    .X(_03487_));
 sky130_fd_sc_hd__o211a_1 _17369_ (.A1(\jtag.dataBSRRegister.data[15] ),
    .A2(net1253),
    .B1(_03487_),
    .C1(net1916),
    .X(_01149_));
 sky130_fd_sc_hd__a221o_1 _17370_ (.A1(\jtag.dataBSRRegister.data[15] ),
    .A2(net1344),
    .B1(net1245),
    .B2(\jtag.managementReadData[16] ),
    .C1(net1249),
    .X(_03488_));
 sky130_fd_sc_hd__o211a_1 _17371_ (.A1(\jtag.dataBSRRegister.data[16] ),
    .A2(net1253),
    .B1(_03488_),
    .C1(net1916),
    .X(_01150_));
 sky130_fd_sc_hd__a221o_1 _17372_ (.A1(\jtag.dataBSRRegister.data[16] ),
    .A2(net1344),
    .B1(net1243),
    .B2(\jtag.managementReadData[17] ),
    .C1(net1247),
    .X(_03489_));
 sky130_fd_sc_hd__o211a_1 _17373_ (.A1(\jtag.dataBSRRegister.data[17] ),
    .A2(net1251),
    .B1(_03489_),
    .C1(net1904),
    .X(_01151_));
 sky130_fd_sc_hd__a221o_1 _17374_ (.A1(\jtag.dataBSRRegister.data[17] ),
    .A2(net1344),
    .B1(net1243),
    .B2(\jtag.managementReadData[18] ),
    .C1(net1247),
    .X(_03490_));
 sky130_fd_sc_hd__o211a_1 _17375_ (.A1(\jtag.dataBSRRegister.data[18] ),
    .A2(net1251),
    .B1(_03490_),
    .C1(net1904),
    .X(_01152_));
 sky130_fd_sc_hd__a221o_1 _17376_ (.A1(\jtag.dataBSRRegister.data[18] ),
    .A2(net1344),
    .B1(net1243),
    .B2(\jtag.managementReadData[19] ),
    .C1(net1247),
    .X(_03491_));
 sky130_fd_sc_hd__o211a_1 _17377_ (.A1(\jtag.dataBSRRegister.data[19] ),
    .A2(net1251),
    .B1(_03491_),
    .C1(net1904),
    .X(_01153_));
 sky130_fd_sc_hd__a221o_4 _17378_ (.A1(\jtag.dataBSRRegister.data[19] ),
    .A2(net1344),
    .B1(net1243),
    .B2(\jtag.managementReadData[20] ),
    .C1(net1247),
    .X(_03492_));
 sky130_fd_sc_hd__o211a_1 _17379_ (.A1(\jtag.dataBSRRegister.data[20] ),
    .A2(net1251),
    .B1(_03492_),
    .C1(net1895),
    .X(_01154_));
 sky130_fd_sc_hd__a221o_1 _17380_ (.A1(\jtag.dataBSRRegister.data[20] ),
    .A2(net1343),
    .B1(net1243),
    .B2(\jtag.managementReadData[21] ),
    .C1(net1247),
    .X(_03493_));
 sky130_fd_sc_hd__o211a_1 _17381_ (.A1(\jtag.dataBSRRegister.data[21] ),
    .A2(net1251),
    .B1(_03493_),
    .C1(net1895),
    .X(_01155_));
 sky130_fd_sc_hd__a221o_1 _17382_ (.A1(\jtag.dataBSRRegister.data[21] ),
    .A2(net1343),
    .B1(net1243),
    .B2(\jtag.managementReadData[22] ),
    .C1(net1246),
    .X(_03494_));
 sky130_fd_sc_hd__o211a_1 _17383_ (.A1(\jtag.dataBSRRegister.data[22] ),
    .A2(net1250),
    .B1(_03494_),
    .C1(net1894),
    .X(_01156_));
 sky130_fd_sc_hd__a221o_1 _17384_ (.A1(\jtag.dataBSRRegister.data[22] ),
    .A2(net1343),
    .B1(net1242),
    .B2(\jtag.managementReadData[23] ),
    .C1(net1246),
    .X(_03495_));
 sky130_fd_sc_hd__o211a_1 _17385_ (.A1(\jtag.dataBSRRegister.data[23] ),
    .A2(net1250),
    .B1(_03495_),
    .C1(net1893),
    .X(_01157_));
 sky130_fd_sc_hd__a221o_1 _17386_ (.A1(\jtag.dataBSRRegister.data[23] ),
    .A2(net1342),
    .B1(net1242),
    .B2(\jtag.managementReadData[24] ),
    .C1(net1246),
    .X(_03496_));
 sky130_fd_sc_hd__o211a_1 _17387_ (.A1(\jtag.dataBSRRegister.data[24] ),
    .A2(net1250),
    .B1(_03496_),
    .C1(net1893),
    .X(_01158_));
 sky130_fd_sc_hd__a221o_1 _17388_ (.A1(\jtag.dataBSRRegister.data[24] ),
    .A2(net1342),
    .B1(net1242),
    .B2(\jtag.managementReadData[25] ),
    .C1(net1246),
    .X(_03497_));
 sky130_fd_sc_hd__o211a_1 _17389_ (.A1(\jtag.dataBSRRegister.data[25] ),
    .A2(net1250),
    .B1(_03497_),
    .C1(net1893),
    .X(_01159_));
 sky130_fd_sc_hd__a221o_1 _17390_ (.A1(\jtag.dataBSRRegister.data[25] ),
    .A2(net1343),
    .B1(net1242),
    .B2(\jtag.managementReadData[26] ),
    .C1(net1246),
    .X(_03498_));
 sky130_fd_sc_hd__o211a_1 _17391_ (.A1(\jtag.dataBSRRegister.data[26] ),
    .A2(net1250),
    .B1(_03498_),
    .C1(net1893),
    .X(_01160_));
 sky130_fd_sc_hd__a221o_1 _17392_ (.A1(\jtag.dataBSRRegister.data[26] ),
    .A2(net1342),
    .B1(net1242),
    .B2(\jtag.managementReadData[27] ),
    .C1(net1246),
    .X(_03499_));
 sky130_fd_sc_hd__o211a_1 _17393_ (.A1(\jtag.dataBSRRegister.data[27] ),
    .A2(net1250),
    .B1(_03499_),
    .C1(net1893),
    .X(_01161_));
 sky130_fd_sc_hd__a221o_1 _17394_ (.A1(\jtag.dataBSRRegister.data[27] ),
    .A2(net1342),
    .B1(net1242),
    .B2(\jtag.managementReadData[28] ),
    .C1(net1246),
    .X(_03500_));
 sky130_fd_sc_hd__o211a_1 _17395_ (.A1(\jtag.dataBSRRegister.data[28] ),
    .A2(net1250),
    .B1(_03500_),
    .C1(net1886),
    .X(_01162_));
 sky130_fd_sc_hd__a221o_1 _17396_ (.A1(\jtag.dataBSRRegister.data[28] ),
    .A2(net1342),
    .B1(net1242),
    .B2(\jtag.managementReadData[29] ),
    .C1(net1246),
    .X(_03501_));
 sky130_fd_sc_hd__o211a_1 _17397_ (.A1(\jtag.dataBSRRegister.data[29] ),
    .A2(net1250),
    .B1(_03501_),
    .C1(net1886),
    .X(_01163_));
 sky130_fd_sc_hd__a221o_1 _17398_ (.A1(\jtag.dataBSRRegister.data[29] ),
    .A2(net1342),
    .B1(net1242),
    .B2(\jtag.managementReadData[30] ),
    .C1(net1246),
    .X(_03502_));
 sky130_fd_sc_hd__o211a_1 _17399_ (.A1(\jtag.dataBSRRegister.data[30] ),
    .A2(net1250),
    .B1(_03502_),
    .C1(net1887),
    .X(_01164_));
 sky130_fd_sc_hd__a221o_1 _17400_ (.A1(\jtag.dataBSRRegister.data[30] ),
    .A2(net1342),
    .B1(net1242),
    .B2(\jtag.managementReadData[31] ),
    .C1(net1246),
    .X(_03503_));
 sky130_fd_sc_hd__o211a_1 _17401_ (.A1(\jtag.dataBSRRegister.data[31] ),
    .A2(net1250),
    .B1(_03503_),
    .C1(net1887),
    .X(_01165_));
 sky130_fd_sc_hd__nand2_2 _17402_ (.A(net1781),
    .B(_08621_),
    .Y(_03504_));
 sky130_fd_sc_hd__a31o_1 _17403_ (.A1(net1781),
    .A2(net1778),
    .A3(_08620_),
    .B1(\jtag.instructionRegister.data[0] ),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_1 _17404_ (.A0(net445),
    .A1(net188),
    .S(net1779),
    .X(_03506_));
 sky130_fd_sc_hd__o211a_1 _17405_ (.A1(_03504_),
    .A2(_03506_),
    .B1(_03505_),
    .C1(net1886),
    .X(_01166_));
 sky130_fd_sc_hd__a31o_1 _17406_ (.A1(net1781),
    .A2(net1778),
    .A3(_08620_),
    .B1(\jtag.instructionRegister.data[1] ),
    .X(_03507_));
 sky130_fd_sc_hd__mux2_1 _17407_ (.A0(net446),
    .A1(\jtag.instructionRegister.data[0] ),
    .S(net1779),
    .X(_03508_));
 sky130_fd_sc_hd__o211a_1 _17408_ (.A1(_03504_),
    .A2(_03508_),
    .B1(_03507_),
    .C1(net1890),
    .X(_01167_));
 sky130_fd_sc_hd__a31o_1 _17409_ (.A1(net1782),
    .A2(net1777),
    .A3(_08620_),
    .B1(\jtag.instructionRegister.data[2] ),
    .X(_03509_));
 sky130_fd_sc_hd__mux2_1 _17410_ (.A0(net447),
    .A1(\jtag.instructionRegister.data[1] ),
    .S(net1779),
    .X(_03510_));
 sky130_fd_sc_hd__o211a_1 _17411_ (.A1(_03504_),
    .A2(_03510_),
    .B1(_03509_),
    .C1(net1886),
    .X(_01168_));
 sky130_fd_sc_hd__a31o_1 _17412_ (.A1(net1782),
    .A2(net1777),
    .A3(_08620_),
    .B1(\jtag.instructionRegister.data[3] ),
    .X(_03511_));
 sky130_fd_sc_hd__mux2_1 _17413_ (.A0(net448),
    .A1(\jtag.instructionRegister.data[2] ),
    .S(net1779),
    .X(_03512_));
 sky130_fd_sc_hd__o211a_1 _17414_ (.A1(_03504_),
    .A2(_03512_),
    .B1(_03511_),
    .C1(net1886),
    .X(_01169_));
 sky130_fd_sc_hd__a31o_1 _17415_ (.A1(net1781),
    .A2(net1778),
    .A3(_08620_),
    .B1(\jtag.instructionRegister.data[4] ),
    .X(_03513_));
 sky130_fd_sc_hd__mux2_1 _17416_ (.A0(net449),
    .A1(\jtag.instructionRegister.data[3] ),
    .S(net1779),
    .X(_03514_));
 sky130_fd_sc_hd__o211a_1 _17417_ (.A1(_03504_),
    .A2(_03514_),
    .B1(_03513_),
    .C1(net1886),
    .X(_01170_));
 sky130_fd_sc_hd__o21ai_1 _17418_ (.A1(_04398_),
    .A2(net187),
    .B1(\jtag.tckState ),
    .Y(_03515_));
 sky130_fd_sc_hd__o211a_1 _17419_ (.A1(net187),
    .A2(\jtag.tckState ),
    .B1(net1890),
    .C1(_03515_),
    .X(_01171_));
 sky130_fd_sc_hd__and2_1 _17420_ (.A(net187),
    .B(net1890),
    .X(_01172_));
 sky130_fd_sc_hd__nor2_1 _17421_ (.A(_08632_),
    .B(_03395_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand2_2 _17422_ (.A(\jtag.state[3] ),
    .B(\jtag.state[2] ),
    .Y(_03517_));
 sky130_fd_sc_hd__and4_1 _17423_ (.A(\jtag.state[3] ),
    .B(\jtag.state[2] ),
    .C(net1777),
    .D(net1780),
    .X(_03518_));
 sky130_fd_sc_hd__o21a_4 _17424_ (.A1(_03516_),
    .A2(_03518_),
    .B1(net1782),
    .X(_03519_));
 sky130_fd_sc_hd__mux2_1 _17425_ (.A0(net445),
    .A1(\jtag.instructionRegister.data[0] ),
    .S(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__and2_1 _17426_ (.A(net1890),
    .B(_03520_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _17427_ (.A0(net446),
    .A1(\jtag.instructionRegister.data[1] ),
    .S(_03519_),
    .X(_03521_));
 sky130_fd_sc_hd__and2_1 _17428_ (.A(net1890),
    .B(_03521_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _17429_ (.A0(net447),
    .A1(\jtag.instructionRegister.data[2] ),
    .S(_03519_),
    .X(_03522_));
 sky130_fd_sc_hd__or2_1 _17430_ (.A(net1961),
    .B(_03522_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _17431_ (.A0(net448),
    .A1(\jtag.instructionRegister.data[3] ),
    .S(_03519_),
    .X(_03523_));
 sky130_fd_sc_hd__and2_1 _17432_ (.A(net1890),
    .B(_03523_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _17433_ (.A0(net449),
    .A1(\jtag.instructionRegister.data[4] ),
    .S(_03519_),
    .X(_03524_));
 sky130_fd_sc_hd__and2_1 _17434_ (.A(net1886),
    .B(_03524_),
    .X(_01177_));
 sky130_fd_sc_hd__o21ai_1 _17435_ (.A1(net1779),
    .A2(_08633_),
    .B1(net1342),
    .Y(_03525_));
 sky130_fd_sc_hd__nor2_1 _17436_ (.A(net1777),
    .B(_04399_),
    .Y(_03526_));
 sky130_fd_sc_hd__a211o_1 _17437_ (.A1(_03394_),
    .A2(_03526_),
    .B1(_03518_),
    .C1(_09060_),
    .X(_03527_));
 sky130_fd_sc_hd__or2_1 _17438_ (.A(net189),
    .B(_08621_),
    .X(_03528_));
 sky130_fd_sc_hd__a31o_1 _17439_ (.A1(\jtag.state[3] ),
    .A2(\jtag.state[2] ),
    .A3(_03526_),
    .B1(_03516_),
    .X(_03529_));
 sky130_fd_sc_hd__o32a_1 _17440_ (.A1(_03527_),
    .A2(_03528_),
    .A3(_03529_),
    .B1(_03525_),
    .B2(_04443_),
    .X(_03530_));
 sky130_fd_sc_hd__and3_1 _17441_ (.A(net1778),
    .B(_04399_),
    .C(_03394_),
    .X(_03531_));
 sky130_fd_sc_hd__nor2_1 _17442_ (.A(net1779),
    .B(_03517_),
    .Y(_03532_));
 sky130_fd_sc_hd__or4_1 _17443_ (.A(_04398_),
    .B(_03530_),
    .C(_03531_),
    .D(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__o211a_1 _17444_ (.A1(net1781),
    .A2(net1779),
    .B1(net1886),
    .C1(_03533_),
    .X(_01178_));
 sky130_fd_sc_hd__a31o_1 _17445_ (.A1(_03395_),
    .A2(_03517_),
    .A3(_03526_),
    .B1(_03528_),
    .X(_03534_));
 sky130_fd_sc_hd__nor2_1 _17446_ (.A(net1777),
    .B(_03517_),
    .Y(_03535_));
 sky130_fd_sc_hd__o32a_1 _17447_ (.A1(_04443_),
    .A2(_03527_),
    .A3(_03535_),
    .B1(_03534_),
    .B2(_03531_),
    .X(_03536_));
 sky130_fd_sc_hd__a31o_1 _17448_ (.A1(\jtag.state[2] ),
    .A2(net1777),
    .A3(_04399_),
    .B1(_04398_),
    .X(_03537_));
 sky130_fd_sc_hd__o221a_1 _17449_ (.A1(net1782),
    .A2(net1777),
    .B1(_03536_),
    .B2(_03537_),
    .C1(net1886),
    .X(_01179_));
 sky130_fd_sc_hd__o211a_1 _17450_ (.A1(_08620_),
    .A2(_03532_),
    .B1(net1777),
    .C1(net189),
    .X(_03538_));
 sky130_fd_sc_hd__or2_1 _17451_ (.A(_04399_),
    .B(_08633_),
    .X(_03539_));
 sky130_fd_sc_hd__nor2_1 _17452_ (.A(net189),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__o21ai_1 _17453_ (.A1(net1777),
    .A2(_03517_),
    .B1(net1782),
    .Y(_03541_));
 sky130_fd_sc_hd__or4_1 _17454_ (.A(_03525_),
    .B(_03538_),
    .C(_03540_),
    .D(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__o211a_1 _17455_ (.A1(net1782),
    .A2(\jtag.state[2] ),
    .B1(net1888),
    .C1(_03542_),
    .X(_01180_));
 sky130_fd_sc_hd__nand2b_1 _17456_ (.A_N(_03531_),
    .B(_03539_),
    .Y(_03543_));
 sky130_fd_sc_hd__and3_1 _17457_ (.A(_04443_),
    .B(_08620_),
    .C(_03526_),
    .X(_03544_));
 sky130_fd_sc_hd__a211o_1 _17458_ (.A1(net1777),
    .A2(_03532_),
    .B1(_03541_),
    .C1(_08621_),
    .X(_03545_));
 sky130_fd_sc_hd__a211o_1 _17459_ (.A1(net189),
    .A2(_03543_),
    .B1(_03544_),
    .C1(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__o211a_1 _17460_ (.A1(\jtag.state[3] ),
    .A2(net1782),
    .B1(net1888),
    .C1(_03546_),
    .X(_01181_));
 sky130_fd_sc_hd__or2_4 _17461_ (.A(_07835_),
    .B(_03367_),
    .X(_03547_));
 sky130_fd_sc_hd__nand2_1 _17462_ (.A(\jtag.managementReadData[0] ),
    .B(net1642),
    .Y(_03548_));
 sky130_fd_sc_hd__a21oi_1 _17463_ (.A1(net804),
    .A2(_03548_),
    .B1(net1980),
    .Y(_01182_));
 sky130_fd_sc_hd__nand2_1 _17464_ (.A(\jtag.managementReadData[1] ),
    .B(net1643),
    .Y(_03549_));
 sky130_fd_sc_hd__a21oi_1 _17465_ (.A1(net805),
    .A2(_03549_),
    .B1(net1982),
    .Y(_01183_));
 sky130_fd_sc_hd__nand2_1 _17466_ (.A(\jtag.managementReadData[2] ),
    .B(net1642),
    .Y(_03550_));
 sky130_fd_sc_hd__a21oi_1 _17467_ (.A1(net804),
    .A2(_03550_),
    .B1(net1985),
    .Y(_01184_));
 sky130_fd_sc_hd__nand2_1 _17468_ (.A(\jtag.managementReadData[3] ),
    .B(net1643),
    .Y(_03551_));
 sky130_fd_sc_hd__a21oi_1 _17469_ (.A1(net805),
    .A2(_03551_),
    .B1(net1987),
    .Y(_01185_));
 sky130_fd_sc_hd__nand2_1 _17470_ (.A(\jtag.managementReadData[4] ),
    .B(net1643),
    .Y(_03552_));
 sky130_fd_sc_hd__a21oi_1 _17471_ (.A1(net805),
    .A2(_03552_),
    .B1(net1996),
    .Y(_01186_));
 sky130_fd_sc_hd__nand2_1 _17472_ (.A(\jtag.managementReadData[5] ),
    .B(net1642),
    .Y(_03553_));
 sky130_fd_sc_hd__a21oi_1 _17473_ (.A1(net804),
    .A2(_03553_),
    .B1(net1996),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_1 _17474_ (.A(\jtag.managementReadData[6] ),
    .B(net1642),
    .Y(_03554_));
 sky130_fd_sc_hd__a21oi_1 _17475_ (.A1(net804),
    .A2(_03554_),
    .B1(net1990),
    .Y(_01188_));
 sky130_fd_sc_hd__nand2_1 _17476_ (.A(\jtag.managementReadData[7] ),
    .B(net1642),
    .Y(_03555_));
 sky130_fd_sc_hd__a21oi_1 _17477_ (.A1(net804),
    .A2(_03555_),
    .B1(net1990),
    .Y(_01189_));
 sky130_fd_sc_hd__nand2_1 _17478_ (.A(\jtag.managementReadData[8] ),
    .B(net1642),
    .Y(_03556_));
 sky130_fd_sc_hd__a21oi_1 _17479_ (.A1(net804),
    .A2(_03556_),
    .B1(net1990),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _17480_ (.A(\jtag.managementReadData[9] ),
    .B(net1642),
    .Y(_03557_));
 sky130_fd_sc_hd__a21oi_1 _17481_ (.A1(net804),
    .A2(_03557_),
    .B1(net1996),
    .Y(_01191_));
 sky130_fd_sc_hd__nand2_1 _17482_ (.A(\jtag.managementReadData[10] ),
    .B(net1642),
    .Y(_03558_));
 sky130_fd_sc_hd__a21oi_1 _17483_ (.A1(net804),
    .A2(_03558_),
    .B1(net1996),
    .Y(_01192_));
 sky130_fd_sc_hd__nand2_1 _17484_ (.A(\jtag.managementReadData[11] ),
    .B(net1642),
    .Y(_03559_));
 sky130_fd_sc_hd__a21oi_1 _17485_ (.A1(net804),
    .A2(_03559_),
    .B1(net1995),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_1 _17486_ (.A(\jtag.managementReadData[12] ),
    .B(net1642),
    .Y(_03560_));
 sky130_fd_sc_hd__a21oi_1 _17487_ (.A1(net804),
    .A2(_03560_),
    .B1(net1985),
    .Y(_01194_));
 sky130_fd_sc_hd__nand2_1 _17488_ (.A(\jtag.managementReadData[13] ),
    .B(net1643),
    .Y(_03561_));
 sky130_fd_sc_hd__a21oi_1 _17489_ (.A1(net805),
    .A2(_03561_),
    .B1(net1981),
    .Y(_01195_));
 sky130_fd_sc_hd__nand2_1 _17490_ (.A(\jtag.managementReadData[14] ),
    .B(net1643),
    .Y(_03562_));
 sky130_fd_sc_hd__a21oi_1 _17491_ (.A1(net805),
    .A2(_03562_),
    .B1(net1977),
    .Y(_01196_));
 sky130_fd_sc_hd__nand2_1 _17492_ (.A(\jtag.managementReadData[15] ),
    .B(net1643),
    .Y(_03563_));
 sky130_fd_sc_hd__a21oi_1 _17493_ (.A1(net805),
    .A2(_03563_),
    .B1(net1976),
    .Y(_01197_));
 sky130_fd_sc_hd__nand2_1 _17494_ (.A(\jtag.managementReadData[16] ),
    .B(net1643),
    .Y(_03564_));
 sky130_fd_sc_hd__a21oi_1 _17495_ (.A1(net805),
    .A2(_03564_),
    .B1(net1976),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_1 _17496_ (.A(\jtag.managementReadData[17] ),
    .B(net1641),
    .Y(_03565_));
 sky130_fd_sc_hd__a21oi_1 _17497_ (.A1(net803),
    .A2(_03565_),
    .B1(net1972),
    .Y(_01199_));
 sky130_fd_sc_hd__nand2_1 _17498_ (.A(\jtag.managementReadData[18] ),
    .B(net1641),
    .Y(_03566_));
 sky130_fd_sc_hd__a21oi_1 _17499_ (.A1(net803),
    .A2(_03566_),
    .B1(net1972),
    .Y(_01200_));
 sky130_fd_sc_hd__nand2_1 _17500_ (.A(\jtag.managementReadData[19] ),
    .B(net1641),
    .Y(_03567_));
 sky130_fd_sc_hd__a21oi_1 _17501_ (.A1(net803),
    .A2(_03567_),
    .B1(net1967),
    .Y(_01201_));
 sky130_fd_sc_hd__nand2_1 _17502_ (.A(\jtag.managementReadData[20] ),
    .B(net1641),
    .Y(_03568_));
 sky130_fd_sc_hd__a21oi_1 _17503_ (.A1(net803),
    .A2(_03568_),
    .B1(net1966),
    .Y(_01202_));
 sky130_fd_sc_hd__nand2_1 _17504_ (.A(\jtag.managementReadData[21] ),
    .B(net1640),
    .Y(_03569_));
 sky130_fd_sc_hd__a21oi_1 _17505_ (.A1(net803),
    .A2(_03569_),
    .B1(net1962),
    .Y(_01203_));
 sky130_fd_sc_hd__nand2_1 _17506_ (.A(\jtag.managementReadData[22] ),
    .B(net1639),
    .Y(_03570_));
 sky130_fd_sc_hd__a21oi_1 _17507_ (.A1(net802),
    .A2(_03570_),
    .B1(net1962),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_1 _17508_ (.A(\jtag.managementReadData[23] ),
    .B(net1640),
    .Y(_03571_));
 sky130_fd_sc_hd__a21oi_1 _17509_ (.A1(net802),
    .A2(_03571_),
    .B1(net1962),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_1 _17510_ (.A(\jtag.managementReadData[24] ),
    .B(net1640),
    .Y(_03572_));
 sky130_fd_sc_hd__a21oi_1 _17511_ (.A1(net802),
    .A2(_03572_),
    .B1(net1961),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_1 _17512_ (.A(\jtag.managementReadData[25] ),
    .B(net1639),
    .Y(_03573_));
 sky130_fd_sc_hd__a21oi_1 _17513_ (.A1(net802),
    .A2(_03573_),
    .B1(net1961),
    .Y(_01207_));
 sky130_fd_sc_hd__nand2_1 _17514_ (.A(\jtag.managementReadData[26] ),
    .B(net1639),
    .Y(_03574_));
 sky130_fd_sc_hd__a21oi_1 _17515_ (.A1(net802),
    .A2(_03574_),
    .B1(net1961),
    .Y(_01208_));
 sky130_fd_sc_hd__nand2_1 _17516_ (.A(\jtag.managementReadData[27] ),
    .B(net1639),
    .Y(_03575_));
 sky130_fd_sc_hd__a21oi_1 _17517_ (.A1(net802),
    .A2(_03575_),
    .B1(net1961),
    .Y(_01209_));
 sky130_fd_sc_hd__nand2_1 _17518_ (.A(\jtag.managementReadData[28] ),
    .B(net1639),
    .Y(_03576_));
 sky130_fd_sc_hd__a21oi_1 _17519_ (.A1(net802),
    .A2(_03576_),
    .B1(net1961),
    .Y(_01210_));
 sky130_fd_sc_hd__nand2_1 _17520_ (.A(\jtag.managementReadData[29] ),
    .B(net1639),
    .Y(_03577_));
 sky130_fd_sc_hd__a21oi_1 _17521_ (.A1(net802),
    .A2(_03577_),
    .B1(net1961),
    .Y(_01211_));
 sky130_fd_sc_hd__nand2_1 _17522_ (.A(\jtag.managementReadData[30] ),
    .B(net1639),
    .Y(_03578_));
 sky130_fd_sc_hd__a21oi_1 _17523_ (.A1(net802),
    .A2(_03578_),
    .B1(net1961),
    .Y(_01212_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(\jtag.managementReadData[31] ),
    .B(net1640),
    .Y(_03579_));
 sky130_fd_sc_hd__a21oi_1 _17525_ (.A1(net802),
    .A2(_03579_),
    .B1(net1961),
    .Y(_01213_));
 sky130_fd_sc_hd__or4b_2 _17526_ (.A(\jtag.managementState[2] ),
    .B(_09062_),
    .C(_04397_),
    .D_N(\jtag.managementState[1] ),
    .X(_03580_));
 sky130_fd_sc_hd__nor2_1 _17527_ (.A(\jtag.dataBSRRegister.data[31] ),
    .B(\jtag.dataBSRRegister.data[30] ),
    .Y(_03581_));
 sky130_fd_sc_hd__or3_1 _17528_ (.A(\jtag.managementState[1] ),
    .B(_09063_),
    .C(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__or3b_1 _17529_ (.A(\jtag.managementState[2] ),
    .B(\jtag.managementState[0] ),
    .C_N(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__a21o_1 _17530_ (.A1(\jtag.managementState[1] ),
    .A2(net1242),
    .B1(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__o21a_1 _17531_ (.A1(net1218),
    .A2(_03581_),
    .B1(_03580_),
    .X(_03585_));
 sky130_fd_sc_hd__nor2_1 _17532_ (.A(net1969),
    .B(_03585_),
    .Y(_01214_));
 sky130_fd_sc_hd__a21o_1 _17533_ (.A1(_04397_),
    .A2(\jtag.dataBSRRegister.data[31] ),
    .B1(net1639),
    .X(_03586_));
 sky130_fd_sc_hd__a31o_1 _17534_ (.A1(_03580_),
    .A2(_03584_),
    .A3(_03586_),
    .B1(net1969),
    .X(_03587_));
 sky130_fd_sc_hd__o21ba_1 _17535_ (.A1(\jtag.managementState[1] ),
    .A2(_03583_),
    .B1_N(_03587_),
    .X(_01215_));
 sky130_fd_sc_hd__and4b_1 _17536_ (.A_N(\jtag.managementState[2] ),
    .B(\jtag.managementState[1] ),
    .C(\jtag.managementState[0] ),
    .D(net1887),
    .X(_03588_));
 sky130_fd_sc_hd__and3_1 _17537_ (.A(_03580_),
    .B(_03584_),
    .C(_03588_),
    .X(_01216_));
 sky130_fd_sc_hd__or3_2 _17538_ (.A(\core.csr.currentInstruction[11] ),
    .B(\core.csr.currentInstruction[9] ),
    .C(_04514_),
    .X(_03589_));
 sky130_fd_sc_hd__nor2_1 _17539_ (.A(_03040_),
    .B(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__and3_4 _17540_ (.A(net675),
    .B(net1072),
    .C(_03590_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_1 _17541_ (.A0(\core.registers[9][0] ),
    .A1(net1035),
    .S(net535),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _17542_ (.A0(\core.registers[9][1] ),
    .A1(net1039),
    .S(net534),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _17543_ (.A0(\core.registers[9][2] ),
    .A1(net1044),
    .S(net534),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _17544_ (.A0(\core.registers[9][3] ),
    .A1(net1050),
    .S(net534),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _17545_ (.A0(\core.registers[9][4] ),
    .A1(net1054),
    .S(net535),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _17546_ (.A0(\core.registers[9][5] ),
    .A1(net1058),
    .S(net534),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _17547_ (.A0(\core.registers[9][6] ),
    .A1(net1061),
    .S(net534),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _17548_ (.A0(\core.registers[9][7] ),
    .A1(net1132),
    .S(net534),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _17549_ (.A0(\core.registers[9][8] ),
    .A1(net957),
    .S(net534),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _17550_ (.A0(\core.registers[9][9] ),
    .A1(net963),
    .S(net533),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _17551_ (.A0(\core.registers[9][10] ),
    .A1(net967),
    .S(net535),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _17552_ (.A0(\core.registers[9][11] ),
    .A1(net970),
    .S(net533),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _17553_ (.A0(\core.registers[9][12] ),
    .A1(net987),
    .S(net535),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _17554_ (.A0(\core.registers[9][13] ),
    .A1(net983),
    .S(net535),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _17555_ (.A0(\core.registers[9][14] ),
    .A1(net977),
    .S(net535),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _17556_ (.A0(\core.registers[9][15] ),
    .A1(net979),
    .S(net534),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _17557_ (.A0(\core.registers[9][16] ),
    .A1(net1125),
    .S(net532),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _17558_ (.A0(\core.registers[9][17] ),
    .A1(net1129),
    .S(net532),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _17559_ (.A0(\core.registers[9][18] ),
    .A1(net1118),
    .S(net533),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _17560_ (.A0(\core.registers[9][19] ),
    .A1(net1120),
    .S(net532),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _17561_ (.A0(\core.registers[9][20] ),
    .A1(net1136),
    .S(net532),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _17562_ (.A0(\core.registers[9][21] ),
    .A1(net1140),
    .S(net532),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _17563_ (.A0(\core.registers[9][22] ),
    .A1(net1145),
    .S(net533),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _17564_ (.A0(\core.registers[9][23] ),
    .A1(net1150),
    .S(net532),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _17565_ (.A0(\core.registers[9][24] ),
    .A1(net1113),
    .S(net532),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _17566_ (.A0(\core.registers[9][25] ),
    .A1(net1110),
    .S(net532),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _17567_ (.A0(\core.registers[9][26] ),
    .A1(net1100),
    .S(net533),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _17568_ (.A0(\core.registers[9][27] ),
    .A1(net1105),
    .S(net532),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _17569_ (.A0(\core.registers[9][28] ),
    .A1(net1097),
    .S(net532),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _17570_ (.A0(\core.registers[9][29] ),
    .A1(net1094),
    .S(net535),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _17571_ (.A0(\core.registers[9][30] ),
    .A1(net1084),
    .S(net534),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _17572_ (.A0(\core.registers[9][31] ),
    .A1(net1088),
    .S(net534),
    .X(_01248_));
 sky130_fd_sc_hd__nor2_1 _17573_ (.A(_04516_),
    .B(_03040_),
    .Y(_03592_));
 sky130_fd_sc_hd__and3_4 _17574_ (.A(net679),
    .B(net1075),
    .C(_03592_),
    .X(_03593_));
 sky130_fd_sc_hd__mux2_1 _17575_ (.A0(\core.registers[1][0] ),
    .A1(net1038),
    .S(net530),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _17576_ (.A0(\core.registers[1][1] ),
    .A1(net1042),
    .S(net531),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _17577_ (.A0(\core.registers[1][2] ),
    .A1(net1045),
    .S(net530),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _17578_ (.A0(\core.registers[1][3] ),
    .A1(net1049),
    .S(net530),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _17579_ (.A0(\core.registers[1][4] ),
    .A1(net1053),
    .S(net530),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _17580_ (.A0(\core.registers[1][5] ),
    .A1(net1058),
    .S(net530),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _17581_ (.A0(\core.registers[1][6] ),
    .A1(net1063),
    .S(net531),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _17582_ (.A0(\core.registers[1][7] ),
    .A1(net1135),
    .S(net531),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _17583_ (.A0(\core.registers[1][8] ),
    .A1(net959),
    .S(net530),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _17584_ (.A0(\core.registers[1][9] ),
    .A1(net965),
    .S(net529),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _17585_ (.A0(\core.registers[1][10] ),
    .A1(net969),
    .S(net530),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _17586_ (.A0(\core.registers[1][11] ),
    .A1(net2011),
    .S(net529),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _17587_ (.A0(\core.registers[1][12] ),
    .A1(net990),
    .S(net529),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _17588_ (.A0(\core.registers[1][13] ),
    .A1(net985),
    .S(net530),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _17589_ (.A0(\core.registers[1][14] ),
    .A1(net978),
    .S(net530),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _17590_ (.A0(\core.registers[1][15] ),
    .A1(net982),
    .S(net530),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _17591_ (.A0(\core.registers[1][16] ),
    .A1(net1126),
    .S(net528),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _17592_ (.A0(\core.registers[1][17] ),
    .A1(net1130),
    .S(net528),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _17593_ (.A0(\core.registers[1][18] ),
    .A1(net1119),
    .S(net529),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _17594_ (.A0(\core.registers[1][19] ),
    .A1(net1122),
    .S(net528),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _17595_ (.A0(\core.registers[1][20] ),
    .A1(net1139),
    .S(net528),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _17596_ (.A0(\core.registers[1][21] ),
    .A1(net1142),
    .S(net528),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _17597_ (.A0(\core.registers[1][22] ),
    .A1(_04703_),
    .S(net529),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _17598_ (.A0(\core.registers[1][23] ),
    .A1(net1152),
    .S(net528),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _17599_ (.A0(\core.registers[1][24] ),
    .A1(net1114),
    .S(net528),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _17600_ (.A0(\core.registers[1][25] ),
    .A1(net1109),
    .S(net528),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _17601_ (.A0(\core.registers[1][26] ),
    .A1(net1103),
    .S(net529),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _17602_ (.A0(\core.registers[1][27] ),
    .A1(net1107),
    .S(net528),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _17603_ (.A0(\core.registers[1][28] ),
    .A1(net1099),
    .S(net528),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _17604_ (.A0(\core.registers[1][29] ),
    .A1(net1093),
    .S(net531),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _17605_ (.A0(\core.registers[1][30] ),
    .A1(net1087),
    .S(net531),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _17606_ (.A0(\core.registers[1][31] ),
    .A1(net1090),
    .S(net531),
    .X(_01280_));
 sky130_fd_sc_hd__nor2_1 _17607_ (.A(_09097_),
    .B(_03589_),
    .Y(_03594_));
 sky130_fd_sc_hd__and3_4 _17608_ (.A(net675),
    .B(net1072),
    .C(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__mux2_1 _17609_ (.A0(\core.registers[10][0] ),
    .A1(net1035),
    .S(net527),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _17610_ (.A0(\core.registers[10][1] ),
    .A1(net1039),
    .S(net526),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _17611_ (.A0(\core.registers[10][2] ),
    .A1(net1043),
    .S(net526),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _17612_ (.A0(\core.registers[10][3] ),
    .A1(net1050),
    .S(net526),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _17613_ (.A0(\core.registers[10][4] ),
    .A1(net1055),
    .S(net527),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _17614_ (.A0(\core.registers[10][5] ),
    .A1(net1057),
    .S(net526),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _17615_ (.A0(\core.registers[10][6] ),
    .A1(net1062),
    .S(net527),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _17616_ (.A0(\core.registers[10][7] ),
    .A1(net1132),
    .S(net526),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _17617_ (.A0(\core.registers[10][8] ),
    .A1(net957),
    .S(net526),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _17618_ (.A0(\core.registers[10][9] ),
    .A1(net963),
    .S(net525),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _17619_ (.A0(\core.registers[10][10] ),
    .A1(net967),
    .S(net527),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _17620_ (.A0(\core.registers[10][11] ),
    .A1(net970),
    .S(net525),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _17621_ (.A0(\core.registers[10][12] ),
    .A1(net987),
    .S(net525),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _17622_ (.A0(\core.registers[10][13] ),
    .A1(net983),
    .S(net527),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _17623_ (.A0(\core.registers[10][14] ),
    .A1(net976),
    .S(net527),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _17624_ (.A0(\core.registers[10][15] ),
    .A1(net979),
    .S(net526),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _17625_ (.A0(\core.registers[10][16] ),
    .A1(net1125),
    .S(net524),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _17626_ (.A0(\core.registers[10][17] ),
    .A1(net1129),
    .S(net524),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _17627_ (.A0(\core.registers[10][18] ),
    .A1(net1116),
    .S(net525),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _17628_ (.A0(\core.registers[10][19] ),
    .A1(net1120),
    .S(net524),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _17629_ (.A0(\core.registers[10][20] ),
    .A1(net1136),
    .S(net524),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _17630_ (.A0(\core.registers[10][21] ),
    .A1(net1141),
    .S(net524),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _17631_ (.A0(\core.registers[10][22] ),
    .A1(net1145),
    .S(net525),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _17632_ (.A0(\core.registers[10][23] ),
    .A1(net1149),
    .S(net524),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _17633_ (.A0(\core.registers[10][24] ),
    .A1(net1112),
    .S(net524),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _17634_ (.A0(\core.registers[10][25] ),
    .A1(net1110),
    .S(net524),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _17635_ (.A0(\core.registers[10][26] ),
    .A1(net1101),
    .S(net525),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _17636_ (.A0(\core.registers[10][27] ),
    .A1(net1104),
    .S(net524),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _17637_ (.A0(\core.registers[10][28] ),
    .A1(net1097),
    .S(net524),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _17638_ (.A0(\core.registers[10][29] ),
    .A1(net1094),
    .S(net526),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _17639_ (.A0(\core.registers[10][30] ),
    .A1(net1084),
    .S(net526),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _17640_ (.A0(\core.registers[10][31] ),
    .A1(net1088),
    .S(net526),
    .X(_01312_));
 sky130_fd_sc_hd__nor2_1 _17641_ (.A(_09093_),
    .B(_03589_),
    .Y(_03596_));
 sky130_fd_sc_hd__and3_4 _17642_ (.A(net675),
    .B(net1072),
    .C(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__mux2_1 _17643_ (.A0(\core.registers[11][0] ),
    .A1(net1035),
    .S(net523),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _17644_ (.A0(\core.registers[11][1] ),
    .A1(net1039),
    .S(net522),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _17645_ (.A0(\core.registers[11][2] ),
    .A1(net1043),
    .S(net522),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _17646_ (.A0(\core.registers[11][3] ),
    .A1(net1050),
    .S(net522),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _17647_ (.A0(\core.registers[11][4] ),
    .A1(net1055),
    .S(net523),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _17648_ (.A0(\core.registers[11][5] ),
    .A1(net1058),
    .S(net522),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _17649_ (.A0(\core.registers[11][6] ),
    .A1(net1062),
    .S(net523),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _17650_ (.A0(\core.registers[11][7] ),
    .A1(net1132),
    .S(net522),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _17651_ (.A0(\core.registers[11][8] ),
    .A1(net957),
    .S(net522),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _17652_ (.A0(\core.registers[11][9] ),
    .A1(net963),
    .S(net521),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _17653_ (.A0(\core.registers[11][10] ),
    .A1(net967),
    .S(net523),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _17654_ (.A0(\core.registers[11][11] ),
    .A1(net970),
    .S(net521),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _17655_ (.A0(\core.registers[11][12] ),
    .A1(net988),
    .S(net521),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _17656_ (.A0(\core.registers[11][13] ),
    .A1(net983),
    .S(net523),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _17657_ (.A0(\core.registers[11][14] ),
    .A1(net976),
    .S(net523),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _17658_ (.A0(\core.registers[11][15] ),
    .A1(net979),
    .S(net522),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _17659_ (.A0(\core.registers[11][16] ),
    .A1(net1125),
    .S(net520),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _17660_ (.A0(\core.registers[11][17] ),
    .A1(net1129),
    .S(net520),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _17661_ (.A0(\core.registers[11][18] ),
    .A1(net1116),
    .S(net521),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _17662_ (.A0(\core.registers[11][19] ),
    .A1(net1120),
    .S(net520),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _17663_ (.A0(\core.registers[11][20] ),
    .A1(net1136),
    .S(net520),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _17664_ (.A0(\core.registers[11][21] ),
    .A1(net1141),
    .S(net520),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _17665_ (.A0(\core.registers[11][22] ),
    .A1(net1145),
    .S(net521),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _17666_ (.A0(\core.registers[11][23] ),
    .A1(net1149),
    .S(net520),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _17667_ (.A0(\core.registers[11][24] ),
    .A1(net1112),
    .S(net520),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _17668_ (.A0(\core.registers[11][25] ),
    .A1(net1110),
    .S(net520),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _17669_ (.A0(\core.registers[11][26] ),
    .A1(net1100),
    .S(net521),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _17670_ (.A0(\core.registers[11][27] ),
    .A1(net1104),
    .S(net520),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _17671_ (.A0(\core.registers[11][28] ),
    .A1(net1096),
    .S(net520),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _17672_ (.A0(\core.registers[11][29] ),
    .A1(net1094),
    .S(net522),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _17673_ (.A0(\core.registers[11][30] ),
    .A1(net1084),
    .S(net522),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _17674_ (.A0(\core.registers[11][31] ),
    .A1(net1089),
    .S(net522),
    .X(_01376_));
 sky130_fd_sc_hd__nor2_1 _17675_ (.A(_04512_),
    .B(_03589_),
    .Y(_03598_));
 sky130_fd_sc_hd__and3_4 _17676_ (.A(net675),
    .B(net1072),
    .C(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__mux2_1 _17677_ (.A0(\core.registers[8][0] ),
    .A1(net1035),
    .S(net519),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _17678_ (.A0(\core.registers[8][1] ),
    .A1(net1039),
    .S(net518),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _17679_ (.A0(\core.registers[8][2] ),
    .A1(net1044),
    .S(net518),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _17680_ (.A0(\core.registers[8][3] ),
    .A1(net1050),
    .S(net518),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _17681_ (.A0(\core.registers[8][4] ),
    .A1(net1054),
    .S(net519),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _17682_ (.A0(\core.registers[8][5] ),
    .A1(net1058),
    .S(net518),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _17683_ (.A0(\core.registers[8][6] ),
    .A1(net1061),
    .S(net518),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _17684_ (.A0(\core.registers[8][7] ),
    .A1(net1132),
    .S(net518),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _17685_ (.A0(\core.registers[8][8] ),
    .A1(net957),
    .S(net518),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _17686_ (.A0(\core.registers[8][9] ),
    .A1(net963),
    .S(net517),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _17687_ (.A0(\core.registers[8][10] ),
    .A1(net967),
    .S(net519),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _17688_ (.A0(\core.registers[8][11] ),
    .A1(net970),
    .S(net517),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _17689_ (.A0(\core.registers[8][12] ),
    .A1(net987),
    .S(net519),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _17690_ (.A0(\core.registers[8][13] ),
    .A1(net983),
    .S(net519),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _17691_ (.A0(\core.registers[8][14] ),
    .A1(net977),
    .S(net519),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _17692_ (.A0(\core.registers[8][15] ),
    .A1(net980),
    .S(net518),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _17693_ (.A0(\core.registers[8][16] ),
    .A1(net1125),
    .S(net516),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _17694_ (.A0(\core.registers[8][17] ),
    .A1(net1129),
    .S(net516),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _17695_ (.A0(\core.registers[8][18] ),
    .A1(net1116),
    .S(net517),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _17696_ (.A0(\core.registers[8][19] ),
    .A1(net1120),
    .S(net516),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _17697_ (.A0(\core.registers[8][20] ),
    .A1(net1136),
    .S(net516),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _17698_ (.A0(\core.registers[8][21] ),
    .A1(net1140),
    .S(net516),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _17699_ (.A0(\core.registers[8][22] ),
    .A1(net1145),
    .S(net517),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _17700_ (.A0(\core.registers[8][23] ),
    .A1(net1150),
    .S(net516),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _17701_ (.A0(\core.registers[8][24] ),
    .A1(net1113),
    .S(net516),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _17702_ (.A0(\core.registers[8][25] ),
    .A1(net1110),
    .S(net516),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _17703_ (.A0(\core.registers[8][26] ),
    .A1(net1100),
    .S(net517),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _17704_ (.A0(\core.registers[8][27] ),
    .A1(net1105),
    .S(net516),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _17705_ (.A0(\core.registers[8][28] ),
    .A1(net1096),
    .S(net516),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _17706_ (.A0(\core.registers[8][29] ),
    .A1(net1094),
    .S(net519),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _17707_ (.A0(\core.registers[8][30] ),
    .A1(net1084),
    .S(net518),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _17708_ (.A0(\core.registers[8][31] ),
    .A1(net1088),
    .S(net518),
    .X(_01408_));
 sky130_fd_sc_hd__or3_2 _17709_ (.A(\core.csr.currentInstruction[11] ),
    .B(\core.csr.currentInstruction[10] ),
    .C(_04515_),
    .X(_03600_));
 sky130_fd_sc_hd__nor2_1 _17710_ (.A(_09093_),
    .B(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__and3_4 _17711_ (.A(net675),
    .B(net1073),
    .C(_03601_),
    .X(_03602_));
 sky130_fd_sc_hd__mux2_1 _17712_ (.A0(\core.registers[7][0] ),
    .A1(net1038),
    .S(net514),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _17713_ (.A0(\core.registers[7][1] ),
    .A1(net1042),
    .S(net514),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _17714_ (.A0(\core.registers[7][2] ),
    .A1(net1045),
    .S(net515),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _17715_ (.A0(\core.registers[7][3] ),
    .A1(net1048),
    .S(net514),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _17716_ (.A0(\core.registers[7][4] ),
    .A1(net1054),
    .S(net514),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _17717_ (.A0(\core.registers[7][5] ),
    .A1(net1057),
    .S(net515),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _17718_ (.A0(\core.registers[7][6] ),
    .A1(net1063),
    .S(net515),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _17719_ (.A0(\core.registers[7][7] ),
    .A1(net1135),
    .S(net515),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _17720_ (.A0(\core.registers[7][8] ),
    .A1(net959),
    .S(net515),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _17721_ (.A0(\core.registers[7][9] ),
    .A1(net964),
    .S(net513),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _17722_ (.A0(\core.registers[7][10] ),
    .A1(net969),
    .S(net514),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _17723_ (.A0(\core.registers[7][11] ),
    .A1(net973),
    .S(net513),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _17724_ (.A0(\core.registers[7][12] ),
    .A1(net990),
    .S(net513),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _17725_ (.A0(\core.registers[7][13] ),
    .A1(net985),
    .S(net514),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _17726_ (.A0(\core.registers[7][14] ),
    .A1(net975),
    .S(net514),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _17727_ (.A0(\core.registers[7][15] ),
    .A1(net982),
    .S(net514),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _17728_ (.A0(\core.registers[7][16] ),
    .A1(net1126),
    .S(net512),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _17729_ (.A0(\core.registers[7][17] ),
    .A1(net1128),
    .S(net512),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _17730_ (.A0(\core.registers[7][18] ),
    .A1(net1118),
    .S(net513),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _17731_ (.A0(\core.registers[7][19] ),
    .A1(net1122),
    .S(net512),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _17732_ (.A0(\core.registers[7][20] ),
    .A1(net1139),
    .S(net512),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _17733_ (.A0(\core.registers[7][21] ),
    .A1(net1143),
    .S(net512),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _17734_ (.A0(\core.registers[7][22] ),
    .A1(net1148),
    .S(net513),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _17735_ (.A0(\core.registers[7][23] ),
    .A1(net1152),
    .S(net512),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _17736_ (.A0(\core.registers[7][24] ),
    .A1(net1114),
    .S(net512),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _17737_ (.A0(\core.registers[7][25] ),
    .A1(net1109),
    .S(net512),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _17738_ (.A0(\core.registers[7][26] ),
    .A1(net1103),
    .S(net513),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _17739_ (.A0(\core.registers[7][27] ),
    .A1(net1107),
    .S(net512),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _17740_ (.A0(\core.registers[7][28] ),
    .A1(net1097),
    .S(net512),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _17741_ (.A0(\core.registers[7][29] ),
    .A1(net1093),
    .S(net514),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _17742_ (.A0(\core.registers[7][30] ),
    .A1(net1087),
    .S(net515),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _17743_ (.A0(\core.registers[7][31] ),
    .A1(net1090),
    .S(net514),
    .X(_01440_));
 sky130_fd_sc_hd__nor2_1 _17744_ (.A(_09097_),
    .B(_03600_),
    .Y(_03603_));
 sky130_fd_sc_hd__and3_4 _17745_ (.A(net675),
    .B(net1073),
    .C(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__mux2_1 _17746_ (.A0(\core.registers[6][0] ),
    .A1(net1037),
    .S(net510),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _17747_ (.A0(\core.registers[6][1] ),
    .A1(net1042),
    .S(net510),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _17748_ (.A0(\core.registers[6][2] ),
    .A1(net1045),
    .S(net511),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _17749_ (.A0(\core.registers[6][3] ),
    .A1(net1049),
    .S(net510),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _17750_ (.A0(\core.registers[6][4] ),
    .A1(net1054),
    .S(net510),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _17751_ (.A0(\core.registers[6][5] ),
    .A1(net1057),
    .S(net511),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _17752_ (.A0(\core.registers[6][6] ),
    .A1(net1063),
    .S(net511),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _17753_ (.A0(\core.registers[6][7] ),
    .A1(net1135),
    .S(net511),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _17754_ (.A0(\core.registers[6][8] ),
    .A1(net959),
    .S(net511),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _17755_ (.A0(\core.registers[6][9] ),
    .A1(net964),
    .S(net509),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _17756_ (.A0(\core.registers[6][10] ),
    .A1(net969),
    .S(net510),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _17757_ (.A0(\core.registers[6][11] ),
    .A1(net973),
    .S(net509),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _17758_ (.A0(\core.registers[6][12] ),
    .A1(net990),
    .S(net509),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _17759_ (.A0(\core.registers[6][13] ),
    .A1(net985),
    .S(net510),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _17760_ (.A0(\core.registers[6][14] ),
    .A1(net975),
    .S(net510),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _17761_ (.A0(\core.registers[6][15] ),
    .A1(net982),
    .S(net510),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _17762_ (.A0(\core.registers[6][16] ),
    .A1(net1126),
    .S(net508),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _17763_ (.A0(\core.registers[6][17] ),
    .A1(net1128),
    .S(net508),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _17764_ (.A0(\core.registers[6][18] ),
    .A1(net1118),
    .S(net509),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _17765_ (.A0(\core.registers[6][19] ),
    .A1(net1122),
    .S(net508),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _17766_ (.A0(\core.registers[6][20] ),
    .A1(net1139),
    .S(net508),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _17767_ (.A0(\core.registers[6][21] ),
    .A1(net1142),
    .S(net508),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _17768_ (.A0(\core.registers[6][22] ),
    .A1(net1148),
    .S(net509),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _17769_ (.A0(\core.registers[6][23] ),
    .A1(net1152),
    .S(net508),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _17770_ (.A0(\core.registers[6][24] ),
    .A1(net1114),
    .S(net508),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _17771_ (.A0(\core.registers[6][25] ),
    .A1(net1109),
    .S(net508),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _17772_ (.A0(\core.registers[6][26] ),
    .A1(net1103),
    .S(net509),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _17773_ (.A0(\core.registers[6][27] ),
    .A1(net1107),
    .S(net508),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _17774_ (.A0(\core.registers[6][28] ),
    .A1(net1097),
    .S(net508),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _17775_ (.A0(\core.registers[6][29] ),
    .A1(net1093),
    .S(net510),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _17776_ (.A0(\core.registers[6][30] ),
    .A1(net1087),
    .S(net511),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _17777_ (.A0(\core.registers[6][31] ),
    .A1(net1090),
    .S(net510),
    .X(_01472_));
 sky130_fd_sc_hd__nor2_1 _17778_ (.A(_09098_),
    .B(_03040_),
    .Y(_03605_));
 sky130_fd_sc_hd__and3_4 _17779_ (.A(net679),
    .B(net1074),
    .C(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__mux2_1 _17780_ (.A0(\core.registers[29][0] ),
    .A1(net1035),
    .S(net506),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _17781_ (.A0(\core.registers[29][1] ),
    .A1(net1041),
    .S(net507),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _17782_ (.A0(\core.registers[29][2] ),
    .A1(net1047),
    .S(net507),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _17783_ (.A0(\core.registers[29][3] ),
    .A1(net1050),
    .S(net506),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _17784_ (.A0(\core.registers[29][4] ),
    .A1(net1056),
    .S(net507),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _17785_ (.A0(\core.registers[29][5] ),
    .A1(net1059),
    .S(net506),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _17786_ (.A0(\core.registers[29][6] ),
    .A1(net1064),
    .S(net506),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _17787_ (.A0(\core.registers[29][7] ),
    .A1(net1134),
    .S(net506),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _17788_ (.A0(\core.registers[29][8] ),
    .A1(net958),
    .S(net507),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _17789_ (.A0(\core.registers[29][9] ),
    .A1(net962),
    .S(net505),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _17790_ (.A0(\core.registers[29][10] ),
    .A1(net966),
    .S(net507),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _17791_ (.A0(\core.registers[29][11] ),
    .A1(net970),
    .S(net505),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _17792_ (.A0(\core.registers[29][12] ),
    .A1(net988),
    .S(net507),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _17793_ (.A0(\core.registers[29][13] ),
    .A1(net983),
    .S(net506),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _17794_ (.A0(\core.registers[29][14] ),
    .A1(net974),
    .S(net507),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _17795_ (.A0(\core.registers[29][15] ),
    .A1(net979),
    .S(net506),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _17796_ (.A0(\core.registers[29][16] ),
    .A1(net1127),
    .S(net504),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _17797_ (.A0(\core.registers[29][17] ),
    .A1(net1131),
    .S(net504),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _17798_ (.A0(\core.registers[29][18] ),
    .A1(net1117),
    .S(net505),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _17799_ (.A0(\core.registers[29][19] ),
    .A1(net1121),
    .S(net504),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _17800_ (.A0(\core.registers[29][20] ),
    .A1(net1136),
    .S(net504),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _17801_ (.A0(\core.registers[29][21] ),
    .A1(net1140),
    .S(net504),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _17802_ (.A0(\core.registers[29][22] ),
    .A1(net1145),
    .S(net505),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _17803_ (.A0(\core.registers[29][23] ),
    .A1(net1150),
    .S(net504),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _17804_ (.A0(\core.registers[29][24] ),
    .A1(net1112),
    .S(net504),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _17805_ (.A0(\core.registers[29][25] ),
    .A1(net1110),
    .S(net504),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _17806_ (.A0(\core.registers[29][26] ),
    .A1(net1100),
    .S(net505),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _17807_ (.A0(\core.registers[29][27] ),
    .A1(net1104),
    .S(net504),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _17808_ (.A0(\core.registers[29][28] ),
    .A1(net1099),
    .S(net504),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _17809_ (.A0(\core.registers[29][29] ),
    .A1(net1095),
    .S(net506),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _17810_ (.A0(\core.registers[29][30] ),
    .A1(net1086),
    .S(net506),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _17811_ (.A0(\core.registers[29][31] ),
    .A1(net1091),
    .S(net506),
    .X(_01504_));
 sky130_fd_sc_hd__nor2_1 _17812_ (.A(_03040_),
    .B(_03600_),
    .Y(_03607_));
 sky130_fd_sc_hd__and3_4 _17813_ (.A(net676),
    .B(net1073),
    .C(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__mux2_1 _17814_ (.A0(\core.registers[5][0] ),
    .A1(net1038),
    .S(net502),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _17815_ (.A0(\core.registers[5][1] ),
    .A1(net1042),
    .S(net502),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _17816_ (.A0(\core.registers[5][2] ),
    .A1(net1045),
    .S(net503),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _17817_ (.A0(\core.registers[5][3] ),
    .A1(net1049),
    .S(net502),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _17818_ (.A0(\core.registers[5][4] ),
    .A1(net1053),
    .S(net502),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _17819_ (.A0(\core.registers[5][5] ),
    .A1(net1058),
    .S(net503),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _17820_ (.A0(\core.registers[5][6] ),
    .A1(net1063),
    .S(net503),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _17821_ (.A0(\core.registers[5][7] ),
    .A1(net1135),
    .S(net503),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _17822_ (.A0(\core.registers[5][8] ),
    .A1(net959),
    .S(net503),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _17823_ (.A0(\core.registers[5][9] ),
    .A1(net964),
    .S(net501),
    .X(_01514_));
 sky130_fd_sc_hd__mux2_1 _17824_ (.A0(\core.registers[5][10] ),
    .A1(net969),
    .S(net502),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _17825_ (.A0(\core.registers[5][11] ),
    .A1(net2011),
    .S(net501),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _17826_ (.A0(\core.registers[5][12] ),
    .A1(net990),
    .S(net501),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _17827_ (.A0(\core.registers[5][13] ),
    .A1(net985),
    .S(net502),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _17828_ (.A0(\core.registers[5][14] ),
    .A1(net978),
    .S(net502),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _17829_ (.A0(\core.registers[5][15] ),
    .A1(net982),
    .S(net502),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _17830_ (.A0(\core.registers[5][16] ),
    .A1(net1126),
    .S(net500),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _17831_ (.A0(\core.registers[5][17] ),
    .A1(net1128),
    .S(net500),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _17832_ (.A0(\core.registers[5][18] ),
    .A1(net1118),
    .S(net501),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _17833_ (.A0(\core.registers[5][19] ),
    .A1(net1122),
    .S(net500),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _17834_ (.A0(\core.registers[5][20] ),
    .A1(net1139),
    .S(net500),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _17835_ (.A0(\core.registers[5][21] ),
    .A1(net1142),
    .S(net500),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _17836_ (.A0(\core.registers[5][22] ),
    .A1(net1147),
    .S(net501),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _17837_ (.A0(\core.registers[5][23] ),
    .A1(net1152),
    .S(net500),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _17838_ (.A0(\core.registers[5][24] ),
    .A1(net1114),
    .S(net500),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _17839_ (.A0(\core.registers[5][25] ),
    .A1(net1111),
    .S(net500),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _17840_ (.A0(\core.registers[5][26] ),
    .A1(net1103),
    .S(net501),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _17841_ (.A0(\core.registers[5][27] ),
    .A1(net1107),
    .S(net500),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _17842_ (.A0(\core.registers[5][28] ),
    .A1(net1097),
    .S(net500),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _17843_ (.A0(\core.registers[5][29] ),
    .A1(net1093),
    .S(net502),
    .X(_01534_));
 sky130_fd_sc_hd__mux2_1 _17844_ (.A0(\core.registers[5][30] ),
    .A1(net1087),
    .S(net503),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _17845_ (.A0(\core.registers[5][31] ),
    .A1(net1090),
    .S(net502),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _17846_ (.A0(\wbSRAMInterface.currentByteSelect[0] ),
    .A1(net247),
    .S(net1350),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _17847_ (.A0(\wbSRAMInterface.currentByteSelect[1] ),
    .A1(net248),
    .S(net1350),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _17848_ (.A0(\wbSRAMInterface.currentByteSelect[2] ),
    .A1(net249),
    .S(net1350),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _17849_ (.A0(\wbSRAMInterface.currentByteSelect[3] ),
    .A1(net250),
    .S(net1350),
    .X(_01540_));
 sky130_fd_sc_hd__nor2_1 _17850_ (.A(_04512_),
    .B(_03600_),
    .Y(_03609_));
 sky130_fd_sc_hd__and3_4 _17851_ (.A(net676),
    .B(net1073),
    .C(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__mux2_1 _17852_ (.A0(\core.registers[4][0] ),
    .A1(net1038),
    .S(net498),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _17853_ (.A0(\core.registers[4][1] ),
    .A1(net1042),
    .S(net498),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _17854_ (.A0(\core.registers[4][2] ),
    .A1(net1045),
    .S(net499),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _17855_ (.A0(\core.registers[4][3] ),
    .A1(net1048),
    .S(net498),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _17856_ (.A0(\core.registers[4][4] ),
    .A1(net1053),
    .S(net498),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _17857_ (.A0(\core.registers[4][5] ),
    .A1(net1058),
    .S(net499),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _17858_ (.A0(\core.registers[4][6] ),
    .A1(net1063),
    .S(net499),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _17859_ (.A0(\core.registers[4][7] ),
    .A1(net1133),
    .S(net499),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _17860_ (.A0(\core.registers[4][8] ),
    .A1(net959),
    .S(net499),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _17861_ (.A0(\core.registers[4][9] ),
    .A1(net964),
    .S(net497),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _17862_ (.A0(\core.registers[4][10] ),
    .A1(_05387_),
    .S(net498),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _17863_ (.A0(\core.registers[4][11] ),
    .A1(net2011),
    .S(net497),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _17864_ (.A0(\core.registers[4][12] ),
    .A1(net990),
    .S(net497),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _17865_ (.A0(\core.registers[4][13] ),
    .A1(net985),
    .S(net498),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _17866_ (.A0(\core.registers[4][14] ),
    .A1(net978),
    .S(net498),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _17867_ (.A0(\core.registers[4][15] ),
    .A1(net982),
    .S(net498),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _17868_ (.A0(\core.registers[4][16] ),
    .A1(net1126),
    .S(net496),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _17869_ (.A0(\core.registers[4][17] ),
    .A1(net1128),
    .S(net496),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _17870_ (.A0(\core.registers[4][18] ),
    .A1(net1118),
    .S(net497),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _17871_ (.A0(\core.registers[4][19] ),
    .A1(net1122),
    .S(net496),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _17872_ (.A0(\core.registers[4][20] ),
    .A1(net1138),
    .S(net496),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _17873_ (.A0(\core.registers[4][21] ),
    .A1(net1143),
    .S(net496),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _17874_ (.A0(\core.registers[4][22] ),
    .A1(net1147),
    .S(net497),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _17875_ (.A0(\core.registers[4][23] ),
    .A1(net1152),
    .S(net496),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _17876_ (.A0(\core.registers[4][24] ),
    .A1(net1115),
    .S(net496),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _17877_ (.A0(\core.registers[4][25] ),
    .A1(net1111),
    .S(net496),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _17878_ (.A0(\core.registers[4][26] ),
    .A1(net1103),
    .S(net497),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _17879_ (.A0(\core.registers[4][27] ),
    .A1(net1107),
    .S(net496),
    .X(_01568_));
 sky130_fd_sc_hd__mux2_1 _17880_ (.A0(\core.registers[4][28] ),
    .A1(net1097),
    .S(net496),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _17881_ (.A0(\core.registers[4][29] ),
    .A1(net1093),
    .S(net498),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _17882_ (.A0(\core.registers[4][30] ),
    .A1(net1087),
    .S(net499),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _17883_ (.A0(\core.registers[4][31] ),
    .A1(net1090),
    .S(net498),
    .X(_01572_));
 sky130_fd_sc_hd__nor2_1 _17884_ (.A(_04516_),
    .B(_09093_),
    .Y(_03611_));
 sky130_fd_sc_hd__and3_4 _17885_ (.A(net679),
    .B(_09085_),
    .C(_03611_),
    .X(_03612_));
 sky130_fd_sc_hd__mux2_1 _17886_ (.A0(\core.registers[3][0] ),
    .A1(net1037),
    .S(net494),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _17887_ (.A0(\core.registers[3][1] ),
    .A1(net1042),
    .S(net494),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _17888_ (.A0(\core.registers[3][2] ),
    .A1(net1045),
    .S(net494),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _17889_ (.A0(\core.registers[3][3] ),
    .A1(net1049),
    .S(net494),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _17890_ (.A0(\core.registers[3][4] ),
    .A1(net1053),
    .S(net494),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _17891_ (.A0(\core.registers[3][5] ),
    .A1(net1060),
    .S(net495),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _17892_ (.A0(\core.registers[3][6] ),
    .A1(net1063),
    .S(net495),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _17893_ (.A0(\core.registers[3][7] ),
    .A1(net1135),
    .S(net495),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _17894_ (.A0(\core.registers[3][8] ),
    .A1(net959),
    .S(net495),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _17895_ (.A0(\core.registers[3][9] ),
    .A1(net965),
    .S(net493),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _17896_ (.A0(\core.registers[3][10] ),
    .A1(net969),
    .S(net494),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _17897_ (.A0(\core.registers[3][11] ),
    .A1(net2011),
    .S(net493),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _17898_ (.A0(\core.registers[3][12] ),
    .A1(net990),
    .S(net493),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _17899_ (.A0(\core.registers[3][13] ),
    .A1(net985),
    .S(net494),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _17900_ (.A0(\core.registers[3][14] ),
    .A1(net975),
    .S(net493),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _17901_ (.A0(\core.registers[3][15] ),
    .A1(net982),
    .S(net494),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _17902_ (.A0(\core.registers[3][16] ),
    .A1(net1126),
    .S(net492),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _17903_ (.A0(\core.registers[3][17] ),
    .A1(net1129),
    .S(net492),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _17904_ (.A0(\core.registers[3][18] ),
    .A1(net1119),
    .S(net493),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _17905_ (.A0(\core.registers[3][19] ),
    .A1(net1123),
    .S(net492),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _17906_ (.A0(\core.registers[3][20] ),
    .A1(net1139),
    .S(net492),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _17907_ (.A0(\core.registers[3][21] ),
    .A1(net1143),
    .S(net492),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _17908_ (.A0(\core.registers[3][22] ),
    .A1(net1148),
    .S(net493),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _17909_ (.A0(\core.registers[3][23] ),
    .A1(net1152),
    .S(net492),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _17910_ (.A0(\core.registers[3][24] ),
    .A1(net1114),
    .S(net492),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _17911_ (.A0(\core.registers[3][25] ),
    .A1(net1109),
    .S(net492),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _17912_ (.A0(\core.registers[3][26] ),
    .A1(_06953_),
    .S(net493),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _17913_ (.A0(\core.registers[3][27] ),
    .A1(net1107),
    .S(net492),
    .X(_01600_));
 sky130_fd_sc_hd__mux2_1 _17914_ (.A0(\core.registers[3][28] ),
    .A1(net1097),
    .S(net492),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _17915_ (.A0(\core.registers[3][29] ),
    .A1(net1092),
    .S(net494),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _17916_ (.A0(\core.registers[3][30] ),
    .A1(net1087),
    .S(net495),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _17917_ (.A0(\core.registers[3][31] ),
    .A1(net1090),
    .S(net494),
    .X(_01604_));
 sky130_fd_sc_hd__nor2_1 _17918_ (.A(_09093_),
    .B(_09098_),
    .Y(_03613_));
 sky130_fd_sc_hd__and3_4 _17919_ (.A(net679),
    .B(net1074),
    .C(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__mux2_1 _17920_ (.A0(\core.registers[31][0] ),
    .A1(net1036),
    .S(net491),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _17921_ (.A0(\core.registers[31][1] ),
    .A1(net1041),
    .S(net491),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _17922_ (.A0(\core.registers[31][2] ),
    .A1(net1043),
    .S(net491),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _17923_ (.A0(\core.registers[31][3] ),
    .A1(net1050),
    .S(net490),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _17924_ (.A0(\core.registers[31][4] ),
    .A1(net1056),
    .S(net491),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _17925_ (.A0(\core.registers[31][5] ),
    .A1(net1059),
    .S(net490),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _17926_ (.A0(\core.registers[31][6] ),
    .A1(net1064),
    .S(net490),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _17927_ (.A0(\core.registers[31][7] ),
    .A1(net1134),
    .S(net490),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _17928_ (.A0(\core.registers[31][8] ),
    .A1(net957),
    .S(net490),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _17929_ (.A0(\core.registers[31][9] ),
    .A1(net962),
    .S(net489),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _17930_ (.A0(\core.registers[31][10] ),
    .A1(net966),
    .S(net491),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _17931_ (.A0(\core.registers[31][11] ),
    .A1(net970),
    .S(net489),
    .X(_01616_));
 sky130_fd_sc_hd__mux2_1 _17932_ (.A0(\core.registers[31][12] ),
    .A1(net988),
    .S(net491),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _17933_ (.A0(\core.registers[31][13] ),
    .A1(net983),
    .S(net490),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _17934_ (.A0(\core.registers[31][14] ),
    .A1(net974),
    .S(net491),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _17935_ (.A0(\core.registers[31][15] ),
    .A1(net979),
    .S(net490),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _17936_ (.A0(\core.registers[31][16] ),
    .A1(net1127),
    .S(net488),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _17937_ (.A0(\core.registers[31][17] ),
    .A1(net1131),
    .S(net488),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _17938_ (.A0(\core.registers[31][18] ),
    .A1(net1117),
    .S(net489),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _17939_ (.A0(\core.registers[31][19] ),
    .A1(net1121),
    .S(net488),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _17940_ (.A0(\core.registers[31][20] ),
    .A1(net1137),
    .S(net488),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _17941_ (.A0(\core.registers[31][21] ),
    .A1(net1141),
    .S(net488),
    .X(_01626_));
 sky130_fd_sc_hd__mux2_1 _17942_ (.A0(\core.registers[31][22] ),
    .A1(net1146),
    .S(net489),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _17943_ (.A0(\core.registers[31][23] ),
    .A1(net1150),
    .S(net488),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _17944_ (.A0(\core.registers[31][24] ),
    .A1(net1113),
    .S(net488),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _17945_ (.A0(\core.registers[31][25] ),
    .A1(net1108),
    .S(net488),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _17946_ (.A0(\core.registers[31][26] ),
    .A1(net1101),
    .S(net489),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _17947_ (.A0(\core.registers[31][27] ),
    .A1(net1104),
    .S(net488),
    .X(_01632_));
 sky130_fd_sc_hd__mux2_1 _17948_ (.A0(\core.registers[31][28] ),
    .A1(net1099),
    .S(net488),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _17949_ (.A0(\core.registers[31][29] ),
    .A1(net1095),
    .S(net490),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _17950_ (.A0(\core.registers[31][30] ),
    .A1(net1086),
    .S(net490),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _17951_ (.A0(\core.registers[31][31] ),
    .A1(net1091),
    .S(net490),
    .X(_01636_));
 sky130_fd_sc_hd__nor2_1 _17952_ (.A(net1989),
    .B(_08764_),
    .Y(_01637_));
 sky130_fd_sc_hd__and2b_1 _17953_ (.A_N(\core.csr.instretTimer.currentValue[0] ),
    .B(\core.pipe2_stall ),
    .X(_03615_));
 sky130_fd_sc_hd__and2b_1 _17954_ (.A_N(\core.pipe2_stall ),
    .B(\core.csr.instretTimer.currentValue[0] ),
    .X(_03616_));
 sky130_fd_sc_hd__nor3_1 _17955_ (.A(net1990),
    .B(_03615_),
    .C(_03616_),
    .Y(_01638_));
 sky130_fd_sc_hd__and2_1 _17956_ (.A(\core.csr.instretTimer.currentValue[1] ),
    .B(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__nor2_1 _17957_ (.A(net1991),
    .B(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__o21a_1 _17958_ (.A1(\core.csr.instretTimer.currentValue[1] ),
    .A2(_03616_),
    .B1(_03618_),
    .X(_01639_));
 sky130_fd_sc_hd__and3_1 _17959_ (.A(\core.csr.instretTimer.currentValue[2] ),
    .B(\core.csr.instretTimer.currentValue[1] ),
    .C(_03616_),
    .X(_03619_));
 sky130_fd_sc_hd__o21ai_1 _17960_ (.A1(\core.csr.instretTimer.currentValue[2] ),
    .A2(_03617_),
    .B1(net1945),
    .Y(_03620_));
 sky130_fd_sc_hd__nor2_1 _17961_ (.A(_03619_),
    .B(_03620_),
    .Y(_01640_));
 sky130_fd_sc_hd__and3_2 _17962_ (.A(\core.csr.instretTimer.currentValue[3] ),
    .B(\core.csr.instretTimer.currentValue[2] ),
    .C(_03617_),
    .X(_03621_));
 sky130_fd_sc_hd__o21ai_1 _17963_ (.A1(\core.csr.instretTimer.currentValue[3] ),
    .A2(_03619_),
    .B1(net1945),
    .Y(_03622_));
 sky130_fd_sc_hd__nor2_1 _17964_ (.A(_03621_),
    .B(_03622_),
    .Y(_01641_));
 sky130_fd_sc_hd__and2_2 _17965_ (.A(\core.csr.instretTimer.currentValue[4] ),
    .B(_03621_),
    .X(_03623_));
 sky130_fd_sc_hd__nor2_1 _17966_ (.A(net1993),
    .B(_03623_),
    .Y(_03624_));
 sky130_fd_sc_hd__o21a_1 _17967_ (.A1(\core.csr.instretTimer.currentValue[4] ),
    .A2(_03621_),
    .B1(_03624_),
    .X(_01642_));
 sky130_fd_sc_hd__a21oi_1 _17968_ (.A1(\core.csr.instretTimer.currentValue[5] ),
    .A2(_03623_),
    .B1(net1992),
    .Y(_03625_));
 sky130_fd_sc_hd__o21a_1 _17969_ (.A1(\core.csr.instretTimer.currentValue[5] ),
    .A2(_03623_),
    .B1(_03625_),
    .X(_01643_));
 sky130_fd_sc_hd__a21oi_1 _17970_ (.A1(\core.csr.instretTimer.currentValue[5] ),
    .A2(_03623_),
    .B1(\core.csr.instretTimer.currentValue[6] ),
    .Y(_03626_));
 sky130_fd_sc_hd__and3_1 _17971_ (.A(\core.csr.instretTimer.currentValue[6] ),
    .B(\core.csr.instretTimer.currentValue[5] ),
    .C(_03623_),
    .X(_03627_));
 sky130_fd_sc_hd__nor3_1 _17972_ (.A(net1992),
    .B(_03626_),
    .C(_03627_),
    .Y(_01644_));
 sky130_fd_sc_hd__and2_1 _17973_ (.A(\core.csr.instretTimer.currentValue[7] ),
    .B(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__o21ai_1 _17974_ (.A1(\core.csr.instretTimer.currentValue[7] ),
    .A2(_03627_),
    .B1(net1957),
    .Y(_03629_));
 sky130_fd_sc_hd__nor2_1 _17975_ (.A(_03628_),
    .B(_03629_),
    .Y(_01645_));
 sky130_fd_sc_hd__and3_1 _17976_ (.A(\core.csr.instretTimer.currentValue[8] ),
    .B(\core.csr.instretTimer.currentValue[7] ),
    .C(_03627_),
    .X(_03630_));
 sky130_fd_sc_hd__nor2_1 _17977_ (.A(net1992),
    .B(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__o21a_1 _17978_ (.A1(\core.csr.instretTimer.currentValue[8] ),
    .A2(_03628_),
    .B1(_03631_),
    .X(_01646_));
 sky130_fd_sc_hd__and2_1 _17979_ (.A(\core.csr.instretTimer.currentValue[9] ),
    .B(_03630_),
    .X(_03632_));
 sky130_fd_sc_hd__nor2_1 _17980_ (.A(net1997),
    .B(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hd__o21a_1 _17981_ (.A1(\core.csr.instretTimer.currentValue[9] ),
    .A2(_03630_),
    .B1(_03633_),
    .X(_01647_));
 sky130_fd_sc_hd__and3_1 _17982_ (.A(\core.csr.instretTimer.currentValue[10] ),
    .B(\core.csr.instretTimer.currentValue[9] ),
    .C(_03630_),
    .X(_03634_));
 sky130_fd_sc_hd__o21ai_1 _17983_ (.A1(\core.csr.instretTimer.currentValue[10] ),
    .A2(_03632_),
    .B1(net1959),
    .Y(_03635_));
 sky130_fd_sc_hd__nor2_1 _17984_ (.A(_03634_),
    .B(_03635_),
    .Y(_01648_));
 sky130_fd_sc_hd__and3_1 _17985_ (.A(\core.csr.instretTimer.currentValue[11] ),
    .B(\core.csr.instretTimer.currentValue[10] ),
    .C(_03632_),
    .X(_03636_));
 sky130_fd_sc_hd__nor2_1 _17986_ (.A(net1997),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__o21a_1 _17987_ (.A1(\core.csr.instretTimer.currentValue[11] ),
    .A2(_03634_),
    .B1(_03637_),
    .X(_01649_));
 sky130_fd_sc_hd__and2_1 _17988_ (.A(\core.csr.instretTimer.currentValue[12] ),
    .B(_03636_),
    .X(_03638_));
 sky130_fd_sc_hd__nor2_1 _17989_ (.A(net1997),
    .B(_03638_),
    .Y(_03639_));
 sky130_fd_sc_hd__o21a_1 _17990_ (.A1(\core.csr.instretTimer.currentValue[12] ),
    .A2(_03636_),
    .B1(_03639_),
    .X(_01650_));
 sky130_fd_sc_hd__and3_2 _17991_ (.A(\core.csr.instretTimer.currentValue[13] ),
    .B(\core.csr.instretTimer.currentValue[12] ),
    .C(_03636_),
    .X(_03640_));
 sky130_fd_sc_hd__nor2_1 _17992_ (.A(net1997),
    .B(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__o21a_1 _17993_ (.A1(\core.csr.instretTimer.currentValue[13] ),
    .A2(_03638_),
    .B1(_03641_),
    .X(_01651_));
 sky130_fd_sc_hd__and2_1 _17994_ (.A(\core.csr.instretTimer.currentValue[14] ),
    .B(_03640_),
    .X(_03642_));
 sky130_fd_sc_hd__nor2_1 _17995_ (.A(net2001),
    .B(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__o21a_1 _17996_ (.A1(\core.csr.instretTimer.currentValue[14] ),
    .A2(_03640_),
    .B1(_03643_),
    .X(_01652_));
 sky130_fd_sc_hd__and3_2 _17997_ (.A(\core.csr.instretTimer.currentValue[15] ),
    .B(\core.csr.instretTimer.currentValue[14] ),
    .C(_03640_),
    .X(_03644_));
 sky130_fd_sc_hd__nor2_1 _17998_ (.A(net2001),
    .B(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__o21a_1 _17999_ (.A1(\core.csr.instretTimer.currentValue[15] ),
    .A2(_03642_),
    .B1(_03645_),
    .X(_01653_));
 sky130_fd_sc_hd__a21oi_1 _18000_ (.A1(\core.csr.instretTimer.currentValue[16] ),
    .A2(_03644_),
    .B1(net1999),
    .Y(_03646_));
 sky130_fd_sc_hd__o21a_1 _18001_ (.A1(\core.csr.instretTimer.currentValue[16] ),
    .A2(_03644_),
    .B1(_03646_),
    .X(_01654_));
 sky130_fd_sc_hd__a21oi_1 _18002_ (.A1(\core.csr.instretTimer.currentValue[16] ),
    .A2(_03644_),
    .B1(\core.csr.instretTimer.currentValue[17] ),
    .Y(_03647_));
 sky130_fd_sc_hd__and3_1 _18003_ (.A(\core.csr.instretTimer.currentValue[17] ),
    .B(\core.csr.instretTimer.currentValue[16] ),
    .C(_03644_),
    .X(_03648_));
 sky130_fd_sc_hd__nor3_1 _18004_ (.A(net1999),
    .B(_03647_),
    .C(_03648_),
    .Y(_01655_));
 sky130_fd_sc_hd__and2_4 _18005_ (.A(\core.csr.instretTimer.currentValue[18] ),
    .B(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__nor2_1 _18006_ (.A(net1999),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hd__o21a_1 _18007_ (.A1(\core.csr.instretTimer.currentValue[18] ),
    .A2(_03648_),
    .B1(_03650_),
    .X(_01656_));
 sky130_fd_sc_hd__a21oi_1 _18008_ (.A1(\core.csr.instretTimer.currentValue[19] ),
    .A2(_03649_),
    .B1(net1973),
    .Y(_03651_));
 sky130_fd_sc_hd__o21a_1 _18009_ (.A1(\core.csr.instretTimer.currentValue[19] ),
    .A2(_03649_),
    .B1(_03651_),
    .X(_01657_));
 sky130_fd_sc_hd__a21oi_1 _18010_ (.A1(\core.csr.instretTimer.currentValue[19] ),
    .A2(_03649_),
    .B1(\core.csr.instretTimer.currentValue[20] ),
    .Y(_03652_));
 sky130_fd_sc_hd__and3_1 _18011_ (.A(\core.csr.instretTimer.currentValue[20] ),
    .B(\core.csr.instretTimer.currentValue[19] ),
    .C(_03649_),
    .X(_03653_));
 sky130_fd_sc_hd__nor3_1 _18012_ (.A(net1973),
    .B(_03652_),
    .C(_03653_),
    .Y(_01658_));
 sky130_fd_sc_hd__and2_2 _18013_ (.A(\core.csr.instretTimer.currentValue[21] ),
    .B(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__nor2_1 _18014_ (.A(net1973),
    .B(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__o21a_1 _18015_ (.A1(\core.csr.instretTimer.currentValue[21] ),
    .A2(_03653_),
    .B1(_03655_),
    .X(_01659_));
 sky130_fd_sc_hd__a21oi_1 _18016_ (.A1(\core.csr.instretTimer.currentValue[22] ),
    .A2(_03654_),
    .B1(net1972),
    .Y(_03656_));
 sky130_fd_sc_hd__o21a_1 _18017_ (.A1(\core.csr.instretTimer.currentValue[22] ),
    .A2(_03654_),
    .B1(_03656_),
    .X(_01660_));
 sky130_fd_sc_hd__a21oi_1 _18018_ (.A1(\core.csr.instretTimer.currentValue[22] ),
    .A2(_03654_),
    .B1(\core.csr.instretTimer.currentValue[23] ),
    .Y(_03657_));
 sky130_fd_sc_hd__and3_2 _18019_ (.A(\core.csr.instretTimer.currentValue[23] ),
    .B(\core.csr.instretTimer.currentValue[22] ),
    .C(_03654_),
    .X(_03658_));
 sky130_fd_sc_hd__nor3_1 _18020_ (.A(net1972),
    .B(_03657_),
    .C(_03658_),
    .Y(_01661_));
 sky130_fd_sc_hd__and2_1 _18021_ (.A(\core.csr.instretTimer.currentValue[24] ),
    .B(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__nor2_1 _18022_ (.A(net1967),
    .B(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__o21a_1 _18023_ (.A1(\core.csr.instretTimer.currentValue[24] ),
    .A2(_03658_),
    .B1(_03660_),
    .X(_01662_));
 sky130_fd_sc_hd__and3_1 _18024_ (.A(\core.csr.instretTimer.currentValue[25] ),
    .B(\core.csr.instretTimer.currentValue[24] ),
    .C(_03658_),
    .X(_03661_));
 sky130_fd_sc_hd__nor2_1 _18025_ (.A(net1967),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__o21a_1 _18026_ (.A1(\core.csr.instretTimer.currentValue[25] ),
    .A2(_03659_),
    .B1(_03662_),
    .X(_01663_));
 sky130_fd_sc_hd__and2_1 _18027_ (.A(\core.csr.instretTimer.currentValue[26] ),
    .B(_03661_),
    .X(_03663_));
 sky130_fd_sc_hd__nor2_1 _18028_ (.A(net1967),
    .B(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__o21a_1 _18029_ (.A1(\core.csr.instretTimer.currentValue[26] ),
    .A2(_03661_),
    .B1(_03664_),
    .X(_01664_));
 sky130_fd_sc_hd__and3_4 _18030_ (.A(\core.csr.instretTimer.currentValue[27] ),
    .B(\core.csr.instretTimer.currentValue[26] ),
    .C(_03661_),
    .X(_03665_));
 sky130_fd_sc_hd__nor2_1 _18031_ (.A(net1967),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__o21a_1 _18032_ (.A1(\core.csr.instretTimer.currentValue[27] ),
    .A2(_03663_),
    .B1(_03666_),
    .X(_01665_));
 sky130_fd_sc_hd__and2_1 _18033_ (.A(\core.csr.instretTimer.currentValue[28] ),
    .B(_03665_),
    .X(_03667_));
 sky130_fd_sc_hd__nor2_1 _18034_ (.A(net1987),
    .B(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__o21a_1 _18035_ (.A1(\core.csr.instretTimer.currentValue[28] ),
    .A2(_03665_),
    .B1(_03668_),
    .X(_01666_));
 sky130_fd_sc_hd__and3_2 _18036_ (.A(\core.csr.instretTimer.currentValue[29] ),
    .B(\core.csr.instretTimer.currentValue[28] ),
    .C(_03665_),
    .X(_03669_));
 sky130_fd_sc_hd__nor2_1 _18037_ (.A(net1987),
    .B(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__o21a_1 _18038_ (.A1(\core.csr.instretTimer.currentValue[29] ),
    .A2(_03667_),
    .B1(_03670_),
    .X(_01667_));
 sky130_fd_sc_hd__and2_4 _18039_ (.A(\core.csr.instretTimer.currentValue[30] ),
    .B(_03669_),
    .X(_03671_));
 sky130_fd_sc_hd__nor2_1 _18040_ (.A(net1995),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__o21a_1 _18041_ (.A1(\core.csr.instretTimer.currentValue[30] ),
    .A2(_03669_),
    .B1(_03672_),
    .X(_01668_));
 sky130_fd_sc_hd__a21oi_1 _18042_ (.A1(\core.csr.instretTimer.currentValue[31] ),
    .A2(_03671_),
    .B1(net1996),
    .Y(_03673_));
 sky130_fd_sc_hd__o21a_1 _18043_ (.A1(\core.csr.instretTimer.currentValue[31] ),
    .A2(_03671_),
    .B1(_03673_),
    .X(_01669_));
 sky130_fd_sc_hd__a21oi_1 _18044_ (.A1(\core.csr.instretTimer.currentValue[31] ),
    .A2(_03671_),
    .B1(\core.csr.instretTimer.currentValue[32] ),
    .Y(_03674_));
 sky130_fd_sc_hd__and3_1 _18045_ (.A(\core.csr.instretTimer.currentValue[32] ),
    .B(\core.csr.instretTimer.currentValue[31] ),
    .C(_03671_),
    .X(_03675_));
 sky130_fd_sc_hd__nor3_1 _18046_ (.A(net1990),
    .B(_03674_),
    .C(_03675_),
    .Y(_01670_));
 sky130_fd_sc_hd__and2_2 _18047_ (.A(\core.csr.instretTimer.currentValue[33] ),
    .B(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__nor2_1 _18048_ (.A(net1990),
    .B(_03676_),
    .Y(_03677_));
 sky130_fd_sc_hd__o21a_1 _18049_ (.A1(\core.csr.instretTimer.currentValue[33] ),
    .A2(_03675_),
    .B1(_03677_),
    .X(_01671_));
 sky130_fd_sc_hd__a21oi_1 _18050_ (.A1(\core.csr.instretTimer.currentValue[34] ),
    .A2(_03676_),
    .B1(net1991),
    .Y(_03678_));
 sky130_fd_sc_hd__o21a_1 _18051_ (.A1(\core.csr.instretTimer.currentValue[34] ),
    .A2(_03676_),
    .B1(_03678_),
    .X(_01672_));
 sky130_fd_sc_hd__a21oi_1 _18052_ (.A1(\core.csr.instretTimer.currentValue[34] ),
    .A2(_03676_),
    .B1(\core.csr.instretTimer.currentValue[35] ),
    .Y(_03679_));
 sky130_fd_sc_hd__and3_2 _18053_ (.A(\core.csr.instretTimer.currentValue[35] ),
    .B(\core.csr.instretTimer.currentValue[34] ),
    .C(_03676_),
    .X(_03680_));
 sky130_fd_sc_hd__nor3_1 _18054_ (.A(net1991),
    .B(_03679_),
    .C(_03680_),
    .Y(_01673_));
 sky130_fd_sc_hd__and2_2 _18055_ (.A(\core.csr.instretTimer.currentValue[36] ),
    .B(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__nor2_1 _18056_ (.A(net1993),
    .B(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__o21a_1 _18057_ (.A1(\core.csr.instretTimer.currentValue[36] ),
    .A2(_03680_),
    .B1(_03682_),
    .X(_01674_));
 sky130_fd_sc_hd__a21oi_1 _18058_ (.A1(\core.csr.instretTimer.currentValue[37] ),
    .A2(_03681_),
    .B1(net1993),
    .Y(_03683_));
 sky130_fd_sc_hd__o21a_1 _18059_ (.A1(\core.csr.instretTimer.currentValue[37] ),
    .A2(_03681_),
    .B1(_03683_),
    .X(_01675_));
 sky130_fd_sc_hd__a21oi_1 _18060_ (.A1(\core.csr.instretTimer.currentValue[37] ),
    .A2(_03681_),
    .B1(\core.csr.instretTimer.currentValue[38] ),
    .Y(_03684_));
 sky130_fd_sc_hd__and3_1 _18061_ (.A(\core.csr.instretTimer.currentValue[38] ),
    .B(\core.csr.instretTimer.currentValue[37] ),
    .C(_03681_),
    .X(_03685_));
 sky130_fd_sc_hd__nor3_1 _18062_ (.A(net1992),
    .B(_03684_),
    .C(_03685_),
    .Y(_01676_));
 sky130_fd_sc_hd__and2_2 _18063_ (.A(\core.csr.instretTimer.currentValue[39] ),
    .B(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__nor2_1 _18064_ (.A(net1992),
    .B(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__o21a_1 _18065_ (.A1(\core.csr.instretTimer.currentValue[39] ),
    .A2(_03685_),
    .B1(_03687_),
    .X(_01677_));
 sky130_fd_sc_hd__a21oi_1 _18066_ (.A1(\core.csr.instretTimer.currentValue[40] ),
    .A2(_03686_),
    .B1(net1993),
    .Y(_03688_));
 sky130_fd_sc_hd__o21a_1 _18067_ (.A1(\core.csr.instretTimer.currentValue[40] ),
    .A2(_03686_),
    .B1(_03688_),
    .X(_01678_));
 sky130_fd_sc_hd__a21oi_1 _18068_ (.A1(\core.csr.instretTimer.currentValue[40] ),
    .A2(_03686_),
    .B1(\core.csr.instretTimer.currentValue[41] ),
    .Y(_03689_));
 sky130_fd_sc_hd__and3_1 _18069_ (.A(\core.csr.instretTimer.currentValue[41] ),
    .B(\core.csr.instretTimer.currentValue[40] ),
    .C(_03686_),
    .X(_03690_));
 sky130_fd_sc_hd__nor3_1 _18070_ (.A(net1997),
    .B(_03689_),
    .C(_03690_),
    .Y(_01679_));
 sky130_fd_sc_hd__and2_2 _18071_ (.A(\core.csr.instretTimer.currentValue[42] ),
    .B(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__nor2_1 _18072_ (.A(net1997),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__o21a_1 _18073_ (.A1(\core.csr.instretTimer.currentValue[42] ),
    .A2(_03690_),
    .B1(_03692_),
    .X(_01680_));
 sky130_fd_sc_hd__a21oi_1 _18074_ (.A1(\core.csr.instretTimer.currentValue[43] ),
    .A2(_03691_),
    .B1(net1997),
    .Y(_03693_));
 sky130_fd_sc_hd__o21a_1 _18075_ (.A1(\core.csr.instretTimer.currentValue[43] ),
    .A2(_03691_),
    .B1(_03693_),
    .X(_01681_));
 sky130_fd_sc_hd__a21oi_1 _18076_ (.A1(\core.csr.instretTimer.currentValue[43] ),
    .A2(_03691_),
    .B1(\core.csr.instretTimer.currentValue[44] ),
    .Y(_03694_));
 sky130_fd_sc_hd__and3_1 _18077_ (.A(\core.csr.instretTimer.currentValue[44] ),
    .B(\core.csr.instretTimer.currentValue[43] ),
    .C(_03691_),
    .X(_03695_));
 sky130_fd_sc_hd__nor3_1 _18078_ (.A(net1997),
    .B(_03694_),
    .C(_03695_),
    .Y(_01682_));
 sky130_fd_sc_hd__and2_2 _18079_ (.A(\core.csr.instretTimer.currentValue[45] ),
    .B(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__nor2_1 _18080_ (.A(net1997),
    .B(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__o21a_1 _18081_ (.A1(\core.csr.instretTimer.currentValue[45] ),
    .A2(_03695_),
    .B1(_03697_),
    .X(_01683_));
 sky130_fd_sc_hd__a21oi_1 _18082_ (.A1(\core.csr.instretTimer.currentValue[46] ),
    .A2(_03696_),
    .B1(net1998),
    .Y(_03698_));
 sky130_fd_sc_hd__o21a_1 _18083_ (.A1(\core.csr.instretTimer.currentValue[46] ),
    .A2(_03696_),
    .B1(_03698_),
    .X(_01684_));
 sky130_fd_sc_hd__a21oi_1 _18084_ (.A1(\core.csr.instretTimer.currentValue[46] ),
    .A2(_03696_),
    .B1(\core.csr.instretTimer.currentValue[47] ),
    .Y(_03699_));
 sky130_fd_sc_hd__and3_1 _18085_ (.A(\core.csr.instretTimer.currentValue[47] ),
    .B(\core.csr.instretTimer.currentValue[46] ),
    .C(_03696_),
    .X(_03700_));
 sky130_fd_sc_hd__nor3_1 _18086_ (.A(net1998),
    .B(_03699_),
    .C(_03700_),
    .Y(_01685_));
 sky130_fd_sc_hd__and2_2 _18087_ (.A(\core.csr.instretTimer.currentValue[48] ),
    .B(_03700_),
    .X(_03701_));
 sky130_fd_sc_hd__nor2_1 _18088_ (.A(net1999),
    .B(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__o21a_1 _18089_ (.A1(\core.csr.instretTimer.currentValue[48] ),
    .A2(_03700_),
    .B1(_03702_),
    .X(_01686_));
 sky130_fd_sc_hd__a21oi_1 _18090_ (.A1(\core.csr.instretTimer.currentValue[49] ),
    .A2(_03701_),
    .B1(net1999),
    .Y(_03703_));
 sky130_fd_sc_hd__o21a_1 _18091_ (.A1(\core.csr.instretTimer.currentValue[49] ),
    .A2(_03701_),
    .B1(_03703_),
    .X(_01687_));
 sky130_fd_sc_hd__a21oi_1 _18092_ (.A1(\core.csr.instretTimer.currentValue[49] ),
    .A2(_03701_),
    .B1(\core.csr.instretTimer.currentValue[50] ),
    .Y(_03704_));
 sky130_fd_sc_hd__and3_4 _18093_ (.A(\core.csr.instretTimer.currentValue[50] ),
    .B(\core.csr.instretTimer.currentValue[49] ),
    .C(_03701_),
    .X(_03705_));
 sky130_fd_sc_hd__nor3_1 _18094_ (.A(net1999),
    .B(_03704_),
    .C(_03705_),
    .Y(_01688_));
 sky130_fd_sc_hd__and2_2 _18095_ (.A(\core.csr.instretTimer.currentValue[51] ),
    .B(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__nor2_1 _18096_ (.A(net1973),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__o21a_1 _18097_ (.A1(\core.csr.instretTimer.currentValue[51] ),
    .A2(_03705_),
    .B1(_03707_),
    .X(_01689_));
 sky130_fd_sc_hd__a21oi_1 _18098_ (.A1(\core.csr.instretTimer.currentValue[52] ),
    .A2(_03706_),
    .B1(net1972),
    .Y(_03708_));
 sky130_fd_sc_hd__o21a_1 _18099_ (.A1(\core.csr.instretTimer.currentValue[52] ),
    .A2(_03706_),
    .B1(_03708_),
    .X(_01690_));
 sky130_fd_sc_hd__a21oi_1 _18100_ (.A1(\core.csr.instretTimer.currentValue[52] ),
    .A2(_03706_),
    .B1(\core.csr.instretTimer.currentValue[53] ),
    .Y(_03709_));
 sky130_fd_sc_hd__and3_1 _18101_ (.A(\core.csr.instretTimer.currentValue[53] ),
    .B(\core.csr.instretTimer.currentValue[52] ),
    .C(_03706_),
    .X(_03710_));
 sky130_fd_sc_hd__nor3_1 _18102_ (.A(net1972),
    .B(_03709_),
    .C(_03710_),
    .Y(_01691_));
 sky130_fd_sc_hd__and2_2 _18103_ (.A(\core.csr.instretTimer.currentValue[54] ),
    .B(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__nor2_1 _18104_ (.A(net1972),
    .B(_03711_),
    .Y(_03712_));
 sky130_fd_sc_hd__o21a_1 _18105_ (.A1(\core.csr.instretTimer.currentValue[54] ),
    .A2(_03710_),
    .B1(_03712_),
    .X(_01692_));
 sky130_fd_sc_hd__a21oi_1 _18106_ (.A1(\core.csr.instretTimer.currentValue[55] ),
    .A2(_03711_),
    .B1(net1972),
    .Y(_03713_));
 sky130_fd_sc_hd__o21a_1 _18107_ (.A1(\core.csr.instretTimer.currentValue[55] ),
    .A2(_03711_),
    .B1(_03713_),
    .X(_01693_));
 sky130_fd_sc_hd__a21oi_1 _18108_ (.A1(\core.csr.instretTimer.currentValue[55] ),
    .A2(_03711_),
    .B1(\core.csr.instretTimer.currentValue[56] ),
    .Y(_03714_));
 sky130_fd_sc_hd__and3_1 _18109_ (.A(\core.csr.instretTimer.currentValue[56] ),
    .B(\core.csr.instretTimer.currentValue[55] ),
    .C(_03711_),
    .X(_03715_));
 sky130_fd_sc_hd__nor3_1 _18110_ (.A(net1967),
    .B(_03714_),
    .C(_03715_),
    .Y(_01694_));
 sky130_fd_sc_hd__and2_2 _18111_ (.A(\core.csr.instretTimer.currentValue[57] ),
    .B(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__nor2_1 _18112_ (.A(net1967),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__o21a_1 _18113_ (.A1(\core.csr.instretTimer.currentValue[57] ),
    .A2(_03715_),
    .B1(_03717_),
    .X(_01695_));
 sky130_fd_sc_hd__a21oi_1 _18114_ (.A1(\core.csr.instretTimer.currentValue[58] ),
    .A2(_03716_),
    .B1(net1967),
    .Y(_03718_));
 sky130_fd_sc_hd__o21a_1 _18115_ (.A1(\core.csr.instretTimer.currentValue[58] ),
    .A2(_03716_),
    .B1(_03718_),
    .X(_01696_));
 sky130_fd_sc_hd__a21oi_1 _18116_ (.A1(\core.csr.instretTimer.currentValue[58] ),
    .A2(_03716_),
    .B1(\core.csr.instretTimer.currentValue[59] ),
    .Y(_03719_));
 sky130_fd_sc_hd__and3_4 _18117_ (.A(\core.csr.instretTimer.currentValue[59] ),
    .B(\core.csr.instretTimer.currentValue[58] ),
    .C(_03716_),
    .X(_03720_));
 sky130_fd_sc_hd__nor3_1 _18118_ (.A(net1968),
    .B(_03719_),
    .C(_03720_),
    .Y(_01697_));
 sky130_fd_sc_hd__and2_1 _18119_ (.A(\core.csr.instretTimer.currentValue[60] ),
    .B(_03720_),
    .X(_03721_));
 sky130_fd_sc_hd__nor2_1 _18120_ (.A(net1995),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__o21a_1 _18121_ (.A1(\core.csr.instretTimer.currentValue[60] ),
    .A2(_03720_),
    .B1(_03722_),
    .X(_01698_));
 sky130_fd_sc_hd__and3_1 _18122_ (.A(\core.csr.instretTimer.currentValue[61] ),
    .B(\core.csr.instretTimer.currentValue[60] ),
    .C(_03720_),
    .X(_03723_));
 sky130_fd_sc_hd__nor2_1 _18123_ (.A(net1995),
    .B(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__o21a_1 _18124_ (.A1(\core.csr.instretTimer.currentValue[61] ),
    .A2(_03721_),
    .B1(_03724_),
    .X(_01699_));
 sky130_fd_sc_hd__and2_1 _18125_ (.A(\core.csr.instretTimer.currentValue[62] ),
    .B(_03723_),
    .X(_03725_));
 sky130_fd_sc_hd__nor2_1 _18126_ (.A(net1995),
    .B(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__o21a_1 _18127_ (.A1(\core.csr.instretTimer.currentValue[62] ),
    .A2(_03723_),
    .B1(_03726_),
    .X(_01700_));
 sky130_fd_sc_hd__a21oi_1 _18128_ (.A1(\core.csr.instretTimer.currentValue[63] ),
    .A2(_03725_),
    .B1(net1995),
    .Y(_03727_));
 sky130_fd_sc_hd__o21a_1 _18129_ (.A1(\core.csr.instretTimer.currentValue[63] ),
    .A2(_03725_),
    .B1(_03727_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_4 _18130_ (.A0(_07876_),
    .A1(\core.csr.currentInstruction[20] ),
    .S(net1789),
    .X(_03728_));
 sky130_fd_sc_hd__mux2_4 _18131_ (.A0(_07843_),
    .A1(\core.csr.currentInstruction[21] ),
    .S(net1789),
    .X(_03729_));
 sky130_fd_sc_hd__nand2b_1 _18132_ (.A_N(_03729_),
    .B(_03728_),
    .Y(_03730_));
 sky130_fd_sc_hd__mux2_2 _18133_ (.A0(_07870_),
    .A1(\core.csr.currentInstruction[22] ),
    .S(net1789),
    .X(_03731_));
 sky130_fd_sc_hd__and2_1 _18134_ (.A(net1789),
    .B(\core.csr.currentInstruction[23] ),
    .X(_03732_));
 sky130_fd_sc_hd__nor2_1 _18135_ (.A(_09264_),
    .B(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__nor2_1 _18136_ (.A(_07868_),
    .B(_09239_),
    .Y(_03734_));
 sky130_fd_sc_hd__a31o_1 _18137_ (.A1(net1789),
    .A2(net1775),
    .A3(net1269),
    .B1(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__and2_1 _18138_ (.A(_03733_),
    .B(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__nand2_1 _18139_ (.A(_03731_),
    .B(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__mux2_2 _18140_ (.A0(_07849_),
    .A1(\core.csr.currentInstruction[26] ),
    .S(net1792),
    .X(_03738_));
 sky130_fd_sc_hd__inv_2 _18141_ (.A(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__a21o_1 _18142_ (.A1(net1794),
    .A2(\core.csr.currentInstruction[29] ),
    .B1(_09246_),
    .X(_03740_));
 sky130_fd_sc_hd__mux2_1 _18143_ (.A0(_07851_),
    .A1(\core.csr.currentInstruction[28] ),
    .S(net1794),
    .X(_03741_));
 sky130_fd_sc_hd__nand2_2 _18144_ (.A(_03740_),
    .B(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__a21o_1 _18145_ (.A1(net1792),
    .A2(\core.csr.currentInstruction[25] ),
    .B1(_09255_),
    .X(_03743_));
 sky130_fd_sc_hd__a21o_1 _18146_ (.A1(net1792),
    .A2(\core.csr.currentInstruction[27] ),
    .B1(_09261_),
    .X(_03744_));
 sky130_fd_sc_hd__or3_1 _18147_ (.A(_03742_),
    .B(_03743_),
    .C(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_1 _18148_ (.A0(_07844_),
    .A1(\core.csr.currentInstruction[24] ),
    .S(net1792),
    .X(_03746_));
 sky130_fd_sc_hd__mux2_1 _18149_ (.A0(_07848_),
    .A1(\core.csr.currentInstruction[31] ),
    .S(net1794),
    .X(_03747_));
 sky130_fd_sc_hd__a21o_1 _18150_ (.A1(net1794),
    .A2(\core.csr.currentInstruction[30] ),
    .B1(_09252_),
    .X(_03748_));
 sky130_fd_sc_hd__nand2_1 _18151_ (.A(_03747_),
    .B(_03748_),
    .Y(_03749_));
 sky130_fd_sc_hd__and3_1 _18152_ (.A(net1790),
    .B(net1775),
    .C(net1269),
    .X(_03750_));
 sky130_fd_sc_hd__o21a_1 _18153_ (.A1(_03734_),
    .A2(_03750_),
    .B1(_03733_),
    .X(_03751_));
 sky130_fd_sc_hd__nand2_2 _18154_ (.A(_03731_),
    .B(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__or2_4 _18155_ (.A(_03730_),
    .B(_03752_),
    .X(_03753_));
 sky130_fd_sc_hd__or4b_2 _18156_ (.A(_03738_),
    .B(_03743_),
    .C(_03744_),
    .D_N(_03746_),
    .X(_03754_));
 sky130_fd_sc_hd__nor4_4 _18157_ (.A(_03742_),
    .B(_03749_),
    .C(_03753_),
    .D(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__nand2b_2 _18158_ (.A_N(net1810),
    .B(net1791),
    .Y(_03756_));
 sky130_fd_sc_hd__o21ai_4 _18159_ (.A1(net1790),
    .A2(_08770_),
    .B1(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__clkinv_2 _18160_ (.A(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__mux2_1 _18161_ (.A0(\core.csr.mconfigptr.currentValue[0] ),
    .A1(_03758_),
    .S(net852),
    .X(_03759_));
 sky130_fd_sc_hd__and2_1 _18162_ (.A(net1954),
    .B(_03759_),
    .X(_01702_));
 sky130_fd_sc_hd__nand2_1 _18163_ (.A(net1790),
    .B(_04401_),
    .Y(_03760_));
 sky130_fd_sc_hd__o21ai_2 _18164_ (.A1(net1790),
    .A2(_08779_),
    .B1(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__inv_2 _18165_ (.A(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__mux2_1 _18166_ (.A0(\core.csr.mconfigptr.currentValue[1] ),
    .A1(_03762_),
    .S(net852),
    .X(_03763_));
 sky130_fd_sc_hd__and2_1 _18167_ (.A(net1958),
    .B(_03763_),
    .X(_01703_));
 sky130_fd_sc_hd__nand2b_4 _18168_ (.A_N(\core.pipe1_resultRegister[2] ),
    .B(net1788),
    .Y(_03764_));
 sky130_fd_sc_hd__o21ai_4 _18169_ (.A1(net1788),
    .A2(_08786_),
    .B1(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__inv_2 _18170_ (.A(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__mux2_1 _18171_ (.A0(\core.csr.mconfigptr.currentValue[2] ),
    .A1(_03766_),
    .S(net852),
    .X(_03767_));
 sky130_fd_sc_hd__and2_1 _18172_ (.A(net1959),
    .B(_03767_),
    .X(_01704_));
 sky130_fd_sc_hd__nand2b_2 _18173_ (.A_N(\core.pipe1_resultRegister[3] ),
    .B(net1791),
    .Y(_03768_));
 sky130_fd_sc_hd__o21ai_4 _18174_ (.A1(net1795),
    .A2(_08795_),
    .B1(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__inv_2 _18175_ (.A(_03769_),
    .Y(_03770_));
 sky130_fd_sc_hd__mux2_1 _18176_ (.A0(\core.csr.mconfigptr.currentValue[3] ),
    .A1(_03770_),
    .S(net852),
    .X(_03771_));
 sky130_fd_sc_hd__and2_1 _18177_ (.A(net1956),
    .B(_03771_),
    .X(_01705_));
 sky130_fd_sc_hd__nand2b_4 _18178_ (.A_N(\core.pipe1_resultRegister[4] ),
    .B(net1791),
    .Y(_03772_));
 sky130_fd_sc_hd__o21ai_4 _18179_ (.A1(net1790),
    .A2(_08804_),
    .B1(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__clkinv_2 _18180_ (.A(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__mux2_1 _18181_ (.A0(\core.csr.mconfigptr.currentValue[4] ),
    .A1(_03774_),
    .S(net853),
    .X(_03775_));
 sky130_fd_sc_hd__and2_1 _18182_ (.A(net1955),
    .B(_03775_),
    .X(_01706_));
 sky130_fd_sc_hd__nand2b_2 _18183_ (.A_N(\core.pipe1_resultRegister[5] ),
    .B(net1788),
    .Y(_03776_));
 sky130_fd_sc_hd__o21ai_4 _18184_ (.A1(net1788),
    .A2(_08814_),
    .B1(_03776_),
    .Y(_03777_));
 sky130_fd_sc_hd__inv_2 _18185_ (.A(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__mux2_1 _18186_ (.A0(\core.csr.mconfigptr.currentValue[5] ),
    .A1(_03778_),
    .S(net853),
    .X(_03779_));
 sky130_fd_sc_hd__and2_1 _18187_ (.A(net1955),
    .B(_03779_),
    .X(_01707_));
 sky130_fd_sc_hd__nand2b_2 _18188_ (.A_N(\core.pipe1_resultRegister[6] ),
    .B(net1791),
    .Y(_03780_));
 sky130_fd_sc_hd__o21ai_4 _18189_ (.A1(net1789),
    .A2(_08821_),
    .B1(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__inv_2 _18190_ (.A(_03781_),
    .Y(_03782_));
 sky130_fd_sc_hd__mux2_1 _18191_ (.A0(\core.csr.mconfigptr.currentValue[6] ),
    .A1(_03782_),
    .S(net852),
    .X(_03783_));
 sky130_fd_sc_hd__and2_1 _18192_ (.A(net1954),
    .B(_03783_),
    .X(_01708_));
 sky130_fd_sc_hd__nand2b_2 _18193_ (.A_N(\core.pipe1_resultRegister[7] ),
    .B(net1788),
    .Y(_03784_));
 sky130_fd_sc_hd__o21ai_4 _18194_ (.A1(net1788),
    .A2(_08831_),
    .B1(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__inv_2 _18195_ (.A(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__mux2_1 _18196_ (.A0(\core.csr.mconfigptr.currentValue[7] ),
    .A1(_03786_),
    .S(net853),
    .X(_03787_));
 sky130_fd_sc_hd__and2_1 _18197_ (.A(net1954),
    .B(_03787_),
    .X(_01709_));
 sky130_fd_sc_hd__nand2b_2 _18198_ (.A_N(\core.pipe1_resultRegister[8] ),
    .B(net1791),
    .Y(_03788_));
 sky130_fd_sc_hd__o21ai_4 _18199_ (.A1(net1795),
    .A2(_08840_),
    .B1(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__inv_2 _18200_ (.A(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__mux2_1 _18201_ (.A0(_04396_),
    .A1(_03789_),
    .S(net852),
    .X(_03791_));
 sky130_fd_sc_hd__nor2_1 _18202_ (.A(net1994),
    .B(_03791_),
    .Y(_01710_));
 sky130_fd_sc_hd__nand2b_4 _18203_ (.A_N(\core.pipe1_resultRegister[9] ),
    .B(net1788),
    .Y(_03792_));
 sky130_fd_sc_hd__o21ai_4 _18204_ (.A1(net1796),
    .A2(_08849_),
    .B1(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__clkinv_4 _18205_ (.A(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__mux2_1 _18206_ (.A0(\core.csr.mconfigptr.currentValue[9] ),
    .A1(_03794_),
    .S(net852),
    .X(_03795_));
 sky130_fd_sc_hd__and2_1 _18207_ (.A(net1958),
    .B(_03795_),
    .X(_01711_));
 sky130_fd_sc_hd__nand2b_4 _18208_ (.A_N(\core.pipe1_resultRegister[10] ),
    .B(net1788),
    .Y(_03796_));
 sky130_fd_sc_hd__o21ai_4 _18209_ (.A1(net1796),
    .A2(_08858_),
    .B1(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__clkinv_4 _18210_ (.A(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__mux2_1 _18211_ (.A0(\core.csr.mconfigptr.currentValue[10] ),
    .A1(_03798_),
    .S(net853),
    .X(_03799_));
 sky130_fd_sc_hd__and2_1 _18212_ (.A(net1959),
    .B(_03799_),
    .X(_01712_));
 sky130_fd_sc_hd__nand2b_4 _18213_ (.A_N(\core.pipe1_resultRegister[11] ),
    .B(net1788),
    .Y(_03800_));
 sky130_fd_sc_hd__o21ai_4 _18214_ (.A1(net1788),
    .A2(_08868_),
    .B1(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__inv_4 _18215_ (.A(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__mux2_1 _18216_ (.A0(\core.csr.mconfigptr.currentValue[11] ),
    .A1(_03802_),
    .S(net852),
    .X(_03803_));
 sky130_fd_sc_hd__and2_1 _18217_ (.A(net1958),
    .B(_03803_),
    .X(_01713_));
 sky130_fd_sc_hd__nand2b_2 _18218_ (.A_N(\core.pipe1_resultRegister[12] ),
    .B(net1786),
    .Y(_03804_));
 sky130_fd_sc_hd__o21ai_4 _18219_ (.A1(net1787),
    .A2(_08877_),
    .B1(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__inv_4 _18220_ (.A(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__mux2_1 _18221_ (.A0(\core.csr.mconfigptr.currentValue[12] ),
    .A1(_03806_),
    .S(net853),
    .X(_03807_));
 sky130_fd_sc_hd__and2_1 _18222_ (.A(net1959),
    .B(_03807_),
    .X(_01714_));
 sky130_fd_sc_hd__nand2b_2 _18223_ (.A_N(\core.pipe1_resultRegister[13] ),
    .B(net1787),
    .Y(_03808_));
 sky130_fd_sc_hd__o21ai_4 _18224_ (.A1(net1787),
    .A2(_08886_),
    .B1(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__inv_4 _18225_ (.A(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__mux2_1 _18226_ (.A0(\core.csr.mconfigptr.currentValue[13] ),
    .A1(_03810_),
    .S(net852),
    .X(_03811_));
 sky130_fd_sc_hd__and2_1 _18227_ (.A(net1954),
    .B(_03811_),
    .X(_01715_));
 sky130_fd_sc_hd__nand2b_4 _18228_ (.A_N(\core.pipe1_resultRegister[14] ),
    .B(net1786),
    .Y(_03812_));
 sky130_fd_sc_hd__o21ai_4 _18229_ (.A1(net1787),
    .A2(_08895_),
    .B1(_03812_),
    .Y(_03813_));
 sky130_fd_sc_hd__clkinv_4 _18230_ (.A(_03813_),
    .Y(_03814_));
 sky130_fd_sc_hd__mux2_1 _18231_ (.A0(\core.csr.mconfigptr.currentValue[14] ),
    .A1(_03814_),
    .S(net853),
    .X(_03815_));
 sky130_fd_sc_hd__and2_1 _18232_ (.A(net1955),
    .B(_03815_),
    .X(_01716_));
 sky130_fd_sc_hd__nand2b_4 _18233_ (.A_N(\core.pipe1_resultRegister[15] ),
    .B(net1786),
    .Y(_03816_));
 sky130_fd_sc_hd__o21ai_4 _18234_ (.A1(net1786),
    .A2(_08904_),
    .B1(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__inv_4 _18235_ (.A(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__mux2_1 _18236_ (.A0(\core.csr.mconfigptr.currentValue[15] ),
    .A1(_03818_),
    .S(net852),
    .X(_03819_));
 sky130_fd_sc_hd__and2_1 _18237_ (.A(net1956),
    .B(_03819_),
    .X(_01717_));
 sky130_fd_sc_hd__nand2b_2 _18238_ (.A_N(\core.pipe1_resultRegister[16] ),
    .B(net1786),
    .Y(_03820_));
 sky130_fd_sc_hd__o21ai_4 _18239_ (.A1(net1786),
    .A2(_08915_),
    .B1(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__inv_2 _18240_ (.A(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__mux2_1 _18241_ (.A0(\core.csr.mconfigptr.currentValue[16] ),
    .A1(_03822_),
    .S(net851),
    .X(_03823_));
 sky130_fd_sc_hd__and2_1 _18242_ (.A(net1917),
    .B(_03823_),
    .X(_01718_));
 sky130_fd_sc_hd__nand2b_2 _18243_ (.A_N(\core.pipe1_resultRegister[17] ),
    .B(net1786),
    .Y(_03824_));
 sky130_fd_sc_hd__o21ai_4 _18244_ (.A1(net1786),
    .A2(_08923_),
    .B1(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__inv_2 _18245_ (.A(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__mux2_1 _18246_ (.A0(\core.csr.mconfigptr.currentValue[17] ),
    .A1(_03826_),
    .S(net850),
    .X(_03827_));
 sky130_fd_sc_hd__and2_1 _18247_ (.A(net1916),
    .B(_03827_),
    .X(_01719_));
 sky130_fd_sc_hd__nand2b_2 _18248_ (.A_N(\core.pipe1_resultRegister[18] ),
    .B(net1786),
    .Y(_03828_));
 sky130_fd_sc_hd__o21ai_4 _18249_ (.A1(net1786),
    .A2(_08932_),
    .B1(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__clkinv_2 _18250_ (.A(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__mux2_1 _18251_ (.A0(\core.csr.mconfigptr.currentValue[18] ),
    .A1(_03830_),
    .S(net851),
    .X(_03831_));
 sky130_fd_sc_hd__and2_1 _18252_ (.A(net1912),
    .B(_03831_),
    .X(_01720_));
 sky130_fd_sc_hd__nand2b_2 _18253_ (.A_N(\core.pipe1_resultRegister[19] ),
    .B(net1785),
    .Y(_03832_));
 sky130_fd_sc_hd__o21ai_4 _18254_ (.A1(net1785),
    .A2(_08943_),
    .B1(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__clkinv_2 _18255_ (.A(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__mux2_1 _18256_ (.A0(\core.csr.mconfigptr.currentValue[19] ),
    .A1(_03834_),
    .S(net850),
    .X(_03835_));
 sky130_fd_sc_hd__and2_1 _18257_ (.A(net1911),
    .B(_03835_),
    .X(_01721_));
 sky130_fd_sc_hd__nand2b_4 _18258_ (.A_N(\core.pipe1_resultRegister[20] ),
    .B(net1783),
    .Y(_03836_));
 sky130_fd_sc_hd__o21ai_4 _18259_ (.A1(net1784),
    .A2(_08952_),
    .B1(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__inv_2 _18260_ (.A(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__mux2_1 _18261_ (.A0(\core.csr.mconfigptr.currentValue[20] ),
    .A1(_03838_),
    .S(net850),
    .X(_03839_));
 sky130_fd_sc_hd__and2_1 _18262_ (.A(net1911),
    .B(_03839_),
    .X(_01722_));
 sky130_fd_sc_hd__nand2b_2 _18263_ (.A_N(\core.pipe1_resultRegister[21] ),
    .B(net1783),
    .Y(_03840_));
 sky130_fd_sc_hd__o21ai_4 _18264_ (.A1(net1784),
    .A2(_08961_),
    .B1(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__inv_2 _18265_ (.A(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__mux2_1 _18266_ (.A0(\core.csr.mconfigptr.currentValue[21] ),
    .A1(_03842_),
    .S(net850),
    .X(_03843_));
 sky130_fd_sc_hd__and2_1 _18267_ (.A(net1911),
    .B(_03843_),
    .X(_01723_));
 sky130_fd_sc_hd__nand2b_2 _18268_ (.A_N(\core.pipe1_resultRegister[22] ),
    .B(net1783),
    .Y(_03844_));
 sky130_fd_sc_hd__o21ai_4 _18269_ (.A1(net1784),
    .A2(_08970_),
    .B1(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__inv_2 _18270_ (.A(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__mux2_1 _18271_ (.A0(\core.csr.mconfigptr.currentValue[22] ),
    .A1(_03846_),
    .S(net850),
    .X(_03847_));
 sky130_fd_sc_hd__and2_1 _18272_ (.A(net1912),
    .B(_03847_),
    .X(_01724_));
 sky130_fd_sc_hd__nand2b_2 _18273_ (.A_N(\core.pipe1_resultRegister[23] ),
    .B(net1783),
    .Y(_03848_));
 sky130_fd_sc_hd__o21ai_4 _18274_ (.A1(net1784),
    .A2(_08979_),
    .B1(_03848_),
    .Y(_03849_));
 sky130_fd_sc_hd__inv_2 _18275_ (.A(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__mux2_1 _18276_ (.A0(\core.csr.mconfigptr.currentValue[23] ),
    .A1(_03850_),
    .S(net850),
    .X(_03851_));
 sky130_fd_sc_hd__and2_1 _18277_ (.A(net1912),
    .B(_03851_),
    .X(_01725_));
 sky130_fd_sc_hd__nand2b_2 _18278_ (.A_N(\core.pipe1_resultRegister[24] ),
    .B(net1783),
    .Y(_03852_));
 sky130_fd_sc_hd__o21ai_4 _18279_ (.A1(net1784),
    .A2(_08990_),
    .B1(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__inv_2 _18280_ (.A(_03853_),
    .Y(_03854_));
 sky130_fd_sc_hd__mux2_1 _18281_ (.A0(\core.csr.mconfigptr.currentValue[24] ),
    .A1(_03854_),
    .S(net850),
    .X(_03855_));
 sky130_fd_sc_hd__and2_1 _18282_ (.A(net1903),
    .B(_03855_),
    .X(_01726_));
 sky130_fd_sc_hd__nand2b_2 _18283_ (.A_N(\core.pipe1_resultRegister[25] ),
    .B(net1783),
    .Y(_03856_));
 sky130_fd_sc_hd__o21ai_4 _18284_ (.A1(net1784),
    .A2(_08998_),
    .B1(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__clkinv_2 _18285_ (.A(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__mux2_1 _18286_ (.A0(\core.csr.mconfigptr.currentValue[25] ),
    .A1(_03858_),
    .S(net850),
    .X(_03859_));
 sky130_fd_sc_hd__and2_1 _18287_ (.A(net1901),
    .B(_03859_),
    .X(_01727_));
 sky130_fd_sc_hd__nand2b_2 _18288_ (.A_N(\core.pipe1_resultRegister[26] ),
    .B(net1783),
    .Y(_03860_));
 sky130_fd_sc_hd__o21ai_4 _18289_ (.A1(net1784),
    .A2(_09007_),
    .B1(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__clkinv_2 _18290_ (.A(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__mux2_1 _18291_ (.A0(\core.csr.mconfigptr.currentValue[26] ),
    .A1(_03862_),
    .S(net850),
    .X(_03863_));
 sky130_fd_sc_hd__and2_1 _18292_ (.A(net1901),
    .B(_03863_),
    .X(_01728_));
 sky130_fd_sc_hd__nand2b_2 _18293_ (.A_N(\core.pipe1_resultRegister[27] ),
    .B(net1785),
    .Y(_03864_));
 sky130_fd_sc_hd__o21ai_4 _18294_ (.A1(net1785),
    .A2(_09016_),
    .B1(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__inv_2 _18295_ (.A(_03865_),
    .Y(_03866_));
 sky130_fd_sc_hd__mux2_1 _18296_ (.A0(\core.csr.mconfigptr.currentValue[27] ),
    .A1(_03866_),
    .S(net850),
    .X(_03867_));
 sky130_fd_sc_hd__and2_1 _18297_ (.A(net1903),
    .B(_03867_),
    .X(_01729_));
 sky130_fd_sc_hd__nand2b_2 _18298_ (.A_N(\core.pipe1_resultRegister[28] ),
    .B(net1783),
    .Y(_03868_));
 sky130_fd_sc_hd__o21ai_4 _18299_ (.A1(net1784),
    .A2(_09023_),
    .B1(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__clkinv_4 _18300_ (.A(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__mux2_1 _18301_ (.A0(\core.csr.mconfigptr.currentValue[28] ),
    .A1(_03870_),
    .S(net851),
    .X(_03871_));
 sky130_fd_sc_hd__and2_1 _18302_ (.A(net1916),
    .B(_03871_),
    .X(_01730_));
 sky130_fd_sc_hd__nand2b_2 _18303_ (.A_N(\core.pipe1_resultRegister[29] ),
    .B(net1785),
    .Y(_03872_));
 sky130_fd_sc_hd__o21ai_4 _18304_ (.A1(net1785),
    .A2(_09034_),
    .B1(_03872_),
    .Y(_03873_));
 sky130_fd_sc_hd__clkinv_4 _18305_ (.A(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__mux2_1 _18306_ (.A0(\core.csr.mconfigptr.currentValue[29] ),
    .A1(_03874_),
    .S(net851),
    .X(_03875_));
 sky130_fd_sc_hd__and2_1 _18307_ (.A(net1917),
    .B(_03875_),
    .X(_01731_));
 sky130_fd_sc_hd__nand2b_2 _18308_ (.A_N(\core.pipe1_resultRegister[30] ),
    .B(net1783),
    .Y(_03876_));
 sky130_fd_sc_hd__o21ai_4 _18309_ (.A1(net1783),
    .A2(_09043_),
    .B1(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__clkinv_8 _18310_ (.A(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__mux2_1 _18311_ (.A0(\core.csr.mconfigptr.currentValue[30] ),
    .A1(_03878_),
    .S(net853),
    .X(_03879_));
 sky130_fd_sc_hd__and2_1 _18312_ (.A(net1936),
    .B(_03879_),
    .X(_01732_));
 sky130_fd_sc_hd__nand2b_2 _18313_ (.A_N(\core.pipe1_resultRegister[31] ),
    .B(net1785),
    .Y(_03880_));
 sky130_fd_sc_hd__o21ai_4 _18314_ (.A1(net1785),
    .A2(_09052_),
    .B1(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__clkinv_4 _18315_ (.A(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__mux2_1 _18316_ (.A0(\core.csr.mconfigptr.currentValue[31] ),
    .A1(_03882_),
    .S(net851),
    .X(_03883_));
 sky130_fd_sc_hd__and2_1 _18317_ (.A(net1932),
    .B(_03883_),
    .X(_01733_));
 sky130_fd_sc_hd__or3_1 _18318_ (.A(_03746_),
    .B(_03747_),
    .C(_03748_),
    .X(_03884_));
 sky130_fd_sc_hd__or3_4 _18319_ (.A(_03739_),
    .B(_03745_),
    .C(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__or2_4 _18320_ (.A(_03728_),
    .B(_03729_),
    .X(_03886_));
 sky130_fd_sc_hd__or3b_1 _18321_ (.A(_03886_),
    .B(_03731_),
    .C_N(_03736_),
    .X(_03887_));
 sky130_fd_sc_hd__or4b_2 _18322_ (.A(_09264_),
    .B(_03731_),
    .C(_03732_),
    .D_N(_03735_),
    .X(_03888_));
 sky130_fd_sc_hd__or3b_4 _18323_ (.A(_03885_),
    .B(_03731_),
    .C_N(_03751_),
    .X(_03889_));
 sky130_fd_sc_hd__nor2_8 _18324_ (.A(_03886_),
    .B(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hd__nand2_1 _18325_ (.A(_03757_),
    .B(net848),
    .Y(_03891_));
 sky130_fd_sc_hd__o211a_1 _18326_ (.A1(\core.csr.traps.mscratch.currentValue[0] ),
    .A2(net848),
    .B1(_03891_),
    .C1(net1953),
    .X(_01734_));
 sky130_fd_sc_hd__nand2_1 _18327_ (.A(_03761_),
    .B(net848),
    .Y(_03892_));
 sky130_fd_sc_hd__o211a_1 _18328_ (.A1(\core.csr.traps.mscratch.currentValue[1] ),
    .A2(net849),
    .B1(_03892_),
    .C1(net1935),
    .X(_01735_));
 sky130_fd_sc_hd__nand2_1 _18329_ (.A(_03765_),
    .B(net848),
    .Y(_03893_));
 sky130_fd_sc_hd__o211a_1 _18330_ (.A1(\core.csr.traps.mscratch.currentValue[2] ),
    .A2(net848),
    .B1(_03893_),
    .C1(net1937),
    .X(_01736_));
 sky130_fd_sc_hd__nand2_1 _18331_ (.A(_03769_),
    .B(net848),
    .Y(_03894_));
 sky130_fd_sc_hd__o211a_1 _18332_ (.A1(\core.csr.traps.mscratch.currentValue[3] ),
    .A2(net848),
    .B1(_03894_),
    .C1(net1934),
    .X(_01737_));
 sky130_fd_sc_hd__nand2_1 _18333_ (.A(_03773_),
    .B(net848),
    .Y(_03895_));
 sky130_fd_sc_hd__o211a_1 _18334_ (.A1(\core.csr.traps.mscratch.currentValue[4] ),
    .A2(net848),
    .B1(_03895_),
    .C1(net1936),
    .X(_01738_));
 sky130_fd_sc_hd__nand2_1 _18335_ (.A(_03777_),
    .B(net847),
    .Y(_03896_));
 sky130_fd_sc_hd__o211a_1 _18336_ (.A1(\core.csr.traps.mscratch.currentValue[5] ),
    .A2(net847),
    .B1(_03896_),
    .C1(net1933),
    .X(_01739_));
 sky130_fd_sc_hd__nand2_1 _18337_ (.A(_03781_),
    .B(net849),
    .Y(_03897_));
 sky130_fd_sc_hd__o211a_1 _18338_ (.A1(\core.csr.traps.mscratch.currentValue[6] ),
    .A2(net849),
    .B1(_03897_),
    .C1(net1953),
    .X(_01740_));
 sky130_fd_sc_hd__nand2_1 _18339_ (.A(_03785_),
    .B(net847),
    .Y(_03898_));
 sky130_fd_sc_hd__o211a_1 _18340_ (.A1(\core.csr.traps.mscratch.currentValue[7] ),
    .A2(net847),
    .B1(_03898_),
    .C1(net1930),
    .X(_01741_));
 sky130_fd_sc_hd__nand2_1 _18341_ (.A(_03789_),
    .B(net848),
    .Y(_03899_));
 sky130_fd_sc_hd__o211a_1 _18342_ (.A1(\core.csr.traps.mscratch.currentValue[8] ),
    .A2(net849),
    .B1(_03899_),
    .C1(net1955),
    .X(_01742_));
 sky130_fd_sc_hd__nand2_1 _18343_ (.A(_03793_),
    .B(net849),
    .Y(_03900_));
 sky130_fd_sc_hd__o211a_1 _18344_ (.A1(\core.csr.traps.mscratch.currentValue[9] ),
    .A2(net849),
    .B1(_03900_),
    .C1(net1930),
    .X(_01743_));
 sky130_fd_sc_hd__nand2_1 _18345_ (.A(_03797_),
    .B(net847),
    .Y(_03901_));
 sky130_fd_sc_hd__o211a_1 _18346_ (.A1(\core.csr.traps.mscratch.currentValue[10] ),
    .A2(net847),
    .B1(_03901_),
    .C1(net1932),
    .X(_01744_));
 sky130_fd_sc_hd__nand2_1 _18347_ (.A(_03801_),
    .B(net847),
    .Y(_03902_));
 sky130_fd_sc_hd__o211a_1 _18348_ (.A1(\core.csr.traps.mscratch.currentValue[11] ),
    .A2(net847),
    .B1(_03902_),
    .C1(net1914),
    .X(_01745_));
 sky130_fd_sc_hd__nand2_1 _18349_ (.A(_03805_),
    .B(net847),
    .Y(_03903_));
 sky130_fd_sc_hd__o211a_1 _18350_ (.A1(\core.csr.traps.mscratch.currentValue[12] ),
    .A2(net847),
    .B1(_03903_),
    .C1(net1917),
    .X(_01746_));
 sky130_fd_sc_hd__nand2_1 _18351_ (.A(_03809_),
    .B(net845),
    .Y(_03904_));
 sky130_fd_sc_hd__o211a_1 _18352_ (.A1(\core.csr.traps.mscratch.currentValue[13] ),
    .A2(net845),
    .B1(_03904_),
    .C1(net1915),
    .X(_01747_));
 sky130_fd_sc_hd__nand2_1 _18353_ (.A(_03813_),
    .B(net845),
    .Y(_03905_));
 sky130_fd_sc_hd__o211a_1 _18354_ (.A1(\core.csr.traps.mscratch.currentValue[14] ),
    .A2(net845),
    .B1(_03905_),
    .C1(net1916),
    .X(_01748_));
 sky130_fd_sc_hd__nand2_1 _18355_ (.A(_03817_),
    .B(net846),
    .Y(_03906_));
 sky130_fd_sc_hd__o211a_1 _18356_ (.A1(\core.csr.traps.mscratch.currentValue[15] ),
    .A2(net846),
    .B1(_03906_),
    .C1(net1912),
    .X(_01749_));
 sky130_fd_sc_hd__nand2_1 _18357_ (.A(_03821_),
    .B(net846),
    .Y(_03907_));
 sky130_fd_sc_hd__o211a_1 _18358_ (.A1(\core.csr.traps.mscratch.currentValue[16] ),
    .A2(net846),
    .B1(_03907_),
    .C1(net1912),
    .X(_01750_));
 sky130_fd_sc_hd__nand2_1 _18359_ (.A(_03825_),
    .B(net845),
    .Y(_03908_));
 sky130_fd_sc_hd__o211a_1 _18360_ (.A1(\core.csr.traps.mscratch.currentValue[17] ),
    .A2(net845),
    .B1(_03908_),
    .C1(net1911),
    .X(_01751_));
 sky130_fd_sc_hd__nand2_1 _18361_ (.A(_03829_),
    .B(net845),
    .Y(_03909_));
 sky130_fd_sc_hd__o211a_1 _18362_ (.A1(\core.csr.traps.mscratch.currentValue[18] ),
    .A2(net845),
    .B1(_03909_),
    .C1(net1911),
    .X(_01752_));
 sky130_fd_sc_hd__nand2_1 _18363_ (.A(_03833_),
    .B(net845),
    .Y(_03910_));
 sky130_fd_sc_hd__o211a_1 _18364_ (.A1(\core.csr.traps.mscratch.currentValue[19] ),
    .A2(net845),
    .B1(_03910_),
    .C1(net1903),
    .X(_01753_));
 sky130_fd_sc_hd__nand2_1 _18365_ (.A(_03837_),
    .B(net843),
    .Y(_03911_));
 sky130_fd_sc_hd__o211a_1 _18366_ (.A1(\core.csr.traps.mscratch.currentValue[20] ),
    .A2(net843),
    .B1(_03911_),
    .C1(net1897),
    .X(_01754_));
 sky130_fd_sc_hd__nand2_1 _18367_ (.A(_03841_),
    .B(net842),
    .Y(_03912_));
 sky130_fd_sc_hd__o211a_1 _18368_ (.A1(\core.csr.traps.mscratch.currentValue[21] ),
    .A2(net842),
    .B1(_03912_),
    .C1(net1895),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_1 _18369_ (.A(_03845_),
    .B(net842),
    .Y(_03913_));
 sky130_fd_sc_hd__o211a_1 _18370_ (.A1(\core.csr.traps.mscratch.currentValue[22] ),
    .A2(net842),
    .B1(_03913_),
    .C1(net1895),
    .X(_01756_));
 sky130_fd_sc_hd__nand2_1 _18371_ (.A(_03849_),
    .B(net843),
    .Y(_03914_));
 sky130_fd_sc_hd__o211a_1 _18372_ (.A1(\core.csr.traps.mscratch.currentValue[23] ),
    .A2(net843),
    .B1(_03914_),
    .C1(net1897),
    .X(_01757_));
 sky130_fd_sc_hd__nand2_1 _18373_ (.A(_03853_),
    .B(net842),
    .Y(_03915_));
 sky130_fd_sc_hd__o211a_1 _18374_ (.A1(\core.csr.traps.mscratch.currentValue[24] ),
    .A2(net842),
    .B1(_03915_),
    .C1(net1896),
    .X(_01758_));
 sky130_fd_sc_hd__nand2_1 _18375_ (.A(_03857_),
    .B(net843),
    .Y(_03916_));
 sky130_fd_sc_hd__o211a_1 _18376_ (.A1(\core.csr.traps.mscratch.currentValue[25] ),
    .A2(net843),
    .B1(_03916_),
    .C1(net1902),
    .X(_01759_));
 sky130_fd_sc_hd__nand2_1 _18377_ (.A(_03861_),
    .B(net844),
    .Y(_03917_));
 sky130_fd_sc_hd__o211a_1 _18378_ (.A1(\core.csr.traps.mscratch.currentValue[26] ),
    .A2(net844),
    .B1(_03917_),
    .C1(net1902),
    .X(_01760_));
 sky130_fd_sc_hd__nand2_1 _18379_ (.A(_03865_),
    .B(net844),
    .Y(_03918_));
 sky130_fd_sc_hd__o211a_1 _18380_ (.A1(\core.csr.traps.mscratch.currentValue[27] ),
    .A2(net844),
    .B1(_03918_),
    .C1(net1903),
    .X(_01761_));
 sky130_fd_sc_hd__nand2_1 _18381_ (.A(_03869_),
    .B(net842),
    .Y(_03919_));
 sky130_fd_sc_hd__o211a_1 _18382_ (.A1(\core.csr.traps.mscratch.currentValue[28] ),
    .A2(net842),
    .B1(_03919_),
    .C1(net1897),
    .X(_01762_));
 sky130_fd_sc_hd__nand2_1 _18383_ (.A(_03873_),
    .B(net844),
    .Y(_03920_));
 sky130_fd_sc_hd__o211a_1 _18384_ (.A1(\core.csr.traps.mscratch.currentValue[29] ),
    .A2(net844),
    .B1(_03920_),
    .C1(net1902),
    .X(_01763_));
 sky130_fd_sc_hd__nand2_1 _18385_ (.A(_03877_),
    .B(net842),
    .Y(_03921_));
 sky130_fd_sc_hd__o211a_1 _18386_ (.A1(\core.csr.traps.mscratch.currentValue[30] ),
    .A2(net842),
    .B1(_03921_),
    .C1(net1896),
    .X(_01764_));
 sky130_fd_sc_hd__nand2_1 _18387_ (.A(_03881_),
    .B(net844),
    .Y(_03922_));
 sky130_fd_sc_hd__o211a_1 _18388_ (.A1(\core.csr.traps.mscratch.currentValue[31] ),
    .A2(net844),
    .B1(_03922_),
    .C1(net1903),
    .X(_01765_));
 sky130_fd_sc_hd__or3_4 _18389_ (.A(_03738_),
    .B(_03745_),
    .C(_03884_),
    .X(_03923_));
 sky130_fd_sc_hd__nor3_4 _18390_ (.A(_03752_),
    .B(_03886_),
    .C(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__mux2_1 _18391_ (.A0(\core.csr.traps.mie.currentValue[0] ),
    .A1(_03758_),
    .S(net894),
    .X(_03925_));
 sky130_fd_sc_hd__and2_1 _18392_ (.A(net1956),
    .B(_03925_),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _18393_ (.A0(\core.csr.traps.mie.currentValue[1] ),
    .A1(_03762_),
    .S(net894),
    .X(_03926_));
 sky130_fd_sc_hd__and2_1 _18394_ (.A(net1958),
    .B(_03926_),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _18395_ (.A0(\core.csr.traps.mie.currentValue[2] ),
    .A1(_03766_),
    .S(_03924_),
    .X(_03927_));
 sky130_fd_sc_hd__and2_1 _18396_ (.A(net1937),
    .B(_03927_),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _18397_ (.A0(\core.csr.traps.mie.currentValue[3] ),
    .A1(_03770_),
    .S(net894),
    .X(_03928_));
 sky130_fd_sc_hd__and2_1 _18398_ (.A(net1954),
    .B(_03928_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _18399_ (.A0(\core.csr.traps.mie.currentValue[4] ),
    .A1(_03774_),
    .S(net894),
    .X(_03929_));
 sky130_fd_sc_hd__and2_1 _18400_ (.A(net1955),
    .B(_03929_),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_1 _18401_ (.A0(\core.csr.traps.mie.currentValue[5] ),
    .A1(_03778_),
    .S(net895),
    .X(_03930_));
 sky130_fd_sc_hd__and2_1 _18402_ (.A(net1955),
    .B(_03930_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _18403_ (.A0(\core.csr.traps.mie.currentValue[6] ),
    .A1(_03782_),
    .S(net894),
    .X(_03931_));
 sky130_fd_sc_hd__and2_1 _18404_ (.A(net1954),
    .B(_03931_),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_1 _18405_ (.A0(\core.csr.traps.mie.currentValue[7] ),
    .A1(_03786_),
    .S(net895),
    .X(_03932_));
 sky130_fd_sc_hd__and2_1 _18406_ (.A(net1954),
    .B(_03932_),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_1 _18407_ (.A0(\core.csr.traps.mie.currentValue[8] ),
    .A1(_03790_),
    .S(net895),
    .X(_03933_));
 sky130_fd_sc_hd__and2_1 _18408_ (.A(net1955),
    .B(_03933_),
    .X(_01774_));
 sky130_fd_sc_hd__mux2_1 _18409_ (.A0(\core.csr.traps.mie.currentValue[9] ),
    .A1(_03794_),
    .S(net895),
    .X(_03934_));
 sky130_fd_sc_hd__and2_1 _18410_ (.A(net1958),
    .B(_03934_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _18411_ (.A0(\core.csr.traps.mie.currentValue[10] ),
    .A1(_03798_),
    .S(net894),
    .X(_03935_));
 sky130_fd_sc_hd__and2_1 _18412_ (.A(net1959),
    .B(_03935_),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _18413_ (.A0(\core.csr.traps.mie.currentValue[11] ),
    .A1(_03802_),
    .S(net894),
    .X(_03936_));
 sky130_fd_sc_hd__and2_1 _18414_ (.A(net1958),
    .B(_03936_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _18415_ (.A0(\core.csr.traps.mie.currentValue[12] ),
    .A1(_03806_),
    .S(net894),
    .X(_03937_));
 sky130_fd_sc_hd__and2_1 _18416_ (.A(net1959),
    .B(_03937_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _18417_ (.A0(\core.csr.traps.mie.currentValue[13] ),
    .A1(_03810_),
    .S(net894),
    .X(_03938_));
 sky130_fd_sc_hd__and2_1 _18418_ (.A(net1954),
    .B(_03938_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _18419_ (.A0(\core.csr.traps.mie.currentValue[14] ),
    .A1(_03814_),
    .S(net895),
    .X(_03939_));
 sky130_fd_sc_hd__and2_1 _18420_ (.A(net1955),
    .B(_03939_),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _18421_ (.A0(\core.csr.traps.mie.currentValue[15] ),
    .A1(_03818_),
    .S(net894),
    .X(_03940_));
 sky130_fd_sc_hd__and2_1 _18422_ (.A(net1956),
    .B(_03940_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _18423_ (.A0(\core.csr.traps.mie.currentValue[16] ),
    .A1(_03822_),
    .S(net893),
    .X(_03941_));
 sky130_fd_sc_hd__and2_1 _18424_ (.A(net1912),
    .B(_03941_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _18425_ (.A0(\core.csr.traps.mie.currentValue[17] ),
    .A1(_03826_),
    .S(net893),
    .X(_03942_));
 sky130_fd_sc_hd__and2_1 _18426_ (.A(net1911),
    .B(_03942_),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _18427_ (.A0(\core.csr.traps.mie.currentValue[18] ),
    .A1(_03830_),
    .S(net893),
    .X(_03943_));
 sky130_fd_sc_hd__and2_1 _18428_ (.A(net1911),
    .B(_03943_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _18429_ (.A0(\core.csr.traps.mie.currentValue[19] ),
    .A1(_03834_),
    .S(net892),
    .X(_03944_));
 sky130_fd_sc_hd__and2_1 _18430_ (.A(net1903),
    .B(_03944_),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _18431_ (.A0(\core.csr.traps.mie.currentValue[20] ),
    .A1(_03838_),
    .S(net892),
    .X(_03945_));
 sky130_fd_sc_hd__and2_1 _18432_ (.A(net1898),
    .B(_03945_),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _18433_ (.A0(\core.csr.traps.mie.currentValue[21] ),
    .A1(_03842_),
    .S(net892),
    .X(_03946_));
 sky130_fd_sc_hd__and2_1 _18434_ (.A(net1896),
    .B(_03946_),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _18435_ (.A0(\core.csr.traps.mie.currentValue[22] ),
    .A1(_03846_),
    .S(net892),
    .X(_03947_));
 sky130_fd_sc_hd__and2_1 _18436_ (.A(net1896),
    .B(_03947_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _18437_ (.A0(\core.csr.traps.mie.currentValue[23] ),
    .A1(_03850_),
    .S(net892),
    .X(_03948_));
 sky130_fd_sc_hd__and2_1 _18438_ (.A(net1896),
    .B(_03948_),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _18439_ (.A0(\core.csr.traps.mie.currentValue[24] ),
    .A1(_03854_),
    .S(net892),
    .X(_03949_));
 sky130_fd_sc_hd__and2_1 _18440_ (.A(net1895),
    .B(_03949_),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _18441_ (.A0(\core.csr.traps.mie.currentValue[25] ),
    .A1(_03858_),
    .S(net892),
    .X(_03950_));
 sky130_fd_sc_hd__and2_1 _18442_ (.A(net1897),
    .B(_03950_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _18443_ (.A0(\core.csr.traps.mie.currentValue[26] ),
    .A1(_03862_),
    .S(net893),
    .X(_03951_));
 sky130_fd_sc_hd__and2_1 _18444_ (.A(net1901),
    .B(_03951_),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _18445_ (.A0(\core.csr.traps.mie.currentValue[27] ),
    .A1(_03866_),
    .S(net893),
    .X(_03952_));
 sky130_fd_sc_hd__and2_1 _18446_ (.A(net1902),
    .B(_03952_),
    .X(_01793_));
 sky130_fd_sc_hd__mux2_1 _18447_ (.A0(\core.csr.traps.mie.currentValue[28] ),
    .A1(_03870_),
    .S(net892),
    .X(_03953_));
 sky130_fd_sc_hd__and2_1 _18448_ (.A(net1898),
    .B(_03953_),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _18449_ (.A0(\core.csr.traps.mie.currentValue[29] ),
    .A1(_03874_),
    .S(net893),
    .X(_03954_));
 sky130_fd_sc_hd__and2_1 _18450_ (.A(net1901),
    .B(_03954_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _18451_ (.A0(\core.csr.traps.mie.currentValue[30] ),
    .A1(_03878_),
    .S(net892),
    .X(_03955_));
 sky130_fd_sc_hd__and2_1 _18452_ (.A(net1895),
    .B(_03955_),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _18453_ (.A0(\core.csr.traps.mie.currentValue[31] ),
    .A1(_03882_),
    .S(net892),
    .X(_03956_));
 sky130_fd_sc_hd__and2_1 _18454_ (.A(net1901),
    .B(_03956_),
    .X(_01797_));
 sky130_fd_sc_hd__o311a_1 _18455_ (.A1(_07437_),
    .A2(_07443_),
    .A3(_07500_),
    .B1(_07468_),
    .C1(net782),
    .X(_03957_));
 sky130_fd_sc_hd__nor2_2 _18456_ (.A(_03885_),
    .B(_03888_),
    .Y(_03958_));
 sky130_fd_sc_hd__nand3b_2 _18457_ (.A_N(_03728_),
    .B(_03729_),
    .C(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__and2_4 _18458_ (.A(net766),
    .B(net839),
    .X(_03960_));
 sky130_fd_sc_hd__nor2_1 _18459_ (.A(net783),
    .B(_03757_),
    .Y(_03961_));
 sky130_fd_sc_hd__mux2_1 _18460_ (.A0(_03961_),
    .A1(\core.csr.traps.mcause.csrReadData[0] ),
    .S(net752),
    .X(_03962_));
 sky130_fd_sc_hd__o21a_1 _18461_ (.A1(_03957_),
    .A2(_03962_),
    .B1(net1935),
    .X(_01798_));
 sky130_fd_sc_hd__or3b_2 _18462_ (.A(net767),
    .B(_07469_),
    .C_N(_07502_),
    .X(_03963_));
 sky130_fd_sc_hd__or2_1 _18463_ (.A(net784),
    .B(_03761_),
    .X(_03964_));
 sky130_fd_sc_hd__o2bb2a_1 _18464_ (.A1_N(\core.csr.traps.mcause.csrReadData[1] ),
    .A2_N(net753),
    .B1(_03964_),
    .B2(net840),
    .X(_03965_));
 sky130_fd_sc_hd__a21oi_1 _18465_ (.A1(_03963_),
    .A2(_03965_),
    .B1(net1984),
    .Y(_01799_));
 sky130_fd_sc_hd__or2_1 _18466_ (.A(net783),
    .B(_03765_),
    .X(_03966_));
 sky130_fd_sc_hd__nor2_1 _18467_ (.A(net752),
    .B(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__a32o_1 _18468_ (.A1(net780),
    .A2(_07470_),
    .A3(net811),
    .B1(net752),
    .B2(\core.csr.traps.mcause.csrReadData[2] ),
    .X(_03968_));
 sky130_fd_sc_hd__o21a_1 _18469_ (.A1(_03967_),
    .A2(_03968_),
    .B1(net1931),
    .X(_01800_));
 sky130_fd_sc_hd__nor2_1 _18470_ (.A(net781),
    .B(_03769_),
    .Y(_03969_));
 sky130_fd_sc_hd__or2_1 _18471_ (.A(net781),
    .B(_03769_),
    .X(_03970_));
 sky130_fd_sc_hd__or2_1 _18472_ (.A(net766),
    .B(_07468_),
    .X(_03971_));
 sky130_fd_sc_hd__nand2_1 _18473_ (.A(_03970_),
    .B(net749),
    .Y(_03972_));
 sky130_fd_sc_hd__mux2_1 _18474_ (.A0(_03972_),
    .A1(\core.csr.traps.mcause.csrReadData[3] ),
    .S(net752),
    .X(_03973_));
 sky130_fd_sc_hd__a31o_1 _18475_ (.A1(net780),
    .A2(_07470_),
    .A3(net444),
    .B1(_03973_),
    .X(_03974_));
 sky130_fd_sc_hd__and2_1 _18476_ (.A(net1931),
    .B(_03974_),
    .X(_01801_));
 sky130_fd_sc_hd__or2_1 _18477_ (.A(net783),
    .B(_03773_),
    .X(_03975_));
 sky130_fd_sc_hd__o2bb2a_1 _18478_ (.A1_N(\core.csr.traps.mcause.csrReadData[4] ),
    .A2_N(net753),
    .B1(_03975_),
    .B2(net840),
    .X(_03976_));
 sky130_fd_sc_hd__nor2_1 _18479_ (.A(net1984),
    .B(_03976_),
    .Y(_01802_));
 sky130_fd_sc_hd__or2_2 _18480_ (.A(net781),
    .B(_03777_),
    .X(_03977_));
 sky130_fd_sc_hd__o2bb2a_1 _18481_ (.A1_N(\core.csr.traps.mcause.csrReadData[5] ),
    .A2_N(net753),
    .B1(_03977_),
    .B2(net840),
    .X(_03978_));
 sky130_fd_sc_hd__nor2_1 _18482_ (.A(net1980),
    .B(_03978_),
    .Y(_01803_));
 sky130_fd_sc_hd__or2_2 _18483_ (.A(net783),
    .B(_03781_),
    .X(_03979_));
 sky130_fd_sc_hd__o2bb2a_1 _18484_ (.A1_N(\core.csr.traps.mcause.csrReadData[6] ),
    .A2_N(net753),
    .B1(_03979_),
    .B2(net840),
    .X(_03980_));
 sky130_fd_sc_hd__nor2_1 _18485_ (.A(net1984),
    .B(_03980_),
    .Y(_01804_));
 sky130_fd_sc_hd__nor2_1 _18486_ (.A(net780),
    .B(_03785_),
    .Y(_03981_));
 sky130_fd_sc_hd__or2_1 _18487_ (.A(net778),
    .B(_03785_),
    .X(_03982_));
 sky130_fd_sc_hd__o2bb2a_1 _18488_ (.A1_N(\core.csr.traps.mcause.csrReadData[7] ),
    .A2_N(net753),
    .B1(_03982_),
    .B2(net841),
    .X(_03983_));
 sky130_fd_sc_hd__nor2_1 _18489_ (.A(net1980),
    .B(_03983_),
    .Y(_01805_));
 sky130_fd_sc_hd__or2_4 _18490_ (.A(net784),
    .B(_03789_),
    .X(_03984_));
 sky130_fd_sc_hd__o2bb2a_1 _18491_ (.A1_N(\core.csr.traps.mcause.csrReadData[8] ),
    .A2_N(net753),
    .B1(_03984_),
    .B2(net841),
    .X(_03985_));
 sky130_fd_sc_hd__nor2_1 _18492_ (.A(net1980),
    .B(_03985_),
    .Y(_01806_));
 sky130_fd_sc_hd__or2_2 _18493_ (.A(net778),
    .B(_03793_),
    .X(_03986_));
 sky130_fd_sc_hd__o2bb2a_1 _18494_ (.A1_N(\core.csr.traps.mcause.csrReadData[9] ),
    .A2_N(net752),
    .B1(_03986_),
    .B2(net840),
    .X(_03987_));
 sky130_fd_sc_hd__nor2_1 _18495_ (.A(net1980),
    .B(_03987_),
    .Y(_01807_));
 sky130_fd_sc_hd__or2_2 _18496_ (.A(net778),
    .B(_03797_),
    .X(_03988_));
 sky130_fd_sc_hd__o2bb2a_1 _18497_ (.A1_N(\core.csr.traps.mcause.csrReadData[10] ),
    .A2_N(net752),
    .B1(_03988_),
    .B2(net840),
    .X(_03989_));
 sky130_fd_sc_hd__nor2_1 _18498_ (.A(net1975),
    .B(_03989_),
    .Y(_01808_));
 sky130_fd_sc_hd__or2_1 _18499_ (.A(net777),
    .B(_03801_),
    .X(_03990_));
 sky130_fd_sc_hd__o2bb2a_1 _18500_ (.A1_N(\core.csr.traps.mcause.csrReadData[11] ),
    .A2_N(net752),
    .B1(_03990_),
    .B2(net840),
    .X(_03991_));
 sky130_fd_sc_hd__nor2_1 _18501_ (.A(net1975),
    .B(_03991_),
    .Y(_01809_));
 sky130_fd_sc_hd__or2_2 _18502_ (.A(net777),
    .B(_03805_),
    .X(_03992_));
 sky130_fd_sc_hd__o2bb2a_1 _18503_ (.A1_N(\core.csr.traps.mcause.csrReadData[12] ),
    .A2_N(net752),
    .B1(_03992_),
    .B2(net840),
    .X(_03993_));
 sky130_fd_sc_hd__nor2_1 _18504_ (.A(net1975),
    .B(_03993_),
    .Y(_01810_));
 sky130_fd_sc_hd__or2_2 _18505_ (.A(net779),
    .B(_03809_),
    .X(_03994_));
 sky130_fd_sc_hd__o2bb2a_1 _18506_ (.A1_N(\core.csr.traps.mcause.csrReadData[13] ),
    .A2_N(net752),
    .B1(_03994_),
    .B2(net840),
    .X(_03995_));
 sky130_fd_sc_hd__nor2_1 _18507_ (.A(net1971),
    .B(_03995_),
    .Y(_01811_));
 sky130_fd_sc_hd__or2_1 _18508_ (.A(net777),
    .B(_03813_),
    .X(_03996_));
 sky130_fd_sc_hd__o2bb2a_1 _18509_ (.A1_N(\core.csr.traps.mcause.csrReadData[14] ),
    .A2_N(net752),
    .B1(_03996_),
    .B2(net840),
    .X(_03997_));
 sky130_fd_sc_hd__nor2_1 _18510_ (.A(net1975),
    .B(_03997_),
    .Y(_01812_));
 sky130_fd_sc_hd__or2_1 _18511_ (.A(net775),
    .B(_03817_),
    .X(_03998_));
 sky130_fd_sc_hd__o2bb2a_1 _18512_ (.A1_N(\core.csr.traps.mcause.csrReadData[15] ),
    .A2_N(net751),
    .B1(_03998_),
    .B2(net839),
    .X(_03999_));
 sky130_fd_sc_hd__nor2_1 _18513_ (.A(net1971),
    .B(_03999_),
    .Y(_01813_));
 sky130_fd_sc_hd__or2_1 _18514_ (.A(net775),
    .B(_03821_),
    .X(_04000_));
 sky130_fd_sc_hd__o2bb2a_1 _18515_ (.A1_N(\core.csr.traps.mcause.csrReadData[16] ),
    .A2_N(net751),
    .B1(_04000_),
    .B2(net839),
    .X(_04001_));
 sky130_fd_sc_hd__nor2_1 _18516_ (.A(net1971),
    .B(_04001_),
    .Y(_01814_));
 sky130_fd_sc_hd__or2_1 _18517_ (.A(net775),
    .B(_03825_),
    .X(_04002_));
 sky130_fd_sc_hd__o2bb2a_1 _18518_ (.A1_N(\core.csr.traps.mcause.csrReadData[17] ),
    .A2_N(net751),
    .B1(_04002_),
    .B2(net839),
    .X(_04003_));
 sky130_fd_sc_hd__nor2_1 _18519_ (.A(net1971),
    .B(_04003_),
    .Y(_01815_));
 sky130_fd_sc_hd__or2_1 _18520_ (.A(net774),
    .B(_03829_),
    .X(_04004_));
 sky130_fd_sc_hd__o2bb2a_1 _18521_ (.A1_N(\core.csr.traps.mcause.csrReadData[18] ),
    .A2_N(net751),
    .B1(_04004_),
    .B2(net839),
    .X(_04005_));
 sky130_fd_sc_hd__nor2_1 _18522_ (.A(net1971),
    .B(_04005_),
    .Y(_01816_));
 sky130_fd_sc_hd__or2_1 _18523_ (.A(net774),
    .B(_03833_),
    .X(_04006_));
 sky130_fd_sc_hd__o2bb2a_1 _18524_ (.A1_N(\core.csr.traps.mcause.csrReadData[19] ),
    .A2_N(net751),
    .B1(_04006_),
    .B2(net839),
    .X(_04007_));
 sky130_fd_sc_hd__nor2_1 _18525_ (.A(net1966),
    .B(_04007_),
    .Y(_01817_));
 sky130_fd_sc_hd__or2_1 _18526_ (.A(net770),
    .B(_03837_),
    .X(_04008_));
 sky130_fd_sc_hd__o2bb2a_1 _18527_ (.A1_N(\core.csr.traps.mcause.csrReadData[20] ),
    .A2_N(net750),
    .B1(_04008_),
    .B2(net838),
    .X(_04009_));
 sky130_fd_sc_hd__nor2_1 _18528_ (.A(net1964),
    .B(_04009_),
    .Y(_01818_));
 sky130_fd_sc_hd__or2_2 _18529_ (.A(net769),
    .B(_03841_),
    .X(_04010_));
 sky130_fd_sc_hd__o2bb2a_1 _18530_ (.A1_N(\core.csr.traps.mcause.csrReadData[21] ),
    .A2_N(net750),
    .B1(_04010_),
    .B2(net838),
    .X(_04011_));
 sky130_fd_sc_hd__nor2_1 _18531_ (.A(net1962),
    .B(_04011_),
    .Y(_01819_));
 sky130_fd_sc_hd__or2_2 _18532_ (.A(net769),
    .B(_03845_),
    .X(_04012_));
 sky130_fd_sc_hd__o2bb2a_1 _18533_ (.A1_N(\core.csr.traps.mcause.csrReadData[22] ),
    .A2_N(net750),
    .B1(_04012_),
    .B2(net838),
    .X(_04013_));
 sky130_fd_sc_hd__nor2_1 _18534_ (.A(net1962),
    .B(_04013_),
    .Y(_01820_));
 sky130_fd_sc_hd__or2_2 _18535_ (.A(net769),
    .B(_03849_),
    .X(_04014_));
 sky130_fd_sc_hd__o2bb2a_1 _18536_ (.A1_N(\core.csr.traps.mcause.csrReadData[23] ),
    .A2_N(net750),
    .B1(_04014_),
    .B2(net838),
    .X(_04015_));
 sky130_fd_sc_hd__nor2_1 _18537_ (.A(net1962),
    .B(_04015_),
    .Y(_01821_));
 sky130_fd_sc_hd__or2_1 _18538_ (.A(net769),
    .B(_03853_),
    .X(_04016_));
 sky130_fd_sc_hd__o2bb2a_1 _18539_ (.A1_N(\core.csr.traps.mcause.csrReadData[24] ),
    .A2_N(net750),
    .B1(_04016_),
    .B2(net838),
    .X(_04017_));
 sky130_fd_sc_hd__nor2_1 _18540_ (.A(net1962),
    .B(_04017_),
    .Y(_01822_));
 sky130_fd_sc_hd__or2_1 _18541_ (.A(net773),
    .B(_03857_),
    .X(_04018_));
 sky130_fd_sc_hd__o2bb2a_1 _18542_ (.A1_N(\core.csr.traps.mcause.csrReadData[25] ),
    .A2_N(net750),
    .B1(_04018_),
    .B2(net838),
    .X(_04019_));
 sky130_fd_sc_hd__nor2_1 _18543_ (.A(net1965),
    .B(_04019_),
    .Y(_01823_));
 sky130_fd_sc_hd__or2_1 _18544_ (.A(net773),
    .B(_03861_),
    .X(_04020_));
 sky130_fd_sc_hd__o2bb2a_1 _18545_ (.A1_N(\core.csr.traps.mcause.csrReadData[26] ),
    .A2_N(net750),
    .B1(_04020_),
    .B2(net838),
    .X(_04021_));
 sky130_fd_sc_hd__nor2_1 _18546_ (.A(net1965),
    .B(_04021_),
    .Y(_01824_));
 sky130_fd_sc_hd__or2_1 _18547_ (.A(net773),
    .B(_03865_),
    .X(_04022_));
 sky130_fd_sc_hd__o2bb2a_1 _18548_ (.A1_N(\core.csr.traps.mcause.csrReadData[27] ),
    .A2_N(net751),
    .B1(_04022_),
    .B2(net839),
    .X(_04023_));
 sky130_fd_sc_hd__nor2_1 _18549_ (.A(net1966),
    .B(_04023_),
    .Y(_01825_));
 sky130_fd_sc_hd__or2_1 _18550_ (.A(net769),
    .B(_03869_),
    .X(_04024_));
 sky130_fd_sc_hd__o2bb2a_1 _18551_ (.A1_N(\core.csr.traps.mcause.csrReadData[28] ),
    .A2_N(net750),
    .B1(_04024_),
    .B2(net838),
    .X(_04025_));
 sky130_fd_sc_hd__nor2_1 _18552_ (.A(net1964),
    .B(_04025_),
    .Y(_01826_));
 sky130_fd_sc_hd__or2_1 _18553_ (.A(net773),
    .B(_03873_),
    .X(_04026_));
 sky130_fd_sc_hd__o2bb2a_1 _18554_ (.A1_N(\core.csr.traps.mcause.csrReadData[29] ),
    .A2_N(net750),
    .B1(_04026_),
    .B2(net838),
    .X(_04027_));
 sky130_fd_sc_hd__nor2_1 _18555_ (.A(net1965),
    .B(_04027_),
    .Y(_01827_));
 sky130_fd_sc_hd__or2_2 _18556_ (.A(net769),
    .B(_03877_),
    .X(_04028_));
 sky130_fd_sc_hd__o2bb2a_1 _18557_ (.A1_N(\core.csr.traps.mcause.csrReadData[30] ),
    .A2_N(net750),
    .B1(_04028_),
    .B2(net838),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_1 _18558_ (.A(net1963),
    .B(_04029_),
    .Y(_01828_));
 sky130_fd_sc_hd__nand2_1 _18559_ (.A(\core.csr.traps.mcause.csrReadData[31] ),
    .B(net751),
    .Y(_04030_));
 sky130_fd_sc_hd__or2_1 _18560_ (.A(net773),
    .B(_03881_),
    .X(_04031_));
 sky130_fd_sc_hd__o211a_1 _18561_ (.A1(net751),
    .A2(_04031_),
    .B1(_04030_),
    .C1(net748),
    .X(_04032_));
 sky130_fd_sc_hd__nor2_1 _18562_ (.A(net1966),
    .B(_04032_),
    .Y(_01829_));
 sky130_fd_sc_hd__or3_4 _18563_ (.A(_03730_),
    .B(_03885_),
    .C(_03888_),
    .X(_04033_));
 sky130_fd_sc_hd__inv_2 _18564_ (.A(net891),
    .Y(_04034_));
 sky130_fd_sc_hd__nor2_8 _18565_ (.A(net783),
    .B(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hd__a22o_1 _18566_ (.A1(net450),
    .A2(net783),
    .B1(_03961_),
    .B2(_04034_),
    .X(_04036_));
 sky130_fd_sc_hd__a21oi_1 _18567_ (.A1(\core.csr.trapReturnVector[0] ),
    .A2(net763),
    .B1(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__nor2_1 _18568_ (.A(net1984),
    .B(_04037_),
    .Y(_01830_));
 sky130_fd_sc_hd__nand2_1 _18569_ (.A(\core.csr.trapReturnVector[1] ),
    .B(net763),
    .Y(_04038_));
 sky130_fd_sc_hd__nand2_2 _18570_ (.A(net461),
    .B(net783),
    .Y(_04039_));
 sky130_fd_sc_hd__o211a_1 _18571_ (.A1(_03964_),
    .A2(net891),
    .B1(_04038_),
    .C1(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__nor2_1 _18572_ (.A(net1984),
    .B(_04040_),
    .Y(_01831_));
 sky130_fd_sc_hd__nand2_1 _18573_ (.A(\core.csr.trapReturnVector[2] ),
    .B(net764),
    .Y(_04041_));
 sky130_fd_sc_hd__nand2_1 _18574_ (.A(net472),
    .B(net781),
    .Y(_04042_));
 sky130_fd_sc_hd__o211a_1 _18575_ (.A1(_03966_),
    .A2(net890),
    .B1(_04041_),
    .C1(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__nor2_1 _18576_ (.A(net1984),
    .B(_04043_),
    .Y(_01832_));
 sky130_fd_sc_hd__nand2_1 _18577_ (.A(\core.csr.trapReturnVector[3] ),
    .B(net764),
    .Y(_04044_));
 sky130_fd_sc_hd__o2bb2a_1 _18578_ (.A1_N(net475),
    .A2_N(net780),
    .B1(_03970_),
    .B2(net891),
    .X(_04045_));
 sky130_fd_sc_hd__a21oi_1 _18579_ (.A1(_04044_),
    .A2(_04045_),
    .B1(net1980),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_1 _18580_ (.A(\core.csr.trapReturnVector[4] ),
    .B(net764),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_2 _18581_ (.A(net476),
    .B(net781),
    .Y(_04047_));
 sky130_fd_sc_hd__o211a_1 _18582_ (.A1(_03975_),
    .A2(net891),
    .B1(_04046_),
    .C1(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__nor2_1 _18583_ (.A(net1984),
    .B(_04048_),
    .Y(_01834_));
 sky130_fd_sc_hd__nand2_1 _18584_ (.A(\core.csr.trapReturnVector[5] ),
    .B(net764),
    .Y(_04049_));
 sky130_fd_sc_hd__nand2_1 _18585_ (.A(net477),
    .B(net780),
    .Y(_04050_));
 sky130_fd_sc_hd__o211a_1 _18586_ (.A1(_03977_),
    .A2(net890),
    .B1(_04049_),
    .C1(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__nor2_1 _18587_ (.A(net1983),
    .B(_04051_),
    .Y(_01835_));
 sky130_fd_sc_hd__nand2_1 _18588_ (.A(\core.csr.trapReturnVector[6] ),
    .B(net763),
    .Y(_04052_));
 sky130_fd_sc_hd__nand2_2 _18589_ (.A(net478),
    .B(net780),
    .Y(_04053_));
 sky130_fd_sc_hd__o211a_1 _18590_ (.A1(_03979_),
    .A2(net890),
    .B1(_04052_),
    .C1(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__nor2_1 _18591_ (.A(net1984),
    .B(_04054_),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_1 _18592_ (.A(\core.csr.trapReturnVector[7] ),
    .B(net764),
    .Y(_04055_));
 sky130_fd_sc_hd__o22a_1 _18593_ (.A1(_04406_),
    .A2(net768),
    .B1(_03982_),
    .B2(net891),
    .X(_04056_));
 sky130_fd_sc_hd__a21oi_1 _18594_ (.A1(_04055_),
    .A2(_04056_),
    .B1(net1980),
    .Y(_01837_));
 sky130_fd_sc_hd__nand2_1 _18595_ (.A(\core.csr.trapReturnVector[8] ),
    .B(net763),
    .Y(_04057_));
 sky130_fd_sc_hd__nand2_1 _18596_ (.A(net480),
    .B(net778),
    .Y(_04058_));
 sky130_fd_sc_hd__o211a_1 _18597_ (.A1(_03984_),
    .A2(net890),
    .B1(_04057_),
    .C1(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__nor2_1 _18598_ (.A(net1980),
    .B(_04059_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2_1 _18599_ (.A(\core.csr.trapReturnVector[9] ),
    .B(net763),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2_1 _18600_ (.A(net481),
    .B(net778),
    .Y(_04061_));
 sky130_fd_sc_hd__o211a_1 _18601_ (.A1(_03986_),
    .A2(net890),
    .B1(_04060_),
    .C1(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__nor2_1 _18602_ (.A(net1975),
    .B(_04062_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _18603_ (.A(\core.csr.trapReturnVector[10] ),
    .B(net763),
    .Y(_04063_));
 sky130_fd_sc_hd__nand2_1 _18604_ (.A(net451),
    .B(net778),
    .Y(_04064_));
 sky130_fd_sc_hd__o211a_1 _18605_ (.A1(_03988_),
    .A2(net890),
    .B1(_04063_),
    .C1(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__nor2_1 _18606_ (.A(net1978),
    .B(_04065_),
    .Y(_01840_));
 sky130_fd_sc_hd__nand2_1 _18607_ (.A(\core.csr.trapReturnVector[11] ),
    .B(net763),
    .Y(_04066_));
 sky130_fd_sc_hd__nand2_1 _18608_ (.A(net452),
    .B(net777),
    .Y(_04067_));
 sky130_fd_sc_hd__o211a_1 _18609_ (.A1(_03990_),
    .A2(net890),
    .B1(_04066_),
    .C1(_04067_),
    .X(_04068_));
 sky130_fd_sc_hd__nor2_1 _18610_ (.A(net1978),
    .B(_04068_),
    .Y(_01841_));
 sky130_fd_sc_hd__nand2_1 _18611_ (.A(\core.csr.trapReturnVector[12] ),
    .B(net763),
    .Y(_04069_));
 sky130_fd_sc_hd__nand2_1 _18612_ (.A(net453),
    .B(net777),
    .Y(_04070_));
 sky130_fd_sc_hd__o211a_1 _18613_ (.A1(_03992_),
    .A2(net890),
    .B1(_04069_),
    .C1(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__nor2_1 _18614_ (.A(net1975),
    .B(_04071_),
    .Y(_01842_));
 sky130_fd_sc_hd__nand2_1 _18615_ (.A(\core.csr.trapReturnVector[13] ),
    .B(net763),
    .Y(_04072_));
 sky130_fd_sc_hd__nand2_1 _18616_ (.A(net454),
    .B(net779),
    .Y(_04073_));
 sky130_fd_sc_hd__o211a_1 _18617_ (.A1(_03994_),
    .A2(net890),
    .B1(_04072_),
    .C1(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__nor2_1 _18618_ (.A(net1975),
    .B(_04074_),
    .Y(_01843_));
 sky130_fd_sc_hd__nand2_1 _18619_ (.A(\core.csr.trapReturnVector[14] ),
    .B(net763),
    .Y(_04075_));
 sky130_fd_sc_hd__nand2_1 _18620_ (.A(net455),
    .B(net775),
    .Y(_04076_));
 sky130_fd_sc_hd__o211a_1 _18621_ (.A1(_03996_),
    .A2(net890),
    .B1(_04075_),
    .C1(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__nor2_1 _18622_ (.A(net1975),
    .B(_04077_),
    .Y(_01844_));
 sky130_fd_sc_hd__nand2_1 _18623_ (.A(\core.csr.trapReturnVector[15] ),
    .B(net762),
    .Y(_04078_));
 sky130_fd_sc_hd__nand2_1 _18624_ (.A(net456),
    .B(net775),
    .Y(_04079_));
 sky130_fd_sc_hd__o211a_1 _18625_ (.A1(_03998_),
    .A2(net889),
    .B1(_04078_),
    .C1(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__nor2_1 _18626_ (.A(net1974),
    .B(_04080_),
    .Y(_01845_));
 sky130_fd_sc_hd__nand2_1 _18627_ (.A(\core.csr.trapReturnVector[16] ),
    .B(net762),
    .Y(_04081_));
 sky130_fd_sc_hd__nand2_1 _18628_ (.A(net457),
    .B(net775),
    .Y(_04082_));
 sky130_fd_sc_hd__o211a_1 _18629_ (.A1(_04000_),
    .A2(net889),
    .B1(_04081_),
    .C1(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__nor2_1 _18630_ (.A(net1974),
    .B(_04083_),
    .Y(_01846_));
 sky130_fd_sc_hd__nand2_1 _18631_ (.A(\core.csr.trapReturnVector[17] ),
    .B(net762),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_1 _18632_ (.A(net458),
    .B(net774),
    .Y(_04085_));
 sky130_fd_sc_hd__o211a_1 _18633_ (.A1(_04002_),
    .A2(net889),
    .B1(_04084_),
    .C1(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__nor2_1 _18634_ (.A(net1971),
    .B(_04086_),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2_1 _18635_ (.A(\core.csr.trapReturnVector[18] ),
    .B(net762),
    .Y(_04087_));
 sky130_fd_sc_hd__nand2_1 _18636_ (.A(net459),
    .B(net774),
    .Y(_04088_));
 sky130_fd_sc_hd__o211a_1 _18637_ (.A1(_04004_),
    .A2(net889),
    .B1(_04087_),
    .C1(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__nor2_1 _18638_ (.A(net1971),
    .B(_04089_),
    .Y(_01848_));
 sky130_fd_sc_hd__nand2_1 _18639_ (.A(\core.csr.trapReturnVector[19] ),
    .B(net762),
    .Y(_04090_));
 sky130_fd_sc_hd__nand2_1 _18640_ (.A(net460),
    .B(net774),
    .Y(_04091_));
 sky130_fd_sc_hd__o211a_1 _18641_ (.A1(_04006_),
    .A2(net889),
    .B1(_04090_),
    .C1(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__nor2_1 _18642_ (.A(net1971),
    .B(_04092_),
    .Y(_01849_));
 sky130_fd_sc_hd__nand2_1 _18643_ (.A(\core.csr.trapReturnVector[20] ),
    .B(net761),
    .Y(_04093_));
 sky130_fd_sc_hd__o2bb2a_1 _18644_ (.A1_N(net462),
    .A2_N(net776),
    .B1(_04008_),
    .B2(net888),
    .X(_04094_));
 sky130_fd_sc_hd__a21oi_1 _18645_ (.A1(_04093_),
    .A2(_04094_),
    .B1(net1965),
    .Y(_01850_));
 sky130_fd_sc_hd__nand2_1 _18646_ (.A(\core.csr.trapReturnVector[21] ),
    .B(net761),
    .Y(_04095_));
 sky130_fd_sc_hd__nand2_1 _18647_ (.A(net463),
    .B(net770),
    .Y(_04096_));
 sky130_fd_sc_hd__o211a_1 _18648_ (.A1(_04010_),
    .A2(net888),
    .B1(_04095_),
    .C1(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__nor2_1 _18649_ (.A(net1963),
    .B(_04097_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand2_1 _18650_ (.A(\core.csr.trapReturnVector[22] ),
    .B(net761),
    .Y(_04098_));
 sky130_fd_sc_hd__nand2_1 _18651_ (.A(net464),
    .B(net769),
    .Y(_04099_));
 sky130_fd_sc_hd__o211a_1 _18652_ (.A1(_04012_),
    .A2(net888),
    .B1(_04098_),
    .C1(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__nor2_1 _18653_ (.A(net1964),
    .B(_04100_),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _18654_ (.A(\core.csr.trapReturnVector[23] ),
    .B(net761),
    .Y(_04101_));
 sky130_fd_sc_hd__nand2_1 _18655_ (.A(net465),
    .B(net770),
    .Y(_04102_));
 sky130_fd_sc_hd__o211a_1 _18656_ (.A1(_04014_),
    .A2(net888),
    .B1(_04101_),
    .C1(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__nor2_1 _18657_ (.A(net1964),
    .B(_04103_),
    .Y(_01853_));
 sky130_fd_sc_hd__nand2_1 _18658_ (.A(\core.csr.trapReturnVector[24] ),
    .B(net761),
    .Y(_04104_));
 sky130_fd_sc_hd__nand2_1 _18659_ (.A(net466),
    .B(net770),
    .Y(_04105_));
 sky130_fd_sc_hd__o211a_1 _18660_ (.A1(_04016_),
    .A2(net888),
    .B1(_04104_),
    .C1(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__nor2_1 _18661_ (.A(net1962),
    .B(_04106_),
    .Y(_01854_));
 sky130_fd_sc_hd__nand2_1 _18662_ (.A(\core.csr.trapReturnVector[25] ),
    .B(net762),
    .Y(_04107_));
 sky130_fd_sc_hd__nand2_1 _18663_ (.A(net467),
    .B(net771),
    .Y(_04108_));
 sky130_fd_sc_hd__o211a_1 _18664_ (.A1(_04018_),
    .A2(net889),
    .B1(_04107_),
    .C1(_04108_),
    .X(_04109_));
 sky130_fd_sc_hd__nor2_1 _18665_ (.A(net1965),
    .B(_04109_),
    .Y(_01855_));
 sky130_fd_sc_hd__nand2_1 _18666_ (.A(\core.csr.trapReturnVector[26] ),
    .B(net761),
    .Y(_04110_));
 sky130_fd_sc_hd__nand2_1 _18667_ (.A(net468),
    .B(net771),
    .Y(_04111_));
 sky130_fd_sc_hd__o211a_1 _18668_ (.A1(_04020_),
    .A2(net888),
    .B1(_04110_),
    .C1(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__nor2_1 _18669_ (.A(net1965),
    .B(_04112_),
    .Y(_01856_));
 sky130_fd_sc_hd__nand2_1 _18670_ (.A(\core.csr.trapReturnVector[27] ),
    .B(net761),
    .Y(_04113_));
 sky130_fd_sc_hd__nand2_1 _18671_ (.A(net469),
    .B(net774),
    .Y(_04114_));
 sky130_fd_sc_hd__o211a_1 _18672_ (.A1(_04022_),
    .A2(net888),
    .B1(_04113_),
    .C1(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__nor2_1 _18673_ (.A(net1966),
    .B(_04115_),
    .Y(_01857_));
 sky130_fd_sc_hd__nand2_1 _18674_ (.A(\core.csr.trapReturnVector[28] ),
    .B(net761),
    .Y(_04116_));
 sky130_fd_sc_hd__nand2_1 _18675_ (.A(net470),
    .B(net770),
    .Y(_04117_));
 sky130_fd_sc_hd__o211a_1 _18676_ (.A1(_04024_),
    .A2(net888),
    .B1(_04116_),
    .C1(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__nor2_1 _18677_ (.A(net1964),
    .B(_04118_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand2_1 _18678_ (.A(\core.csr.trapReturnVector[29] ),
    .B(net761),
    .Y(_04119_));
 sky130_fd_sc_hd__nand2_1 _18679_ (.A(net471),
    .B(net772),
    .Y(_04120_));
 sky130_fd_sc_hd__o211a_1 _18680_ (.A1(_04026_),
    .A2(net888),
    .B1(_04119_),
    .C1(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__nor2_1 _18681_ (.A(net1965),
    .B(_04121_),
    .Y(_01859_));
 sky130_fd_sc_hd__nand2_1 _18682_ (.A(\core.csr.trapReturnVector[30] ),
    .B(net761),
    .Y(_04122_));
 sky130_fd_sc_hd__nand2_1 _18683_ (.A(net473),
    .B(net770),
    .Y(_04123_));
 sky130_fd_sc_hd__o211a_1 _18684_ (.A1(_04028_),
    .A2(net888),
    .B1(_04122_),
    .C1(_04123_),
    .X(_04124_));
 sky130_fd_sc_hd__nor2_1 _18685_ (.A(net1963),
    .B(_04124_),
    .Y(_01860_));
 sky130_fd_sc_hd__nand2_1 _18686_ (.A(\core.csr.trapReturnVector[31] ),
    .B(net762),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _18687_ (.A(net474),
    .B(net772),
    .Y(_04126_));
 sky130_fd_sc_hd__o211a_1 _18688_ (.A1(_04031_),
    .A2(net889),
    .B1(_04125_),
    .C1(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__nor2_1 _18689_ (.A(net1966),
    .B(_04127_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_8 _18690_ (.A(_03753_),
    .B(_03923_),
    .Y(_04128_));
 sky130_fd_sc_hd__mux2_1 _18691_ (.A0(\core.csr.traps.mtvec.csrReadData[0] ),
    .A1(_03758_),
    .S(net837),
    .X(_04129_));
 sky130_fd_sc_hd__and2_1 _18692_ (.A(net1953),
    .B(_04129_),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _18693_ (.A0(\core.csr.traps.mtvec.csrReadData[1] ),
    .A1(_03762_),
    .S(net837),
    .X(_04130_));
 sky130_fd_sc_hd__and2_1 _18694_ (.A(net1935),
    .B(_04130_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _18695_ (.A0(_04394_),
    .A1(_03765_),
    .S(net837),
    .X(_04131_));
 sky130_fd_sc_hd__nor2_1 _18696_ (.A(net1984),
    .B(_04131_),
    .Y(_01864_));
 sky130_fd_sc_hd__mux2_1 _18697_ (.A0(\core.csr.traps.mtvec.csrReadData[3] ),
    .A1(_03770_),
    .S(net836),
    .X(_04132_));
 sky130_fd_sc_hd__and2_1 _18698_ (.A(net1934),
    .B(_04132_),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _18699_ (.A0(\core.csr.traps.mtvec.csrReadData[4] ),
    .A1(_03774_),
    .S(net837),
    .X(_04133_));
 sky130_fd_sc_hd__and2_1 _18700_ (.A(net1936),
    .B(_04133_),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _18701_ (.A0(\core.csr.traps.mtvec.csrReadData[5] ),
    .A1(_03778_),
    .S(net836),
    .X(_04134_));
 sky130_fd_sc_hd__and2_1 _18702_ (.A(net1933),
    .B(_04134_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _18703_ (.A0(_04393_),
    .A1(_03781_),
    .S(net836),
    .X(_04135_));
 sky130_fd_sc_hd__nor2_1 _18704_ (.A(net1996),
    .B(_04135_),
    .Y(_01868_));
 sky130_fd_sc_hd__mux2_1 _18705_ (.A0(\core.csr.traps.mtvec.csrReadData[7] ),
    .A1(_03786_),
    .S(net836),
    .X(_04136_));
 sky130_fd_sc_hd__and2_1 _18706_ (.A(net1932),
    .B(_04136_),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _18707_ (.A0(\core.csr.traps.mtvec.csrReadData[8] ),
    .A1(_03790_),
    .S(net837),
    .X(_04137_));
 sky130_fd_sc_hd__and2_1 _18708_ (.A(net1955),
    .B(_04137_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _18709_ (.A0(\core.csr.traps.mtvec.csrReadData[9] ),
    .A1(_03794_),
    .S(net836),
    .X(_04138_));
 sky130_fd_sc_hd__and2_1 _18710_ (.A(net1930),
    .B(_04138_),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _18711_ (.A0(\core.csr.traps.mtvec.csrReadData[10] ),
    .A1(_03798_),
    .S(net836),
    .X(_04139_));
 sky130_fd_sc_hd__and2_1 _18712_ (.A(net1932),
    .B(_04139_),
    .X(_01872_));
 sky130_fd_sc_hd__mux2_1 _18713_ (.A0(\core.csr.traps.mtvec.csrReadData[11] ),
    .A1(_03802_),
    .S(net836),
    .X(_04140_));
 sky130_fd_sc_hd__and2_1 _18714_ (.A(net1914),
    .B(_04140_),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _18715_ (.A0(\core.csr.traps.mtvec.csrReadData[12] ),
    .A1(_03806_),
    .S(net836),
    .X(_04141_));
 sky130_fd_sc_hd__and2_1 _18716_ (.A(net1916),
    .B(_04141_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _18717_ (.A0(\core.csr.traps.mtvec.csrReadData[13] ),
    .A1(_03810_),
    .S(net836),
    .X(_04142_));
 sky130_fd_sc_hd__and2_1 _18718_ (.A(net1917),
    .B(_04142_),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _18719_ (.A0(\core.csr.traps.mtvec.csrReadData[14] ),
    .A1(_03814_),
    .S(net836),
    .X(_04143_));
 sky130_fd_sc_hd__and2_1 _18720_ (.A(net1916),
    .B(_04143_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _18721_ (.A0(\core.csr.traps.mtvec.csrReadData[15] ),
    .A1(_03818_),
    .S(net835),
    .X(_04144_));
 sky130_fd_sc_hd__and2_1 _18722_ (.A(net1912),
    .B(_04144_),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _18723_ (.A0(\core.csr.traps.mtvec.csrReadData[16] ),
    .A1(_03822_),
    .S(net835),
    .X(_04145_));
 sky130_fd_sc_hd__and2_1 _18724_ (.A(net1912),
    .B(_04145_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _18725_ (.A0(\core.csr.traps.mtvec.csrReadData[17] ),
    .A1(_03826_),
    .S(net835),
    .X(_04146_));
 sky130_fd_sc_hd__and2_1 _18726_ (.A(net1918),
    .B(_04146_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _18727_ (.A0(\core.csr.traps.mtvec.csrReadData[18] ),
    .A1(_03830_),
    .S(net835),
    .X(_04147_));
 sky130_fd_sc_hd__and2_1 _18728_ (.A(net1911),
    .B(_04147_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _18729_ (.A0(\core.csr.traps.mtvec.csrReadData[19] ),
    .A1(_03834_),
    .S(net835),
    .X(_04148_));
 sky130_fd_sc_hd__and2_1 _18730_ (.A(net1903),
    .B(_04148_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _18731_ (.A0(\core.csr.traps.mtvec.csrReadData[20] ),
    .A1(_03838_),
    .S(net834),
    .X(_04149_));
 sky130_fd_sc_hd__and2_1 _18732_ (.A(net1897),
    .B(_04149_),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _18733_ (.A0(\core.csr.traps.mtvec.csrReadData[21] ),
    .A1(_03842_),
    .S(net834),
    .X(_04150_));
 sky130_fd_sc_hd__and2_1 _18734_ (.A(net1896),
    .B(_04150_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _18735_ (.A0(\core.csr.traps.mtvec.csrReadData[22] ),
    .A1(_03846_),
    .S(net834),
    .X(_04151_));
 sky130_fd_sc_hd__and2_1 _18736_ (.A(net1898),
    .B(_04151_),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _18737_ (.A0(\core.csr.traps.mtvec.csrReadData[23] ),
    .A1(_03850_),
    .S(net834),
    .X(_04152_));
 sky130_fd_sc_hd__and2_1 _18738_ (.A(net1897),
    .B(_04152_),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _18739_ (.A0(\core.csr.traps.mtvec.csrReadData[24] ),
    .A1(_03854_),
    .S(net834),
    .X(_04153_));
 sky130_fd_sc_hd__and2_1 _18740_ (.A(net1895),
    .B(_04153_),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _18741_ (.A0(\core.csr.traps.mtvec.csrReadData[25] ),
    .A1(_03858_),
    .S(net834),
    .X(_04154_));
 sky130_fd_sc_hd__and2_1 _18742_ (.A(net1897),
    .B(_04154_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _18743_ (.A0(\core.csr.traps.mtvec.csrReadData[26] ),
    .A1(_03862_),
    .S(net834),
    .X(_04155_));
 sky130_fd_sc_hd__and2_1 _18744_ (.A(net1901),
    .B(_04155_),
    .X(_01888_));
 sky130_fd_sc_hd__mux2_1 _18745_ (.A0(\core.csr.traps.mtvec.csrReadData[27] ),
    .A1(_03866_),
    .S(net835),
    .X(_04156_));
 sky130_fd_sc_hd__and2_1 _18746_ (.A(net1901),
    .B(_04156_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _18747_ (.A0(\core.csr.traps.mtvec.csrReadData[28] ),
    .A1(_03870_),
    .S(net834),
    .X(_04157_));
 sky130_fd_sc_hd__and2_1 _18748_ (.A(net1897),
    .B(_04157_),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _18749_ (.A0(\core.csr.traps.mtvec.csrReadData[29] ),
    .A1(_03874_),
    .S(net835),
    .X(_04158_));
 sky130_fd_sc_hd__and2_1 _18750_ (.A(net1902),
    .B(_04158_),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _18751_ (.A0(\core.csr.traps.mtvec.csrReadData[30] ),
    .A1(_03878_),
    .S(net834),
    .X(_04159_));
 sky130_fd_sc_hd__and2_1 _18752_ (.A(net1894),
    .B(_04159_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _18753_ (.A0(\core.csr.traps.mtvec.csrReadData[31] ),
    .A1(_03882_),
    .S(net834),
    .X(_04160_));
 sky130_fd_sc_hd__and2_1 _18754_ (.A(net1902),
    .B(_04160_),
    .X(_01893_));
 sky130_fd_sc_hd__nor2_2 _18755_ (.A(_03887_),
    .B(_03923_),
    .Y(_04161_));
 sky130_fd_sc_hd__nor2_1 _18756_ (.A(net781),
    .B(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hd__a22o_1 _18757_ (.A1(net1774),
    .A2(_07422_),
    .B1(_03969_),
    .B2(_04161_),
    .X(_04163_));
 sky130_fd_sc_hd__a21o_1 _18758_ (.A1(\core.csr.traps.machineInterruptEnable ),
    .A2(_04162_),
    .B1(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__o311a_1 _18759_ (.A1(\core.csr.traps.machinePreviousInterruptEnable ),
    .A2(net1762),
    .A3(_07433_),
    .B1(_04164_),
    .C1(net1931),
    .X(_01894_));
 sky130_fd_sc_hd__and2_4 _18760_ (.A(\core.csr.traps.machineInterruptEnable ),
    .B(net781),
    .X(_04165_));
 sky130_fd_sc_hd__a21o_1 _18761_ (.A1(_03981_),
    .A2(_04161_),
    .B1(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__a21o_1 _18762_ (.A1(\core.csr.traps.machinePreviousInterruptEnable ),
    .A2(_04162_),
    .B1(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__o211a_1 _18763_ (.A1(net1762),
    .A2(_07433_),
    .B1(_04167_),
    .C1(net1931),
    .X(_01895_));
 sky130_fd_sc_hd__o2bb2a_1 _18764_ (.A1_N(\core.csr.currentInstruction[0] ),
    .A2_N(net1019),
    .B1(_07504_),
    .B2(net831),
    .X(_04168_));
 sky130_fd_sc_hd__or4_4 _18765_ (.A(net1730),
    .B(net1861),
    .C(_07416_),
    .D(_07501_),
    .X(_04169_));
 sky130_fd_sc_hd__o21ai_1 _18766_ (.A1(\core.csr.instruction_memoryAddress[1] ),
    .A2(_04168_),
    .B1(net1163),
    .Y(_04170_));
 sky130_fd_sc_hd__or2_1 _18767_ (.A(net766),
    .B(net1076),
    .X(_04171_));
 sky130_fd_sc_hd__o22a_1 _18768_ (.A1(net450),
    .A2(net1163),
    .B1(_04170_),
    .B2(\core.csr.instruction_memoryAddress[0] ),
    .X(_04172_));
 sky130_fd_sc_hd__a31oi_4 _18769_ (.A1(_03728_),
    .A2(_03729_),
    .A3(_03958_),
    .B1(net783),
    .Y(_04173_));
 sky130_fd_sc_hd__mux2_1 _18770_ (.A0(_03961_),
    .A1(\core.csr.traps.mtval.csrReadData[0] ),
    .S(net760),
    .X(_04174_));
 sky130_fd_sc_hd__a21oi_1 _18771_ (.A1(net783),
    .A2(_04172_),
    .B1(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__nor2_1 _18772_ (.A(net1988),
    .B(_04175_),
    .Y(_01896_));
 sky130_fd_sc_hd__o2bb2a_1 _18773_ (.A1_N(\core.csr.currentInstruction[1] ),
    .A2_N(net1019),
    .B1(_07504_),
    .B2(_07475_),
    .X(_04176_));
 sky130_fd_sc_hd__o21ai_1 _18774_ (.A1(\core.csr.instruction_memoryAddress[0] ),
    .A2(_04176_),
    .B1(net1163),
    .Y(_04177_));
 sky130_fd_sc_hd__a2bb2o_2 _18775_ (.A1_N(\core.csr.instruction_memoryAddress[1] ),
    .A2_N(_04177_),
    .B1(net745),
    .B2(_04039_),
    .X(_04178_));
 sky130_fd_sc_hd__mux2_1 _18776_ (.A0(_03964_),
    .A1(_04392_),
    .S(net760),
    .X(_04179_));
 sky130_fd_sc_hd__a21oi_1 _18777_ (.A1(_04178_),
    .A2(_04179_),
    .B1(net1988),
    .Y(_01897_));
 sky130_fd_sc_hd__a221o_1 _18778_ (.A1(\core.csr.currentInstruction[2] ),
    .A2(net1019),
    .B1(net811),
    .B2(_08382_),
    .C1(net1645),
    .X(_04180_));
 sky130_fd_sc_hd__o21ai_2 _18779_ (.A1(\core.csr.instruction_memoryAddress[2] ),
    .A2(net1650),
    .B1(_04180_),
    .Y(_04181_));
 sky130_fd_sc_hd__a22o_1 _18780_ (.A1(_04042_),
    .A2(net745),
    .B1(_04181_),
    .B2(net1163),
    .X(_04182_));
 sky130_fd_sc_hd__nand2_1 _18781_ (.A(\core.csr.traps.mtval.csrReadData[2] ),
    .B(net759),
    .Y(_04183_));
 sky130_fd_sc_hd__o211a_1 _18782_ (.A1(_03966_),
    .A2(net760),
    .B1(_04182_),
    .C1(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__nor2_1 _18783_ (.A(net1984),
    .B(_04184_),
    .Y(_01898_));
 sky130_fd_sc_hd__or2_1 _18784_ (.A(\core.csr.instruction_memoryAddress[3] ),
    .B(net1649),
    .X(_04185_));
 sky130_fd_sc_hd__a221o_1 _18785_ (.A1(\core.csr.currentInstruction[3] ),
    .A2(net1020),
    .B1(net811),
    .B2(_08395_),
    .C1(net1646),
    .X(_04186_));
 sky130_fd_sc_hd__a21o_1 _18786_ (.A1(_04185_),
    .A2(_04186_),
    .B1(net1077),
    .X(_04187_));
 sky130_fd_sc_hd__o211a_1 _18787_ (.A1(net475),
    .A2(net1163),
    .B1(_04187_),
    .C1(net780),
    .X(_04188_));
 sky130_fd_sc_hd__mux2_1 _18788_ (.A0(_03969_),
    .A1(\core.csr.traps.mtval.csrReadData[3] ),
    .S(net759),
    .X(_04189_));
 sky130_fd_sc_hd__o21a_1 _18789_ (.A1(_04188_),
    .A2(_04189_),
    .B1(net1931),
    .X(_01899_));
 sky130_fd_sc_hd__o2bb2a_1 _18790_ (.A1_N(\core.csr.currentInstruction[4] ),
    .A2_N(net1020),
    .B1(_07504_),
    .B2(_08421_),
    .X(_04190_));
 sky130_fd_sc_hd__mux2_2 _18791_ (.A0(_04408_),
    .A1(_04190_),
    .S(net1650),
    .X(_04191_));
 sky130_fd_sc_hd__a22o_1 _18792_ (.A1(_04047_),
    .A2(net745),
    .B1(_04191_),
    .B2(net1163),
    .X(_04192_));
 sky130_fd_sc_hd__nand2_1 _18793_ (.A(\core.csr.traps.mtval.csrReadData[4] ),
    .B(net760),
    .Y(_04193_));
 sky130_fd_sc_hd__o211a_1 _18794_ (.A1(_03975_),
    .A2(net759),
    .B1(_04192_),
    .C1(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__nor2_1 _18795_ (.A(net1987),
    .B(_04194_),
    .Y(_01900_));
 sky130_fd_sc_hd__o2bb2a_1 _18796_ (.A1_N(\core.csr.currentInstruction[5] ),
    .A2_N(net1020),
    .B1(_07504_),
    .B2(_08435_),
    .X(_04195_));
 sky130_fd_sc_hd__mux2_1 _18797_ (.A0(_04407_),
    .A1(_04195_),
    .S(net1649),
    .X(_04196_));
 sky130_fd_sc_hd__a22o_1 _18798_ (.A1(_04050_),
    .A2(net746),
    .B1(_04196_),
    .B2(net1163),
    .X(_04197_));
 sky130_fd_sc_hd__nand2_1 _18799_ (.A(\core.csr.traps.mtval.csrReadData[5] ),
    .B(net759),
    .Y(_04198_));
 sky130_fd_sc_hd__o211a_1 _18800_ (.A1(_03977_),
    .A2(net759),
    .B1(_04197_),
    .C1(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__nor2_1 _18801_ (.A(net1982),
    .B(_04199_),
    .Y(_01901_));
 sky130_fd_sc_hd__a22o_1 _18802_ (.A1(\core.csr.currentInstruction[6] ),
    .A2(net1019),
    .B1(net811),
    .B2(_08437_),
    .X(_04200_));
 sky130_fd_sc_hd__nand2_1 _18803_ (.A(net1650),
    .B(_04200_),
    .Y(_04201_));
 sky130_fd_sc_hd__a21oi_1 _18804_ (.A1(\core.csr.instruction_memoryAddress[6] ),
    .A2(net1646),
    .B1(net1077),
    .Y(_04202_));
 sky130_fd_sc_hd__a22o_2 _18805_ (.A1(_04053_),
    .A2(net746),
    .B1(_04201_),
    .B2(_04202_),
    .X(_04203_));
 sky130_fd_sc_hd__nand2_1 _18806_ (.A(\core.csr.traps.mtval.csrReadData[6] ),
    .B(net759),
    .Y(_04204_));
 sky130_fd_sc_hd__o211a_1 _18807_ (.A1(_03979_),
    .A2(net759),
    .B1(_04203_),
    .C1(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__nor2_1 _18808_ (.A(net1988),
    .B(_04205_),
    .Y(_01902_));
 sky130_fd_sc_hd__a22o_1 _18809_ (.A1(\core.csr.currentInstruction[7] ),
    .A2(net1019),
    .B1(net811),
    .B2(_08463_),
    .X(_04206_));
 sky130_fd_sc_hd__mux2_1 _18810_ (.A0(\core.csr.instruction_memoryAddress[7] ),
    .A1(_04206_),
    .S(net1649),
    .X(_04207_));
 sky130_fd_sc_hd__mux2_1 _18811_ (.A0(net479),
    .A1(_04207_),
    .S(_04169_),
    .X(_04208_));
 sky130_fd_sc_hd__mux2_1 _18812_ (.A0(_03981_),
    .A1(\core.csr.traps.mtval.csrReadData[7] ),
    .S(net759),
    .X(_04209_));
 sky130_fd_sc_hd__a21oi_1 _18813_ (.A1(net780),
    .A2(_04208_),
    .B1(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__nor2_1 _18814_ (.A(net1983),
    .B(_04210_),
    .Y(_01903_));
 sky130_fd_sc_hd__a22o_1 _18815_ (.A1(\core.csr.currentInstruction[8] ),
    .A2(net1019),
    .B1(net811),
    .B2(_08464_),
    .X(_04211_));
 sky130_fd_sc_hd__nand2_1 _18816_ (.A(net1650),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__a21oi_1 _18817_ (.A1(\core.csr.instruction_memoryAddress[8] ),
    .A2(net1645),
    .B1(net1077),
    .Y(_04213_));
 sky130_fd_sc_hd__a22o_1 _18818_ (.A1(_04058_),
    .A2(net746),
    .B1(_04212_),
    .B2(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__nand2_1 _18819_ (.A(\core.csr.traps.mtval.csrReadData[8] ),
    .B(net759),
    .Y(_04215_));
 sky130_fd_sc_hd__o211a_1 _18820_ (.A1(_03984_),
    .A2(net759),
    .B1(_04214_),
    .C1(_04215_),
    .X(_04216_));
 sky130_fd_sc_hd__nor2_1 _18821_ (.A(net1981),
    .B(_04216_),
    .Y(_01904_));
 sky130_fd_sc_hd__a22o_1 _18822_ (.A1(\core.csr.currentInstruction[9] ),
    .A2(net1019),
    .B1(net811),
    .B2(_08489_),
    .X(_04217_));
 sky130_fd_sc_hd__nand2_1 _18823_ (.A(net1650),
    .B(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__a21oi_1 _18824_ (.A1(\core.csr.instruction_memoryAddress[9] ),
    .A2(net1645),
    .B1(net1077),
    .Y(_04219_));
 sky130_fd_sc_hd__a22o_1 _18825_ (.A1(_04061_),
    .A2(net745),
    .B1(_04218_),
    .B2(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__nand2_1 _18826_ (.A(\core.csr.traps.mtval.csrReadData[9] ),
    .B(net758),
    .Y(_04221_));
 sky130_fd_sc_hd__o211a_1 _18827_ (.A1(_03986_),
    .A2(net758),
    .B1(_04220_),
    .C1(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__nor2_1 _18828_ (.A(net1978),
    .B(_04222_),
    .Y(_01905_));
 sky130_fd_sc_hd__a22o_1 _18829_ (.A1(\core.csr.currentInstruction[10] ),
    .A2(net1019),
    .B1(net811),
    .B2(_08503_),
    .X(_04223_));
 sky130_fd_sc_hd__nand2_1 _18830_ (.A(net1650),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__a21oi_1 _18831_ (.A1(\core.csr.instruction_memoryAddress[10] ),
    .A2(net1646),
    .B1(net1078),
    .Y(_04225_));
 sky130_fd_sc_hd__a22o_1 _18832_ (.A1(_04064_),
    .A2(net745),
    .B1(_04224_),
    .B2(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__nand2_1 _18833_ (.A(\core.csr.traps.mtval.csrReadData[10] ),
    .B(net758),
    .Y(_04227_));
 sky130_fd_sc_hd__o211a_1 _18834_ (.A1(_03988_),
    .A2(net758),
    .B1(_04226_),
    .C1(_04227_),
    .X(_04228_));
 sky130_fd_sc_hd__nor2_1 _18835_ (.A(net1977),
    .B(_04228_),
    .Y(_01906_));
 sky130_fd_sc_hd__a22o_1 _18836_ (.A1(\core.csr.currentInstruction[11] ),
    .A2(net1019),
    .B1(_07503_),
    .B2(_08367_),
    .X(_04229_));
 sky130_fd_sc_hd__nand2_1 _18837_ (.A(net1649),
    .B(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__a21oi_1 _18838_ (.A1(\core.csr.instruction_memoryAddress[11] ),
    .A2(net1645),
    .B1(net1078),
    .Y(_04231_));
 sky130_fd_sc_hd__a22o_1 _18839_ (.A1(_04067_),
    .A2(net745),
    .B1(_04230_),
    .B2(_04231_),
    .X(_04232_));
 sky130_fd_sc_hd__nand2_1 _18840_ (.A(\core.csr.traps.mtval.csrReadData[11] ),
    .B(net760),
    .Y(_04233_));
 sky130_fd_sc_hd__o211a_1 _18841_ (.A1(_03990_),
    .A2(net760),
    .B1(_04232_),
    .C1(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__nor2_1 _18842_ (.A(net1978),
    .B(_04234_),
    .Y(_01907_));
 sky130_fd_sc_hd__a22o_1 _18843_ (.A1(\core.csr.currentInstruction[12] ),
    .A2(net1018),
    .B1(net810),
    .B2(_08333_),
    .X(_04235_));
 sky130_fd_sc_hd__nand2_1 _18844_ (.A(net1649),
    .B(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__a21oi_1 _18845_ (.A1(\core.csr.instruction_memoryAddress[12] ),
    .A2(net1645),
    .B1(net1077),
    .Y(_04237_));
 sky130_fd_sc_hd__a22o_1 _18846_ (.A1(_04070_),
    .A2(net745),
    .B1(_04236_),
    .B2(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__nand2_1 _18847_ (.A(\core.csr.traps.mtval.csrReadData[12] ),
    .B(net758),
    .Y(_04239_));
 sky130_fd_sc_hd__o211a_1 _18848_ (.A1(_03992_),
    .A2(net758),
    .B1(_04238_),
    .C1(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__nor2_1 _18849_ (.A(net1975),
    .B(_04240_),
    .Y(_01908_));
 sky130_fd_sc_hd__a22o_1 _18850_ (.A1(net1885),
    .A2(net1018),
    .B1(net810),
    .B2(_08332_),
    .X(_04241_));
 sky130_fd_sc_hd__nand2_1 _18851_ (.A(net1649),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__a21oi_1 _18852_ (.A1(\core.csr.instruction_memoryAddress[13] ),
    .A2(net1645),
    .B1(net1077),
    .Y(_04243_));
 sky130_fd_sc_hd__a22o_1 _18853_ (.A1(_04073_),
    .A2(net745),
    .B1(_04242_),
    .B2(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__nand2_1 _18854_ (.A(\core.csr.traps.mtval.csrReadData[13] ),
    .B(net758),
    .Y(_04245_));
 sky130_fd_sc_hd__o211a_1 _18855_ (.A1(_03994_),
    .A2(net758),
    .B1(_04244_),
    .C1(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__nor2_1 _18856_ (.A(net1975),
    .B(_04246_),
    .Y(_01909_));
 sky130_fd_sc_hd__a22o_1 _18857_ (.A1(\core.csr.currentInstruction[14] ),
    .A2(net1018),
    .B1(net810),
    .B2(_08331_),
    .X(_04247_));
 sky130_fd_sc_hd__nand2_1 _18858_ (.A(net1649),
    .B(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__a21oi_1 _18859_ (.A1(\core.csr.instruction_memoryAddress[14] ),
    .A2(net1645),
    .B1(net1077),
    .Y(_04249_));
 sky130_fd_sc_hd__a22o_1 _18860_ (.A1(_04076_),
    .A2(net745),
    .B1(_04248_),
    .B2(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__nand2_1 _18861_ (.A(\core.csr.traps.mtval.csrReadData[14] ),
    .B(net758),
    .Y(_04251_));
 sky130_fd_sc_hd__o211a_1 _18862_ (.A1(_03996_),
    .A2(net758),
    .B1(_04250_),
    .C1(_04251_),
    .X(_04252_));
 sky130_fd_sc_hd__nor2_1 _18863_ (.A(net1976),
    .B(_04252_),
    .Y(_01910_));
 sky130_fd_sc_hd__a22o_1 _18864_ (.A1(\core.csr.currentInstruction[15] ),
    .A2(net1018),
    .B1(net810),
    .B2(_08330_),
    .X(_04253_));
 sky130_fd_sc_hd__nand2_1 _18865_ (.A(net1649),
    .B(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__a21oi_1 _18866_ (.A1(\core.csr.instruction_memoryAddress[15] ),
    .A2(net1645),
    .B1(net1077),
    .Y(_04255_));
 sky130_fd_sc_hd__a22o_1 _18867_ (.A1(_04079_),
    .A2(net745),
    .B1(_04254_),
    .B2(_04255_),
    .X(_04256_));
 sky130_fd_sc_hd__nand2_1 _18868_ (.A(\core.csr.traps.mtval.csrReadData[15] ),
    .B(net757),
    .Y(_04257_));
 sky130_fd_sc_hd__o211a_1 _18869_ (.A1(_03998_),
    .A2(net757),
    .B1(_04256_),
    .C1(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__nor2_1 _18870_ (.A(net1974),
    .B(_04258_),
    .Y(_01911_));
 sky130_fd_sc_hd__a22o_1 _18871_ (.A1(\core.csr.currentInstruction[16] ),
    .A2(net1017),
    .B1(net809),
    .B2(_08329_),
    .X(_04259_));
 sky130_fd_sc_hd__nand2_1 _18872_ (.A(net1649),
    .B(_04259_),
    .Y(_04260_));
 sky130_fd_sc_hd__a21oi_1 _18873_ (.A1(\core.csr.instruction_memoryAddress[16] ),
    .A2(net1645),
    .B1(net1077),
    .Y(_04261_));
 sky130_fd_sc_hd__a22o_1 _18874_ (.A1(_04082_),
    .A2(net744),
    .B1(_04260_),
    .B2(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__nand2_1 _18875_ (.A(\core.csr.traps.mtval.csrReadData[16] ),
    .B(net757),
    .Y(_04263_));
 sky130_fd_sc_hd__o211a_1 _18876_ (.A1(_04000_),
    .A2(net757),
    .B1(_04262_),
    .C1(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__nor2_1 _18877_ (.A(net1974),
    .B(_04264_),
    .Y(_01912_));
 sky130_fd_sc_hd__a22o_1 _18878_ (.A1(\core.csr.currentInstruction[17] ),
    .A2(net1016),
    .B1(net808),
    .B2(_08328_),
    .X(_04265_));
 sky130_fd_sc_hd__nand2_1 _18879_ (.A(net1647),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__a21oi_1 _18880_ (.A1(\core.csr.instruction_memoryAddress[17] ),
    .A2(net1646),
    .B1(net1077),
    .Y(_04267_));
 sky130_fd_sc_hd__a22o_1 _18881_ (.A1(_04085_),
    .A2(net743),
    .B1(_04266_),
    .B2(_04267_),
    .X(_04268_));
 sky130_fd_sc_hd__nand2_1 _18882_ (.A(\core.csr.traps.mtval.csrReadData[17] ),
    .B(net756),
    .Y(_04269_));
 sky130_fd_sc_hd__o211a_1 _18883_ (.A1(_04002_),
    .A2(net756),
    .B1(_04268_),
    .C1(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__nor2_1 _18884_ (.A(net1971),
    .B(_04270_),
    .Y(_01913_));
 sky130_fd_sc_hd__a22o_1 _18885_ (.A1(\core.csr.currentInstruction[18] ),
    .A2(net1016),
    .B1(net808),
    .B2(_08327_),
    .X(_04271_));
 sky130_fd_sc_hd__nand2_1 _18886_ (.A(net1647),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__a21oi_1 _18887_ (.A1(\core.csr.instruction_memoryAddress[18] ),
    .A2(net1644),
    .B1(net1076),
    .Y(_04273_));
 sky130_fd_sc_hd__a22o_1 _18888_ (.A1(_04088_),
    .A2(net744),
    .B1(_04272_),
    .B2(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__nand2_1 _18889_ (.A(\core.csr.traps.mtval.csrReadData[18] ),
    .B(net756),
    .Y(_04275_));
 sky130_fd_sc_hd__o211a_1 _18890_ (.A1(_04004_),
    .A2(net756),
    .B1(_04274_),
    .C1(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__nor2_1 _18891_ (.A(net1971),
    .B(_04276_),
    .Y(_01914_));
 sky130_fd_sc_hd__a22o_1 _18892_ (.A1(\core.csr.currentInstruction[19] ),
    .A2(net1016),
    .B1(net808),
    .B2(_08326_),
    .X(_04277_));
 sky130_fd_sc_hd__nand2_1 _18893_ (.A(net1648),
    .B(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__a21oi_1 _18894_ (.A1(\core.csr.instruction_memoryAddress[19] ),
    .A2(net1644),
    .B1(net1076),
    .Y(_04279_));
 sky130_fd_sc_hd__a22o_1 _18895_ (.A1(_04091_),
    .A2(net744),
    .B1(_04278_),
    .B2(_04279_),
    .X(_04280_));
 sky130_fd_sc_hd__nand2_1 _18896_ (.A(\core.csr.traps.mtval.csrReadData[19] ),
    .B(net756),
    .Y(_04281_));
 sky130_fd_sc_hd__o211a_1 _18897_ (.A1(_04006_),
    .A2(net756),
    .B1(_04280_),
    .C1(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__nor2_1 _18898_ (.A(net1966),
    .B(_04282_),
    .Y(_01915_));
 sky130_fd_sc_hd__a22o_1 _18899_ (.A1(\core.csr.currentInstruction[20] ),
    .A2(net1016),
    .B1(net809),
    .B2(_08325_),
    .X(_04283_));
 sky130_fd_sc_hd__mux2_1 _18900_ (.A0(\core.csr.instruction_memoryAddress[20] ),
    .A1(_04283_),
    .S(net1647),
    .X(_04284_));
 sky130_fd_sc_hd__mux2_1 _18901_ (.A0(net462),
    .A1(_04284_),
    .S(net1163),
    .X(_04285_));
 sky130_fd_sc_hd__nand2_1 _18902_ (.A(net776),
    .B(_04285_),
    .Y(_04286_));
 sky130_fd_sc_hd__nand2_1 _18903_ (.A(\core.csr.traps.mtval.csrReadData[20] ),
    .B(net755),
    .Y(_04287_));
 sky130_fd_sc_hd__o211a_1 _18904_ (.A1(_04008_),
    .A2(net755),
    .B1(_04286_),
    .C1(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__nor2_1 _18905_ (.A(net1968),
    .B(_04288_),
    .Y(_01916_));
 sky130_fd_sc_hd__a22o_1 _18906_ (.A1(\core.csr.currentInstruction[21] ),
    .A2(net1016),
    .B1(net809),
    .B2(_08323_),
    .X(_04289_));
 sky130_fd_sc_hd__nand2_2 _18907_ (.A(net1647),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__a21oi_1 _18908_ (.A1(\core.csr.instruction_memoryAddress[21] ),
    .A2(net1644),
    .B1(net1076),
    .Y(_04291_));
 sky130_fd_sc_hd__a22o_1 _18909_ (.A1(_04096_),
    .A2(net743),
    .B1(_04290_),
    .B2(_04291_),
    .X(_04292_));
 sky130_fd_sc_hd__nand2_1 _18910_ (.A(\core.csr.traps.mtval.csrReadData[21] ),
    .B(net754),
    .Y(_04293_));
 sky130_fd_sc_hd__o211a_1 _18911_ (.A1(_04010_),
    .A2(net754),
    .B1(_04292_),
    .C1(_04293_),
    .X(_04294_));
 sky130_fd_sc_hd__nor2_1 _18912_ (.A(net1963),
    .B(_04294_),
    .Y(_01917_));
 sky130_fd_sc_hd__o2bb2a_2 _18913_ (.A1_N(\core.csr.currentInstruction[22] ),
    .A2_N(net1017),
    .B1(_07504_),
    .B2(_08322_),
    .X(_04295_));
 sky130_fd_sc_hd__mux2_1 _18914_ (.A0(_04405_),
    .A1(_04295_),
    .S(net1648),
    .X(_04296_));
 sky130_fd_sc_hd__a22o_1 _18915_ (.A1(_04099_),
    .A2(net743),
    .B1(_04296_),
    .B2(net1163),
    .X(_04297_));
 sky130_fd_sc_hd__nand2_1 _18916_ (.A(\core.csr.traps.mtval.csrReadData[22] ),
    .B(net754),
    .Y(_04298_));
 sky130_fd_sc_hd__o211a_1 _18917_ (.A1(_04012_),
    .A2(net754),
    .B1(_04297_),
    .C1(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__nor2_1 _18918_ (.A(net1963),
    .B(_04299_),
    .Y(_01918_));
 sky130_fd_sc_hd__a22o_1 _18919_ (.A1(\core.csr.currentInstruction[23] ),
    .A2(net1016),
    .B1(net808),
    .B2(_08321_),
    .X(_04300_));
 sky130_fd_sc_hd__nand2_2 _18920_ (.A(net1647),
    .B(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__a21oi_1 _18921_ (.A1(\core.csr.instruction_memoryAddress[23] ),
    .A2(net1644),
    .B1(net1076),
    .Y(_04302_));
 sky130_fd_sc_hd__a22o_1 _18922_ (.A1(_04102_),
    .A2(net743),
    .B1(_04301_),
    .B2(_04302_),
    .X(_04303_));
 sky130_fd_sc_hd__nand2_1 _18923_ (.A(\core.csr.traps.mtval.csrReadData[23] ),
    .B(net754),
    .Y(_04304_));
 sky130_fd_sc_hd__o211a_1 _18924_ (.A1(_04014_),
    .A2(net754),
    .B1(_04303_),
    .C1(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__nor2_1 _18925_ (.A(net1962),
    .B(_04305_),
    .Y(_01919_));
 sky130_fd_sc_hd__a22o_1 _18926_ (.A1(\core.csr.currentInstruction[24] ),
    .A2(net1016),
    .B1(net808),
    .B2(_08342_),
    .X(_04306_));
 sky130_fd_sc_hd__nand2_2 _18927_ (.A(net1647),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21oi_1 _18928_ (.A1(\core.csr.instruction_memoryAddress[24] ),
    .A2(net1644),
    .B1(net1076),
    .Y(_04308_));
 sky130_fd_sc_hd__a22o_1 _18929_ (.A1(_04105_),
    .A2(net743),
    .B1(_04307_),
    .B2(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__nand2_1 _18930_ (.A(\core.csr.traps.mtval.csrReadData[24] ),
    .B(net754),
    .Y(_04310_));
 sky130_fd_sc_hd__o211a_1 _18931_ (.A1(_04016_),
    .A2(net754),
    .B1(_04309_),
    .C1(_04310_),
    .X(_04311_));
 sky130_fd_sc_hd__nor2_1 _18932_ (.A(net1962),
    .B(_04311_),
    .Y(_01920_));
 sky130_fd_sc_hd__a22o_1 _18933_ (.A1(\core.csr.currentInstruction[25] ),
    .A2(net1016),
    .B1(net808),
    .B2(_08341_),
    .X(_04312_));
 sky130_fd_sc_hd__nand2_1 _18934_ (.A(net1648),
    .B(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__a21oi_1 _18935_ (.A1(\core.csr.instruction_memoryAddress[25] ),
    .A2(net1644),
    .B1(net1076),
    .Y(_04314_));
 sky130_fd_sc_hd__a22o_1 _18936_ (.A1(_04108_),
    .A2(net743),
    .B1(_04313_),
    .B2(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__nand2_1 _18937_ (.A(\core.csr.traps.mtval.csrReadData[25] ),
    .B(net757),
    .Y(_04316_));
 sky130_fd_sc_hd__o211a_1 _18938_ (.A1(_04018_),
    .A2(net755),
    .B1(_04315_),
    .C1(_04316_),
    .X(_04317_));
 sky130_fd_sc_hd__nor2_1 _18939_ (.A(net1965),
    .B(_04317_),
    .Y(_01921_));
 sky130_fd_sc_hd__a22o_1 _18940_ (.A1(\core.csr.currentInstruction[26] ),
    .A2(net1016),
    .B1(net808),
    .B2(_08340_),
    .X(_04318_));
 sky130_fd_sc_hd__nand2_1 _18941_ (.A(net1647),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__a21oi_1 _18942_ (.A1(\core.csr.instruction_memoryAddress[26] ),
    .A2(net1644),
    .B1(net1078),
    .Y(_04320_));
 sky130_fd_sc_hd__a22o_1 _18943_ (.A1(_04111_),
    .A2(net743),
    .B1(_04319_),
    .B2(_04320_),
    .X(_04321_));
 sky130_fd_sc_hd__nand2_1 _18944_ (.A(\core.csr.traps.mtval.csrReadData[26] ),
    .B(net755),
    .Y(_04322_));
 sky130_fd_sc_hd__o211a_1 _18945_ (.A1(_04020_),
    .A2(net755),
    .B1(_04321_),
    .C1(_04322_),
    .X(_04323_));
 sky130_fd_sc_hd__nor2_1 _18946_ (.A(net1965),
    .B(_04323_),
    .Y(_01922_));
 sky130_fd_sc_hd__a22o_1 _18947_ (.A1(\core.csr.currentInstruction[27] ),
    .A2(net1017),
    .B1(net808),
    .B2(_08339_),
    .X(_04324_));
 sky130_fd_sc_hd__nand2_1 _18948_ (.A(net1647),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__a21oi_1 _18949_ (.A1(\core.csr.instruction_memoryAddress[27] ),
    .A2(net1646),
    .B1(net1078),
    .Y(_04326_));
 sky130_fd_sc_hd__a22o_1 _18950_ (.A1(_04114_),
    .A2(net744),
    .B1(_04325_),
    .B2(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__nand2_1 _18951_ (.A(\core.csr.traps.mtval.csrReadData[27] ),
    .B(net756),
    .Y(_04328_));
 sky130_fd_sc_hd__o211a_1 _18952_ (.A1(_04022_),
    .A2(net756),
    .B1(_04327_),
    .C1(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__nor2_1 _18953_ (.A(net1966),
    .B(_04329_),
    .Y(_01923_));
 sky130_fd_sc_hd__a22o_2 _18954_ (.A1(\core.csr.currentInstruction[28] ),
    .A2(net1016),
    .B1(net808),
    .B2(_08094_),
    .X(_04330_));
 sky130_fd_sc_hd__nand2_1 _18955_ (.A(net1648),
    .B(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__a21oi_1 _18956_ (.A1(\core.csr.instruction_memoryAddress[28] ),
    .A2(net1644),
    .B1(net1076),
    .Y(_04332_));
 sky130_fd_sc_hd__a22o_1 _18957_ (.A1(_04117_),
    .A2(net743),
    .B1(_04331_),
    .B2(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__nand2_1 _18958_ (.A(\core.csr.traps.mtval.csrReadData[28] ),
    .B(net755),
    .Y(_04334_));
 sky130_fd_sc_hd__o211a_1 _18959_ (.A1(_04024_),
    .A2(net755),
    .B1(_04333_),
    .C1(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__nor2_1 _18960_ (.A(net1964),
    .B(_04335_),
    .Y(_01924_));
 sky130_fd_sc_hd__o2bb2a_1 _18961_ (.A1_N(\core.csr.currentInstruction[29] ),
    .A2_N(net1017),
    .B1(_07504_),
    .B2(_08093_),
    .X(_04336_));
 sky130_fd_sc_hd__mux2_2 _18962_ (.A0(_04404_),
    .A1(_04336_),
    .S(net1647),
    .X(_04337_));
 sky130_fd_sc_hd__a22o_1 _18963_ (.A1(_04120_),
    .A2(net743),
    .B1(_04337_),
    .B2(net1163),
    .X(_04338_));
 sky130_fd_sc_hd__nand2_1 _18964_ (.A(\core.csr.traps.mtval.csrReadData[29] ),
    .B(net755),
    .Y(_04339_));
 sky130_fd_sc_hd__o211a_1 _18965_ (.A1(_04026_),
    .A2(net755),
    .B1(_04338_),
    .C1(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__nor2_1 _18966_ (.A(net1965),
    .B(_04340_),
    .Y(_01925_));
 sky130_fd_sc_hd__a22o_1 _18967_ (.A1(\core.csr.currentInstruction[30] ),
    .A2(net1017),
    .B1(net808),
    .B2(_08089_),
    .X(_04341_));
 sky130_fd_sc_hd__nand2_4 _18968_ (.A(net1649),
    .B(_04341_),
    .Y(_04342_));
 sky130_fd_sc_hd__a21oi_1 _18969_ (.A1(\core.csr.instruction_memoryAddress[30] ),
    .A2(net1644),
    .B1(net1076),
    .Y(_04343_));
 sky130_fd_sc_hd__a22o_1 _18970_ (.A1(_04123_),
    .A2(net743),
    .B1(_04342_),
    .B2(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__nand2_1 _18971_ (.A(\core.csr.traps.mtval.csrReadData[30] ),
    .B(net754),
    .Y(_04345_));
 sky130_fd_sc_hd__o211a_1 _18972_ (.A1(_04028_),
    .A2(net754),
    .B1(_04344_),
    .C1(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__nor2_1 _18973_ (.A(net1963),
    .B(_04346_),
    .Y(_01926_));
 sky130_fd_sc_hd__a22o_1 _18974_ (.A1(\core.csr.currentInstruction[31] ),
    .A2(net1017),
    .B1(net809),
    .B2(_08091_),
    .X(_04347_));
 sky130_fd_sc_hd__nand2_1 _18975_ (.A(net1647),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__a21oi_2 _18976_ (.A1(\core.csr.instruction_memoryAddress[31] ),
    .A2(net1644),
    .B1(net1076),
    .Y(_04349_));
 sky130_fd_sc_hd__a22o_1 _18977_ (.A1(_04126_),
    .A2(net744),
    .B1(_04348_),
    .B2(_04349_),
    .X(_04350_));
 sky130_fd_sc_hd__nand2_1 _18978_ (.A(\core.csr.traps.mtval.csrReadData[31] ),
    .B(net756),
    .Y(_04351_));
 sky130_fd_sc_hd__o211a_1 _18979_ (.A1(_04031_),
    .A2(net756),
    .B1(_04350_),
    .C1(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__nor2_1 _18980_ (.A(net1966),
    .B(_04352_),
    .Y(_01927_));
 sky130_fd_sc_hd__or3_4 _18981_ (.A(_03737_),
    .B(_03885_),
    .C(_03886_),
    .X(_04353_));
 sky130_fd_sc_hd__and2_2 _18982_ (.A(net749),
    .B(net832),
    .X(_04354_));
 sky130_fd_sc_hd__nand2_1 _18983_ (.A(net749),
    .B(net833),
    .Y(_04355_));
 sky130_fd_sc_hd__or2_1 _18984_ (.A(\core.csr.traps.mip.csrReadData[0] ),
    .B(net735),
    .X(_04356_));
 sky130_fd_sc_hd__and2_2 _18985_ (.A(net1932),
    .B(net749),
    .X(_04357_));
 sky130_fd_sc_hd__o211a_1 _18986_ (.A1(_03758_),
    .A2(net832),
    .B1(_04356_),
    .C1(net730),
    .X(_01928_));
 sky130_fd_sc_hd__or2_1 _18987_ (.A(\core.csr.traps.mip.csrReadData[1] ),
    .B(net735),
    .X(_04358_));
 sky130_fd_sc_hd__o211a_1 _18988_ (.A1(_03762_),
    .A2(net833),
    .B1(net730),
    .C1(_04358_),
    .X(_01929_));
 sky130_fd_sc_hd__or2_1 _18989_ (.A(\core.csr.traps.mip.csrReadData[2] ),
    .B(net734),
    .X(_04359_));
 sky130_fd_sc_hd__o211a_1 _18990_ (.A1(_03766_),
    .A2(net833),
    .B1(net731),
    .C1(_04359_),
    .X(_01930_));
 sky130_fd_sc_hd__or2_1 _18991_ (.A(\core.csr.traps.mip.csrReadData[3] ),
    .B(net734),
    .X(_04360_));
 sky130_fd_sc_hd__o211a_1 _18992_ (.A1(_03770_),
    .A2(net833),
    .B1(net731),
    .C1(_04360_),
    .X(_01931_));
 sky130_fd_sc_hd__or2_1 _18993_ (.A(\core.csr.traps.mip.csrReadData[4] ),
    .B(net734),
    .X(_04361_));
 sky130_fd_sc_hd__o211a_1 _18994_ (.A1(_03774_),
    .A2(net833),
    .B1(net731),
    .C1(_04361_),
    .X(_01932_));
 sky130_fd_sc_hd__or2_1 _18995_ (.A(\core.csr.traps.mip.csrReadData[5] ),
    .B(net735),
    .X(_04362_));
 sky130_fd_sc_hd__o211a_1 _18996_ (.A1(_03778_),
    .A2(net833),
    .B1(net731),
    .C1(_04362_),
    .X(_01933_));
 sky130_fd_sc_hd__or2_1 _18997_ (.A(\core.csr.traps.mip.csrReadData[6] ),
    .B(net735),
    .X(_04363_));
 sky130_fd_sc_hd__o211a_1 _18998_ (.A1(_03782_),
    .A2(net833),
    .B1(net731),
    .C1(_04363_),
    .X(_01934_));
 sky130_fd_sc_hd__or2_1 _18999_ (.A(\core.csr.traps.mip.csrReadData[7] ),
    .B(net734),
    .X(_04364_));
 sky130_fd_sc_hd__o211a_1 _19000_ (.A1(_03786_),
    .A2(net832),
    .B1(net730),
    .C1(_04364_),
    .X(_01935_));
 sky130_fd_sc_hd__or2_1 _19001_ (.A(\core.csr.traps.mip.csrReadData[8] ),
    .B(net734),
    .X(_04365_));
 sky130_fd_sc_hd__o211a_1 _19002_ (.A1(_03790_),
    .A2(net833),
    .B1(net731),
    .C1(_04365_),
    .X(_01936_));
 sky130_fd_sc_hd__or2_1 _19003_ (.A(\core.csr.traps.mip.csrReadData[9] ),
    .B(net734),
    .X(_04366_));
 sky130_fd_sc_hd__o211a_1 _19004_ (.A1(_03794_),
    .A2(net832),
    .B1(net730),
    .C1(_04366_),
    .X(_01937_));
 sky130_fd_sc_hd__or2_1 _19005_ (.A(\core.csr.traps.mip.csrReadData[10] ),
    .B(net734),
    .X(_04367_));
 sky130_fd_sc_hd__o211a_1 _19006_ (.A1(_03798_),
    .A2(net832),
    .B1(net730),
    .C1(_04367_),
    .X(_01938_));
 sky130_fd_sc_hd__or2_1 _19007_ (.A(\core.csr.traps.mip.csrReadData[11] ),
    .B(net734),
    .X(_04368_));
 sky130_fd_sc_hd__o211a_1 _19008_ (.A1(_03802_),
    .A2(net832),
    .B1(net730),
    .C1(_04368_),
    .X(_01939_));
 sky130_fd_sc_hd__or2_1 _19009_ (.A(\core.csr.traps.mip.csrReadData[12] ),
    .B(net734),
    .X(_04369_));
 sky130_fd_sc_hd__o211a_1 _19010_ (.A1(_03806_),
    .A2(net832),
    .B1(net730),
    .C1(_04369_),
    .X(_01940_));
 sky130_fd_sc_hd__or2_1 _19011_ (.A(\core.csr.traps.mip.csrReadData[13] ),
    .B(net733),
    .X(_04370_));
 sky130_fd_sc_hd__o211a_1 _19012_ (.A1(_03810_),
    .A2(net832),
    .B1(net730),
    .C1(_04370_),
    .X(_01941_));
 sky130_fd_sc_hd__or2_1 _19013_ (.A(\core.csr.traps.mip.csrReadData[14] ),
    .B(net734),
    .X(_04371_));
 sky130_fd_sc_hd__o211a_1 _19014_ (.A1(_03814_),
    .A2(net832),
    .B1(net730),
    .C1(_04371_),
    .X(_01942_));
 sky130_fd_sc_hd__or2_1 _19015_ (.A(\core.csr.traps.mip.csrReadData[15] ),
    .B(net733),
    .X(_04372_));
 sky130_fd_sc_hd__o211a_1 _19016_ (.A1(_03818_),
    .A2(net832),
    .B1(net730),
    .C1(_04372_),
    .X(_01943_));
 sky130_fd_sc_hd__o21a_4 _19017_ (.A1(_07463_),
    .A2(_07467_),
    .B1(_04165_),
    .X(_04373_));
 sky130_fd_sc_hd__a221o_1 _19018_ (.A1(_03822_),
    .A2(net748),
    .B1(_04373_),
    .B2(_07456_),
    .C1(net737),
    .X(_04374_));
 sky130_fd_sc_hd__o211a_1 _19019_ (.A1(\core.csr.traps.mip.csrReadData[16] ),
    .A2(net733),
    .B1(_04374_),
    .C1(net1912),
    .X(_01944_));
 sky130_fd_sc_hd__a221o_1 _19020_ (.A1(_03826_),
    .A2(net748),
    .B1(_04373_),
    .B2(_07453_),
    .C1(net737),
    .X(_04375_));
 sky130_fd_sc_hd__o211a_1 _19021_ (.A1(\core.csr.traps.mip.csrReadData[17] ),
    .A2(net733),
    .B1(_04375_),
    .C1(net1911),
    .X(_01945_));
 sky130_fd_sc_hd__a221o_1 _19022_ (.A1(_03830_),
    .A2(net748),
    .B1(net742),
    .B2(_07461_),
    .C1(net736),
    .X(_04376_));
 sky130_fd_sc_hd__o211a_1 _19023_ (.A1(\core.csr.traps.mip.csrReadData[18] ),
    .A2(net733),
    .B1(_04376_),
    .C1(net1911),
    .X(_01946_));
 sky130_fd_sc_hd__a221o_1 _19024_ (.A1(_03834_),
    .A2(net748),
    .B1(_04165_),
    .B2(_07462_),
    .C1(net737),
    .X(_04377_));
 sky130_fd_sc_hd__o211a_1 _19025_ (.A1(\core.csr.traps.mip.csrReadData[19] ),
    .A2(net733),
    .B1(_04377_),
    .C1(net1903),
    .X(_01947_));
 sky130_fd_sc_hd__a221o_1 _19026_ (.A1(_03838_),
    .A2(net747),
    .B1(net742),
    .B2(_07447_),
    .C1(net736),
    .X(_04378_));
 sky130_fd_sc_hd__o211a_1 _19027_ (.A1(\core.csr.traps.mip.csrReadData[20] ),
    .A2(net733),
    .B1(_04378_),
    .C1(net1897),
    .X(_01948_));
 sky130_fd_sc_hd__a221o_1 _19028_ (.A1(_03842_),
    .A2(net747),
    .B1(net742),
    .B2(_07449_),
    .C1(net736),
    .X(_04379_));
 sky130_fd_sc_hd__o211a_1 _19029_ (.A1(\core.csr.traps.mip.csrReadData[21] ),
    .A2(net732),
    .B1(_04379_),
    .C1(net1895),
    .X(_01949_));
 sky130_fd_sc_hd__a221o_1 _19030_ (.A1(_03846_),
    .A2(net747),
    .B1(net742),
    .B2(_07458_),
    .C1(net736),
    .X(_04380_));
 sky130_fd_sc_hd__o211a_1 _19031_ (.A1(\core.csr.traps.mip.csrReadData[22] ),
    .A2(net732),
    .B1(_04380_),
    .C1(net1896),
    .X(_01950_));
 sky130_fd_sc_hd__a221o_1 _19032_ (.A1(_03850_),
    .A2(net747),
    .B1(_04165_),
    .B2(_07448_),
    .C1(net736),
    .X(_04381_));
 sky130_fd_sc_hd__o211a_1 _19033_ (.A1(\core.csr.traps.mip.csrReadData[23] ),
    .A2(net732),
    .B1(_04381_),
    .C1(net1895),
    .X(_01951_));
 sky130_fd_sc_hd__a221o_1 _19034_ (.A1(_03854_),
    .A2(net747),
    .B1(net742),
    .B2(_07450_),
    .C1(net736),
    .X(_04382_));
 sky130_fd_sc_hd__o211a_1 _19035_ (.A1(\core.csr.traps.mip.csrReadData[24] ),
    .A2(net732),
    .B1(_04382_),
    .C1(net1896),
    .X(_01952_));
 sky130_fd_sc_hd__a221o_1 _19036_ (.A1(_03858_),
    .A2(net747),
    .B1(net742),
    .B2(_07457_),
    .C1(net736),
    .X(_04383_));
 sky130_fd_sc_hd__o211a_1 _19037_ (.A1(\core.csr.traps.mip.csrReadData[25] ),
    .A2(net732),
    .B1(_04383_),
    .C1(net1897),
    .X(_01953_));
 sky130_fd_sc_hd__a221o_1 _19038_ (.A1(_03862_),
    .A2(net747),
    .B1(net742),
    .B2(_07459_),
    .C1(net736),
    .X(_04384_));
 sky130_fd_sc_hd__o211a_1 _19039_ (.A1(\core.csr.traps.mip.csrReadData[26] ),
    .A2(net732),
    .B1(_04384_),
    .C1(net1901),
    .X(_01954_));
 sky130_fd_sc_hd__a221o_1 _19040_ (.A1(_03866_),
    .A2(net748),
    .B1(_04373_),
    .B2(_07452_),
    .C1(net737),
    .X(_04385_));
 sky130_fd_sc_hd__o211a_1 _19041_ (.A1(\core.csr.traps.mip.csrReadData[27] ),
    .A2(net732),
    .B1(_04385_),
    .C1(net1903),
    .X(_01955_));
 sky130_fd_sc_hd__a221o_1 _19042_ (.A1(_03870_),
    .A2(net747),
    .B1(net742),
    .B2(_07455_),
    .C1(net736),
    .X(_04386_));
 sky130_fd_sc_hd__o211a_1 _19043_ (.A1(\core.csr.traps.mip.csrReadData[28] ),
    .A2(net732),
    .B1(_04386_),
    .C1(net1898),
    .X(_01956_));
 sky130_fd_sc_hd__a221o_1 _19044_ (.A1(_03874_),
    .A2(net747),
    .B1(_04373_),
    .B2(_07454_),
    .C1(net737),
    .X(_04387_));
 sky130_fd_sc_hd__o211a_1 _19045_ (.A1(\core.csr.traps.mip.csrReadData[29] ),
    .A2(net733),
    .B1(_04387_),
    .C1(net1902),
    .X(_01957_));
 sky130_fd_sc_hd__a221o_1 _19046_ (.A1(_03878_),
    .A2(net747),
    .B1(net742),
    .B2(_07451_),
    .C1(net736),
    .X(_04388_));
 sky130_fd_sc_hd__o211a_1 _19047_ (.A1(\core.csr.traps.mip.csrReadData[30] ),
    .A2(net732),
    .B1(_04388_),
    .C1(net1895),
    .X(_01958_));
 sky130_fd_sc_hd__a221o_1 _19048_ (.A1(_03882_),
    .A2(net748),
    .B1(net742),
    .B2(_07460_),
    .C1(net737),
    .X(_04389_));
 sky130_fd_sc_hd__o211a_1 _19049_ (.A1(\core.csr.traps.mip.csrReadData[31] ),
    .A2(net732),
    .B1(_04389_),
    .C1(net1903),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_1 _19050_ (.A0(\core.pipe2_stall ),
    .A1(net1884),
    .S(net686),
    .X(_04390_));
 sky130_fd_sc_hd__or2_1 _19051_ (.A(net1994),
    .B(_04390_),
    .X(_01960_));
 sky130_fd_sc_hd__clkbuf_2 _19052_ (.A(\core.registers[0][0] ),
    .X(_01313_));
 sky130_fd_sc_hd__clkbuf_2 _19053_ (.A(\core.registers[0][1] ),
    .X(_01314_));
 sky130_fd_sc_hd__clkbuf_2 _19054_ (.A(\core.registers[0][2] ),
    .X(_01315_));
 sky130_fd_sc_hd__clkbuf_2 _19055_ (.A(\core.registers[0][3] ),
    .X(_01316_));
 sky130_fd_sc_hd__clkbuf_2 _19056_ (.A(\core.registers[0][4] ),
    .X(_01317_));
 sky130_fd_sc_hd__clkbuf_2 _19057_ (.A(\core.registers[0][5] ),
    .X(_01318_));
 sky130_fd_sc_hd__clkbuf_2 _19058_ (.A(\core.registers[0][6] ),
    .X(_01319_));
 sky130_fd_sc_hd__clkbuf_2 _19059_ (.A(\core.registers[0][7] ),
    .X(_01320_));
 sky130_fd_sc_hd__clkbuf_2 _19060_ (.A(\core.registers[0][8] ),
    .X(_01321_));
 sky130_fd_sc_hd__clkbuf_2 _19061_ (.A(\core.registers[0][9] ),
    .X(_01322_));
 sky130_fd_sc_hd__clkbuf_2 _19062_ (.A(\core.registers[0][10] ),
    .X(_01323_));
 sky130_fd_sc_hd__clkbuf_2 _19063_ (.A(\core.registers[0][11] ),
    .X(_01324_));
 sky130_fd_sc_hd__clkbuf_2 _19064_ (.A(\core.registers[0][12] ),
    .X(_01325_));
 sky130_fd_sc_hd__clkbuf_2 _19065_ (.A(\core.registers[0][13] ),
    .X(_01326_));
 sky130_fd_sc_hd__clkbuf_2 _19066_ (.A(\core.registers[0][14] ),
    .X(_01327_));
 sky130_fd_sc_hd__clkbuf_2 _19067_ (.A(\core.registers[0][15] ),
    .X(_01328_));
 sky130_fd_sc_hd__clkbuf_2 _19068_ (.A(\core.registers[0][16] ),
    .X(_01329_));
 sky130_fd_sc_hd__clkbuf_2 _19069_ (.A(\core.registers[0][17] ),
    .X(_01330_));
 sky130_fd_sc_hd__clkbuf_2 _19070_ (.A(\core.registers[0][18] ),
    .X(_01331_));
 sky130_fd_sc_hd__clkbuf_2 _19071_ (.A(\core.registers[0][19] ),
    .X(_01332_));
 sky130_fd_sc_hd__clkbuf_2 _19072_ (.A(\core.registers[0][20] ),
    .X(_01333_));
 sky130_fd_sc_hd__clkbuf_2 _19073_ (.A(\core.registers[0][21] ),
    .X(_01334_));
 sky130_fd_sc_hd__clkbuf_2 _19074_ (.A(\core.registers[0][22] ),
    .X(_01335_));
 sky130_fd_sc_hd__clkbuf_2 _19075_ (.A(\core.registers[0][23] ),
    .X(_01336_));
 sky130_fd_sc_hd__clkbuf_2 _19076_ (.A(\core.registers[0][24] ),
    .X(_01337_));
 sky130_fd_sc_hd__clkbuf_2 _19077_ (.A(\core.registers[0][25] ),
    .X(_01338_));
 sky130_fd_sc_hd__clkbuf_2 _19078_ (.A(\core.registers[0][26] ),
    .X(_01339_));
 sky130_fd_sc_hd__clkbuf_2 _19079_ (.A(\core.registers[0][27] ),
    .X(_01340_));
 sky130_fd_sc_hd__clkbuf_2 _19080_ (.A(\core.registers[0][28] ),
    .X(_01341_));
 sky130_fd_sc_hd__clkbuf_2 _19081_ (.A(\core.registers[0][29] ),
    .X(_01342_));
 sky130_fd_sc_hd__clkbuf_2 _19082_ (.A(\core.registers[0][30] ),
    .X(_01343_));
 sky130_fd_sc_hd__clkbuf_2 _19083_ (.A(\core.registers[0][31] ),
    .X(_01344_));
 sky130_fd_sc_hd__dfxtp_2 _19084_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00000_),
    .Q(\core.csr.currentInstruction[0] ));
 sky130_fd_sc_hd__dfxtp_2 _19085_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00001_),
    .Q(\core.csr.currentInstruction[1] ));
 sky130_fd_sc_hd__dfxtp_4 _19086_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00002_),
    .Q(\core.csr.currentInstruction[2] ));
 sky130_fd_sc_hd__dfxtp_4 _19087_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00003_),
    .Q(\core.csr.currentInstruction[3] ));
 sky130_fd_sc_hd__dfxtp_4 _19088_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00004_),
    .Q(\core.csr.currentInstruction[4] ));
 sky130_fd_sc_hd__dfxtp_4 _19089_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00005_),
    .Q(\core.csr.currentInstruction[5] ));
 sky130_fd_sc_hd__dfxtp_4 _19090_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00006_),
    .Q(\core.csr.currentInstruction[6] ));
 sky130_fd_sc_hd__dfxtp_4 _19091_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00007_),
    .Q(\core.csr.currentInstruction[7] ));
 sky130_fd_sc_hd__dfxtp_4 _19092_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00008_),
    .Q(\core.csr.currentInstruction[8] ));
 sky130_fd_sc_hd__dfxtp_4 _19093_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00009_),
    .Q(\core.csr.currentInstruction[9] ));
 sky130_fd_sc_hd__dfxtp_4 _19094_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00010_),
    .Q(\core.csr.currentInstruction[10] ));
 sky130_fd_sc_hd__dfxtp_4 _19095_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00011_),
    .Q(\core.csr.currentInstruction[11] ));
 sky130_fd_sc_hd__dfxtp_4 _19096_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00012_),
    .Q(\core.csr.currentInstruction[12] ));
 sky130_fd_sc_hd__dfxtp_2 _19097_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00013_),
    .Q(\core.csr.currentInstruction[13] ));
 sky130_fd_sc_hd__dfxtp_4 _19098_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00014_),
    .Q(\core.csr.currentInstruction[14] ));
 sky130_fd_sc_hd__dfxtp_4 _19099_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00015_),
    .Q(\core.csr.currentInstruction[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19100_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00016_),
    .Q(\core.csr.currentInstruction[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19101_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00017_),
    .Q(\core.csr.currentInstruction[17] ));
 sky130_fd_sc_hd__dfxtp_2 _19102_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00018_),
    .Q(\core.csr.currentInstruction[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19103_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00019_),
    .Q(\core.csr.currentInstruction[19] ));
 sky130_fd_sc_hd__dfxtp_4 _19104_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00020_),
    .Q(\core.csr.currentInstruction[20] ));
 sky130_fd_sc_hd__dfxtp_4 _19105_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00021_),
    .Q(\core.csr.currentInstruction[21] ));
 sky130_fd_sc_hd__dfxtp_4 _19106_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00022_),
    .Q(\core.csr.currentInstruction[22] ));
 sky130_fd_sc_hd__dfxtp_4 _19107_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_00023_),
    .Q(\core.csr.currentInstruction[23] ));
 sky130_fd_sc_hd__dfxtp_4 _19108_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00024_),
    .Q(\core.csr.currentInstruction[24] ));
 sky130_fd_sc_hd__dfxtp_4 _19109_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00025_),
    .Q(\core.csr.currentInstruction[25] ));
 sky130_fd_sc_hd__dfxtp_4 _19110_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00026_),
    .Q(\core.csr.currentInstruction[26] ));
 sky130_fd_sc_hd__dfxtp_4 _19111_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00027_),
    .Q(\core.csr.currentInstruction[27] ));
 sky130_fd_sc_hd__dfxtp_4 _19112_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00028_),
    .Q(\core.csr.currentInstruction[28] ));
 sky130_fd_sc_hd__dfxtp_4 _19113_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00029_),
    .Q(\core.csr.currentInstruction[29] ));
 sky130_fd_sc_hd__dfxtp_4 _19114_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00030_),
    .Q(\core.csr.currentInstruction[30] ));
 sky130_fd_sc_hd__dfxtp_4 _19115_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00031_),
    .Q(\core.csr.currentInstruction[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19116_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00032_),
    .Q(\core.pipe1_operation.currentPipeStall ));
 sky130_fd_sc_hd__dfxtp_4 _19117_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00033_),
    .Q(\core.csr.instruction_memoryAddress[0] ));
 sky130_fd_sc_hd__dfxtp_4 _19118_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00034_),
    .Q(\core.csr.instruction_memoryAddress[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19119_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00035_),
    .Q(\core.csr.instruction_memoryAddress[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19120_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00036_),
    .Q(\core.csr.instruction_memoryAddress[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19121_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00037_),
    .Q(\core.csr.instruction_memoryAddress[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19122_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00038_),
    .Q(\core.csr.instruction_memoryAddress[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19123_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00039_),
    .Q(\core.csr.instruction_memoryAddress[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19124_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00040_),
    .Q(\core.csr.instruction_memoryAddress[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19125_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00041_),
    .Q(\core.csr.instruction_memoryAddress[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19126_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00042_),
    .Q(\core.csr.instruction_memoryAddress[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19127_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_00043_),
    .Q(\core.csr.instruction_memoryAddress[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19128_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00044_),
    .Q(\core.csr.instruction_memoryAddress[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19129_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_00045_),
    .Q(\core.csr.instruction_memoryAddress[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19130_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_00046_),
    .Q(\core.csr.instruction_memoryAddress[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19131_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_00047_),
    .Q(\core.csr.instruction_memoryAddress[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19132_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_00048_),
    .Q(\core.csr.instruction_memoryAddress[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19133_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00049_),
    .Q(\core.csr.instruction_memoryAddress[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19134_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00050_),
    .Q(\core.csr.instruction_memoryAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19135_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00051_),
    .Q(\core.csr.instruction_memoryAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19136_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00052_),
    .Q(\core.csr.instruction_memoryAddress[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19137_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00053_),
    .Q(\core.csr.instruction_memoryAddress[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19138_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00054_),
    .Q(\core.csr.instruction_memoryAddress[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19139_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_00055_),
    .Q(\core.csr.instruction_memoryAddress[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19140_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00056_),
    .Q(\core.csr.instruction_memoryAddress[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19141_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00057_),
    .Q(\core.csr.instruction_memoryAddress[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19142_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00058_),
    .Q(\core.csr.instruction_memoryAddress[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19143_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00059_),
    .Q(\core.csr.instruction_memoryAddress[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19144_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_00060_),
    .Q(\core.csr.instruction_memoryAddress[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19145_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00061_),
    .Q(\core.csr.instruction_memoryAddress[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19146_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_00062_),
    .Q(\core.csr.instruction_memoryAddress[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19147_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_00063_),
    .Q(\core.csr.instruction_memoryAddress[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19148_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_00064_),
    .Q(\core.csr.instruction_memoryAddress[31] ));
 sky130_fd_sc_hd__dfxtp_2 _19149_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00065_),
    .Q(\core.pipe0_fetch.currentPipeStall ));
 sky130_fd_sc_hd__dfxtp_2 _19150_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00066_),
    .Q(\core.pipe0_currentInstruction[0] ));
 sky130_fd_sc_hd__dfxtp_2 _19151_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00067_),
    .Q(\core.pipe0_currentInstruction[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19152_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00068_),
    .Q(\core.pipe0_currentInstruction[2] ));
 sky130_fd_sc_hd__dfxtp_4 _19153_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00069_),
    .Q(\core.pipe0_currentInstruction[3] ));
 sky130_fd_sc_hd__dfxtp_4 _19154_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00070_),
    .Q(\core.pipe0_currentInstruction[4] ));
 sky130_fd_sc_hd__dfxtp_4 _19155_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00071_),
    .Q(\core.pipe0_currentInstruction[5] ));
 sky130_fd_sc_hd__dfxtp_4 _19156_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00072_),
    .Q(\core.pipe0_currentInstruction[6] ));
 sky130_fd_sc_hd__dfxtp_4 _19157_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00073_),
    .Q(\core.pipe0_currentInstruction[7] ));
 sky130_fd_sc_hd__dfxtp_4 _19158_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00074_),
    .Q(\core.pipe0_currentInstruction[8] ));
 sky130_fd_sc_hd__dfxtp_4 _19159_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00075_),
    .Q(\core.pipe0_currentInstruction[9] ));
 sky130_fd_sc_hd__dfxtp_4 _19160_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00076_),
    .Q(\core.pipe0_currentInstruction[10] ));
 sky130_fd_sc_hd__dfxtp_4 _19161_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00077_),
    .Q(\core.pipe0_currentInstruction[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19162_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00078_),
    .Q(\core.pipe0_currentInstruction[12] ));
 sky130_fd_sc_hd__dfxtp_4 _19163_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00079_),
    .Q(\core.pipe0_currentInstruction[13] ));
 sky130_fd_sc_hd__dfxtp_4 _19164_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00080_),
    .Q(\core.pipe0_currentInstruction[14] ));
 sky130_fd_sc_hd__dfxtp_4 _19165_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00081_),
    .Q(\core.pipe0_currentInstruction[15] ));
 sky130_fd_sc_hd__dfxtp_4 _19166_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00082_),
    .Q(\core.pipe0_currentInstruction[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19167_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00083_),
    .Q(\core.pipe0_currentInstruction[17] ));
 sky130_fd_sc_hd__dfxtp_4 _19168_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00084_),
    .Q(\core.pipe0_currentInstruction[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19169_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00085_),
    .Q(\core.pipe0_currentInstruction[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19170_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00086_),
    .Q(\core.pipe0_currentInstruction[20] ));
 sky130_fd_sc_hd__dfxtp_4 _19171_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00087_),
    .Q(\core.pipe0_currentInstruction[21] ));
 sky130_fd_sc_hd__dfxtp_4 _19172_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00088_),
    .Q(\core.pipe0_currentInstruction[22] ));
 sky130_fd_sc_hd__dfxtp_4 _19173_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00089_),
    .Q(\core.pipe0_currentInstruction[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19174_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00090_),
    .Q(\core.pipe0_currentInstruction[24] ));
 sky130_fd_sc_hd__dfxtp_4 _19175_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00091_),
    .Q(\core.pipe0_currentInstruction[25] ));
 sky130_fd_sc_hd__dfxtp_4 _19176_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00092_),
    .Q(\core.pipe0_currentInstruction[26] ));
 sky130_fd_sc_hd__dfxtp_4 _19177_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00093_),
    .Q(\core.pipe0_currentInstruction[27] ));
 sky130_fd_sc_hd__dfxtp_2 _19178_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00094_),
    .Q(\core.pipe0_currentInstruction[28] ));
 sky130_fd_sc_hd__dfxtp_4 _19179_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00095_),
    .Q(\core.pipe0_currentInstruction[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19180_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00096_),
    .Q(\core.pipe0_currentInstruction[30] ));
 sky130_fd_sc_hd__dfxtp_4 _19181_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00097_),
    .Q(\core.pipe0_currentInstruction[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19182_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00098_),
    .Q(\core.pipe0_fetch.cachedInstruction[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19183_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00099_),
    .Q(\core.pipe0_fetch.cachedInstruction[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19184_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00100_),
    .Q(\core.pipe0_fetch.cachedInstruction[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19185_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00101_),
    .Q(\core.pipe0_fetch.cachedInstruction[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19186_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00102_),
    .Q(\core.pipe0_fetch.cachedInstruction[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19187_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00103_),
    .Q(\core.pipe0_fetch.cachedInstruction[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19188_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00104_),
    .Q(\core.pipe0_fetch.cachedInstruction[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19189_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00105_),
    .Q(\core.pipe0_fetch.cachedInstruction[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19190_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00106_),
    .Q(\core.pipe0_fetch.cachedInstruction[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19191_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00107_),
    .Q(\core.pipe0_fetch.cachedInstruction[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19192_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00108_),
    .Q(\core.pipe0_fetch.cachedInstruction[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19193_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00109_),
    .Q(\core.pipe0_fetch.cachedInstruction[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19194_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00110_),
    .Q(\core.pipe0_fetch.cachedInstruction[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19195_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00111_),
    .Q(\core.pipe0_fetch.cachedInstruction[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19196_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00112_),
    .Q(\core.pipe0_fetch.cachedInstruction[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19197_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00113_),
    .Q(\core.pipe0_fetch.cachedInstruction[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19198_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00114_),
    .Q(\core.pipe0_fetch.cachedInstruction[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19199_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00115_),
    .Q(\core.pipe0_fetch.cachedInstruction[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19200_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00116_),
    .Q(\core.pipe0_fetch.cachedInstruction[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19201_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00117_),
    .Q(\core.pipe0_fetch.cachedInstruction[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19202_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00118_),
    .Q(\core.pipe0_fetch.cachedInstruction[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19203_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00119_),
    .Q(\core.pipe0_fetch.cachedInstruction[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19204_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_00120_),
    .Q(\core.pipe0_fetch.cachedInstruction[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19205_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00121_),
    .Q(\core.pipe0_fetch.cachedInstruction[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19206_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00122_),
    .Q(\core.pipe0_fetch.cachedInstruction[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19207_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00123_),
    .Q(\core.pipe0_fetch.cachedInstruction[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19208_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00124_),
    .Q(\core.pipe0_fetch.cachedInstruction[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19209_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00125_),
    .Q(\core.pipe0_fetch.cachedInstruction[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19210_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00126_),
    .Q(\core.pipe0_fetch.cachedInstruction[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19211_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_00127_),
    .Q(\core.pipe0_fetch.cachedInstruction[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19212_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00128_),
    .Q(\core.pipe0_fetch.cachedInstruction[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19213_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00129_),
    .Q(\core.pipe0_fetch.cachedInstruction[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19214_ (.CLK(clknet_4_12__leaf_wb_clk_i),
    .D(_00130_),
    .Q(\core.pipe0_fetch.instructionCached ));
 sky130_fd_sc_hd__dfxtp_2 _19215_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_00131_),
    .Q(\core.fetchProgramCounter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _19216_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_00132_),
    .Q(\core.fetchProgramCounter[1] ));
 sky130_fd_sc_hd__dfxtp_4 _19217_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_00133_),
    .Q(\core.fetchProgramCounter[2] ));
 sky130_fd_sc_hd__dfxtp_4 _19218_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_00134_),
    .Q(\core.fetchProgramCounter[3] ));
 sky130_fd_sc_hd__dfxtp_4 _19219_ (.CLK(clknet_leaf_135_wb_clk_i),
    .D(_00135_),
    .Q(\core.fetchProgramCounter[4] ));
 sky130_fd_sc_hd__dfxtp_4 _19220_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00136_),
    .Q(\core.fetchProgramCounter[5] ));
 sky130_fd_sc_hd__dfxtp_4 _19221_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00137_),
    .Q(\core.fetchProgramCounter[6] ));
 sky130_fd_sc_hd__dfxtp_4 _19222_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00138_),
    .Q(\core.fetchProgramCounter[7] ));
 sky130_fd_sc_hd__dfxtp_2 _19223_ (.CLK(clknet_leaf_137_wb_clk_i),
    .D(_00139_),
    .Q(\core.fetchProgramCounter[8] ));
 sky130_fd_sc_hd__dfxtp_4 _19224_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00140_),
    .Q(\core.fetchProgramCounter[9] ));
 sky130_fd_sc_hd__dfxtp_4 _19225_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00141_),
    .Q(\core.fetchProgramCounter[10] ));
 sky130_fd_sc_hd__dfxtp_2 _19226_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00142_),
    .Q(\core.fetchProgramCounter[11] ));
 sky130_fd_sc_hd__dfxtp_4 _19227_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00143_),
    .Q(\core.fetchProgramCounter[12] ));
 sky130_fd_sc_hd__dfxtp_4 _19228_ (.CLK(clknet_leaf_143_wb_clk_i),
    .D(_00144_),
    .Q(\core.fetchProgramCounter[13] ));
 sky130_fd_sc_hd__dfxtp_4 _19229_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00145_),
    .Q(\core.fetchProgramCounter[14] ));
 sky130_fd_sc_hd__dfxtp_4 _19230_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00146_),
    .Q(\core.fetchProgramCounter[15] ));
 sky130_fd_sc_hd__dfxtp_2 _19231_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_00147_),
    .Q(\core.fetchProgramCounter[16] ));
 sky130_fd_sc_hd__dfxtp_2 _19232_ (.CLK(clknet_leaf_145_wb_clk_i),
    .D(_00148_),
    .Q(\core.fetchProgramCounter[17] ));
 sky130_fd_sc_hd__dfxtp_2 _19233_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00149_),
    .Q(\core.fetchProgramCounter[18] ));
 sky130_fd_sc_hd__dfxtp_2 _19234_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_00150_),
    .Q(\core.fetchProgramCounter[19] ));
 sky130_fd_sc_hd__dfxtp_4 _19235_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00151_),
    .Q(\core.fetchProgramCounter[20] ));
 sky130_fd_sc_hd__dfxtp_4 _19236_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00152_),
    .Q(\core.fetchProgramCounter[21] ));
 sky130_fd_sc_hd__dfxtp_4 _19237_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00153_),
    .Q(\core.fetchProgramCounter[22] ));
 sky130_fd_sc_hd__dfxtp_4 _19238_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00154_),
    .Q(\core.fetchProgramCounter[23] ));
 sky130_fd_sc_hd__dfxtp_4 _19239_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00155_),
    .Q(\core.fetchProgramCounter[24] ));
 sky130_fd_sc_hd__dfxtp_4 _19240_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00156_),
    .Q(\core.fetchProgramCounter[25] ));
 sky130_fd_sc_hd__dfxtp_4 _19241_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00157_),
    .Q(\core.fetchProgramCounter[26] ));
 sky130_fd_sc_hd__dfxtp_2 _19242_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_00158_),
    .Q(\core.fetchProgramCounter[27] ));
 sky130_fd_sc_hd__dfxtp_4 _19243_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00159_),
    .Q(\core.fetchProgramCounter[28] ));
 sky130_fd_sc_hd__dfxtp_4 _19244_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00160_),
    .Q(\core.fetchProgramCounter[29] ));
 sky130_fd_sc_hd__dfxtp_4 _19245_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00161_),
    .Q(\core.fetchProgramCounter[30] ));
 sky130_fd_sc_hd__dfxtp_4 _19246_ (.CLK(clknet_leaf_178_wb_clk_i),
    .D(_00162_),
    .Q(\core.fetchProgramCounter[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19247_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00163_),
    .Q(\jtag.managementAddress[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19248_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00164_),
    .Q(\jtag.managementAddress[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19249_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00165_),
    .Q(\jtag.managementAddress[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19250_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00166_),
    .Q(\jtag.managementAddress[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19251_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_00167_),
    .Q(\jtag.managementAddress[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19252_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00168_),
    .Q(\jtag.managementAddress[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19253_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00169_),
    .Q(\jtag.managementAddress[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19254_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_00170_),
    .Q(\jtag.managementAddress[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19255_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00171_),
    .Q(\jtag.managementAddress[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19256_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00172_),
    .Q(\jtag.managementAddress[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19257_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_00173_),
    .Q(\jtag.managementAddress[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19258_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00174_),
    .Q(\jtag.managementAddress[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19259_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00175_),
    .Q(\jtag.managementAddress[12] ));
 sky130_fd_sc_hd__dfxtp_2 _19260_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00176_),
    .Q(\jtag.managementAddress[13] ));
 sky130_fd_sc_hd__dfxtp_4 _19261_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_00177_),
    .Q(\jtag.managementAddress[14] ));
 sky130_fd_sc_hd__dfxtp_2 _19262_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00178_),
    .Q(\jtag.managementAddress[15] ));
 sky130_fd_sc_hd__dfxtp_2 _19263_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00179_),
    .Q(\jtag.managementAddress[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19264_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_00180_),
    .Q(\jtag.managementAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19265_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_00181_),
    .Q(\jtag.managementAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19266_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_00182_),
    .Q(\jtag.managementAddress[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19267_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00183_),
    .Q(\core.registers[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19268_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00184_),
    .Q(\core.registers[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19269_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00185_),
    .Q(\core.registers[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19270_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00186_),
    .Q(\core.registers[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19271_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00187_),
    .Q(\core.registers[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19272_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00188_),
    .Q(\core.registers[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19273_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00189_),
    .Q(\core.registers[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19274_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00190_),
    .Q(\core.registers[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19275_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_00191_),
    .Q(\core.registers[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19276_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_00192_),
    .Q(\core.registers[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19277_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_00193_),
    .Q(\core.registers[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19278_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00194_),
    .Q(\core.registers[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19279_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00195_),
    .Q(\core.registers[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19280_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00196_),
    .Q(\core.registers[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19281_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00197_),
    .Q(\core.registers[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19282_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00198_),
    .Q(\core.registers[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19283_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_00199_),
    .Q(\core.registers[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19284_ (.CLK(clknet_leaf_203_wb_clk_i),
    .D(_00200_),
    .Q(\core.registers[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19285_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00201_),
    .Q(\core.registers[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19286_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00202_),
    .Q(\core.registers[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19287_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_00203_),
    .Q(\core.registers[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19288_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_00204_),
    .Q(\core.registers[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19289_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00205_),
    .Q(\core.registers[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19290_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00206_),
    .Q(\core.registers[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19291_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00207_),
    .Q(\core.registers[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19292_ (.CLK(clknet_leaf_212_wb_clk_i),
    .D(_00208_),
    .Q(\core.registers[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19293_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00209_),
    .Q(\core.registers[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19294_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00210_),
    .Q(\core.registers[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19295_ (.CLK(clknet_leaf_203_wb_clk_i),
    .D(_00211_),
    .Q(\core.registers[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19296_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00212_),
    .Q(\core.registers[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19297_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00213_),
    .Q(\core.registers[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19298_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_00214_),
    .Q(\core.registers[20][31] ));
 sky130_fd_sc_hd__dfxtp_2 _19299_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00215_),
    .Q(\core.memoryOperationCompleted ));
 sky130_fd_sc_hd__dfxtp_1 _19300_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00216_),
    .Q(\core.useCachedLoad ));
 sky130_fd_sc_hd__dfxtp_1 _19301_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_00217_),
    .Q(\core.management_pipeStartup ));
 sky130_fd_sc_hd__dfxtp_1 _19302_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00218_),
    .Q(\core.registers[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19303_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00219_),
    .Q(\core.registers[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19304_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00220_),
    .Q(\core.registers[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19305_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00221_),
    .Q(\core.registers[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19306_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00222_),
    .Q(\core.registers[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19307_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00223_),
    .Q(\core.registers[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19308_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00224_),
    .Q(\core.registers[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19309_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00225_),
    .Q(\core.registers[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19310_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00226_),
    .Q(\core.registers[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19311_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00227_),
    .Q(\core.registers[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19312_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00228_),
    .Q(\core.registers[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19313_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00229_),
    .Q(\core.registers[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19314_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00230_),
    .Q(\core.registers[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19315_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_00231_),
    .Q(\core.registers[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19316_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00232_),
    .Q(\core.registers[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19317_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00233_),
    .Q(\core.registers[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19318_ (.CLK(clknet_leaf_206_wb_clk_i),
    .D(_00234_),
    .Q(\core.registers[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19319_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_00235_),
    .Q(\core.registers[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19320_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00236_),
    .Q(\core.registers[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19321_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00237_),
    .Q(\core.registers[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19322_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00238_),
    .Q(\core.registers[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19323_ (.CLK(clknet_leaf_204_wb_clk_i),
    .D(_00239_),
    .Q(\core.registers[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19324_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00240_),
    .Q(\core.registers[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19325_ (.CLK(clknet_leaf_212_wb_clk_i),
    .D(_00241_),
    .Q(\core.registers[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19326_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00242_),
    .Q(\core.registers[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19327_ (.CLK(clknet_leaf_212_wb_clk_i),
    .D(_00243_),
    .Q(\core.registers[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19328_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00244_),
    .Q(\core.registers[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19329_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00245_),
    .Q(\core.registers[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19330_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00246_),
    .Q(\core.registers[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19331_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00247_),
    .Q(\core.registers[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19332_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00248_),
    .Q(\core.registers[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19333_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00249_),
    .Q(\core.registers[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19334_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00250_),
    .Q(\core.registers[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19335_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00251_),
    .Q(\core.registers[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19336_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00252_),
    .Q(\core.registers[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19337_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00253_),
    .Q(\core.registers[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19338_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00254_),
    .Q(\core.registers[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19339_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00255_),
    .Q(\core.registers[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19340_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00256_),
    .Q(\core.registers[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19341_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00257_),
    .Q(\core.registers[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19342_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00258_),
    .Q(\core.registers[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19343_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00259_),
    .Q(\core.registers[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19344_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00260_),
    .Q(\core.registers[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19345_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00261_),
    .Q(\core.registers[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19346_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00262_),
    .Q(\core.registers[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19347_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00263_),
    .Q(\core.registers[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19348_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00264_),
    .Q(\core.registers[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19349_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00265_),
    .Q(\core.registers[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19350_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_00266_),
    .Q(\core.registers[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19351_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00267_),
    .Q(\core.registers[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19352_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_00268_),
    .Q(\core.registers[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19353_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00269_),
    .Q(\core.registers[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19354_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00270_),
    .Q(\core.registers[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19355_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_00271_),
    .Q(\core.registers[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19356_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00272_),
    .Q(\core.registers[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19357_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00273_),
    .Q(\core.registers[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19358_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00274_),
    .Q(\core.registers[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19359_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_00275_),
    .Q(\core.registers[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19360_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_00276_),
    .Q(\core.registers[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19361_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00277_),
    .Q(\core.registers[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19362_ (.CLK(clknet_leaf_208_wb_clk_i),
    .D(_00278_),
    .Q(\core.registers[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19363_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00279_),
    .Q(\core.registers[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19364_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00280_),
    .Q(\core.registers[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19365_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00281_),
    .Q(\core.registers[30][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19366_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00282_),
    .Q(\core.registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19367_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00283_),
    .Q(\core.registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19368_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_00284_),
    .Q(\core.registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19369_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00285_),
    .Q(\core.registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19370_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00286_),
    .Q(\core.registers[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19371_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00287_),
    .Q(\core.registers[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19372_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00288_),
    .Q(\core.registers[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19373_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_00289_),
    .Q(\core.registers[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19374_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00290_),
    .Q(\core.registers[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19375_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00291_),
    .Q(\core.registers[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19376_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00292_),
    .Q(\core.registers[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19377_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_00293_),
    .Q(\core.registers[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19378_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00294_),
    .Q(\core.registers[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19379_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00295_),
    .Q(\core.registers[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19380_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_00296_),
    .Q(\core.registers[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19381_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_00297_),
    .Q(\core.registers[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19382_ (.CLK(clknet_leaf_206_wb_clk_i),
    .D(_00298_),
    .Q(\core.registers[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19383_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_00299_),
    .Q(\core.registers[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19384_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_00300_),
    .Q(\core.registers[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19385_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00301_),
    .Q(\core.registers[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19386_ (.CLK(clknet_leaf_208_wb_clk_i),
    .D(_00302_),
    .Q(\core.registers[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19387_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_00303_),
    .Q(\core.registers[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19388_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00304_),
    .Q(\core.registers[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19389_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00305_),
    .Q(\core.registers[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19390_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_00306_),
    .Q(\core.registers[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19391_ (.CLK(clknet_leaf_211_wb_clk_i),
    .D(_00307_),
    .Q(\core.registers[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19392_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_00308_),
    .Q(\core.registers[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19393_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00309_),
    .Q(\core.registers[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19394_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_00310_),
    .Q(\core.registers[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19395_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_00311_),
    .Q(\core.registers[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19396_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00312_),
    .Q(\core.registers[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19397_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_00313_),
    .Q(\core.registers[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19398_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00314_),
    .Q(\core.registers[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19399_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00315_),
    .Q(\core.registers[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19400_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00316_),
    .Q(\core.registers[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19401_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00317_),
    .Q(\core.registers[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19402_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00318_),
    .Q(\core.registers[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19403_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00319_),
    .Q(\core.registers[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19404_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00320_),
    .Q(\core.registers[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19405_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00321_),
    .Q(\core.registers[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19406_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00322_),
    .Q(\core.registers[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19407_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00323_),
    .Q(\core.registers[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19408_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00324_),
    .Q(\core.registers[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19409_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00325_),
    .Q(\core.registers[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19410_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00326_),
    .Q(\core.registers[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19411_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00327_),
    .Q(\core.registers[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19412_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_00328_),
    .Q(\core.registers[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19413_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00329_),
    .Q(\core.registers[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19414_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_00330_),
    .Q(\core.registers[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19415_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00331_),
    .Q(\core.registers[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19416_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00332_),
    .Q(\core.registers[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19417_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00333_),
    .Q(\core.registers[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19418_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_00334_),
    .Q(\core.registers[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19419_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_00335_),
    .Q(\core.registers[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19420_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00336_),
    .Q(\core.registers[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19421_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00337_),
    .Q(\core.registers[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19422_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00338_),
    .Q(\core.registers[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19423_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_00339_),
    .Q(\core.registers[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19424_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00340_),
    .Q(\core.registers[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19425_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00341_),
    .Q(\core.registers[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19426_ (.CLK(clknet_leaf_208_wb_clk_i),
    .D(_00342_),
    .Q(\core.registers[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19427_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00343_),
    .Q(\core.registers[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19428_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00344_),
    .Q(\core.registers[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19429_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00345_),
    .Q(\core.registers[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19430_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00346_),
    .Q(\core.registers[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19431_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00347_),
    .Q(\core.registers[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19432_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00348_),
    .Q(\core.registers[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19433_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00349_),
    .Q(\core.registers[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19434_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00350_),
    .Q(\core.registers[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19435_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00351_),
    .Q(\core.registers[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19436_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00352_),
    .Q(\core.registers[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19437_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00353_),
    .Q(\core.registers[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19438_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00354_),
    .Q(\core.registers[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19439_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_00355_),
    .Q(\core.registers[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19440_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00356_),
    .Q(\core.registers[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19441_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00357_),
    .Q(\core.registers[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19442_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00358_),
    .Q(\core.registers[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19443_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00359_),
    .Q(\core.registers[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19444_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00360_),
    .Q(\core.registers[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19445_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00361_),
    .Q(\core.registers[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19446_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_00362_),
    .Q(\core.registers[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19447_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00363_),
    .Q(\core.registers[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19448_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00364_),
    .Q(\core.registers[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19449_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00365_),
    .Q(\core.registers[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19450_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00366_),
    .Q(\core.registers[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19451_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_00367_),
    .Q(\core.registers[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19452_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00368_),
    .Q(\core.registers[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19453_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00369_),
    .Q(\core.registers[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19454_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00370_),
    .Q(\core.registers[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19455_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00371_),
    .Q(\core.registers[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19456_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00372_),
    .Q(\core.registers[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19457_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00373_),
    .Q(\core.registers[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19458_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00374_),
    .Q(\core.registers[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19459_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00375_),
    .Q(\core.registers[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19460_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00376_),
    .Q(\core.registers[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19461_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00377_),
    .Q(\core.registers[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19462_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00378_),
    .Q(\core.registers[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19463_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00379_),
    .Q(\core.registers[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19464_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00380_),
    .Q(\core.registers[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19465_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00381_),
    .Q(\core.registers[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19466_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00382_),
    .Q(\core.registers[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19467_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_00383_),
    .Q(\core.registers[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19468_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00384_),
    .Q(\core.registers[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19469_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00385_),
    .Q(\core.registers[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19470_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00386_),
    .Q(\core.registers[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19471_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_00387_),
    .Q(\core.registers[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19472_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00388_),
    .Q(\core.registers[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19473_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00389_),
    .Q(\core.registers[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19474_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00390_),
    .Q(\core.registers[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19475_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00391_),
    .Q(\core.registers[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19476_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00392_),
    .Q(\core.registers[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19477_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00393_),
    .Q(\core.registers[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19478_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00394_),
    .Q(\core.registers[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19479_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00395_),
    .Q(\core.registers[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19480_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00396_),
    .Q(\core.registers[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19481_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00397_),
    .Q(\core.registers[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19482_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00398_),
    .Q(\core.registers[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19483_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_00399_),
    .Q(\core.registers[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19484_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00400_),
    .Q(\core.registers[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19485_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00401_),
    .Q(\core.registers[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19486_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00402_),
    .Q(\core.registers[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19487_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00403_),
    .Q(\core.registers[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19488_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00404_),
    .Q(\core.registers[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19489_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00405_),
    .Q(\core.registers[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19490_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00406_),
    .Q(\core.registers[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19491_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00407_),
    .Q(\core.registers[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19492_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00408_),
    .Q(\core.registers[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19493_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00409_),
    .Q(\core.registers[26][31] ));
 sky130_fd_sc_hd__dfxtp_4 _19494_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_00410_),
    .Q(net450));
 sky130_fd_sc_hd__dfxtp_4 _19495_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_00411_),
    .Q(net461));
 sky130_fd_sc_hd__dfxtp_4 _19496_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00412_),
    .Q(net472));
 sky130_fd_sc_hd__dfxtp_4 _19497_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00413_),
    .Q(net475));
 sky130_fd_sc_hd__dfxtp_4 _19498_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_00414_),
    .Q(net476));
 sky130_fd_sc_hd__dfxtp_4 _19499_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00415_),
    .Q(net477));
 sky130_fd_sc_hd__dfxtp_4 _19500_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_00416_),
    .Q(net478));
 sky130_fd_sc_hd__dfxtp_4 _19501_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00417_),
    .Q(net479));
 sky130_fd_sc_hd__dfxtp_4 _19502_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_00418_),
    .Q(net480));
 sky130_fd_sc_hd__dfxtp_4 _19503_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_00419_),
    .Q(net481));
 sky130_fd_sc_hd__dfxtp_4 _19504_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_00420_),
    .Q(net451));
 sky130_fd_sc_hd__dfxtp_4 _19505_ (.CLK(clknet_leaf_142_wb_clk_i),
    .D(_00421_),
    .Q(net452));
 sky130_fd_sc_hd__dfxtp_4 _19506_ (.CLK(clknet_leaf_149_wb_clk_i),
    .D(_00422_),
    .Q(net453));
 sky130_fd_sc_hd__dfxtp_4 _19507_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_00423_),
    .Q(net454));
 sky130_fd_sc_hd__dfxtp_4 _19508_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_00424_),
    .Q(net455));
 sky130_fd_sc_hd__dfxtp_4 _19509_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_00425_),
    .Q(net456));
 sky130_fd_sc_hd__dfxtp_4 _19510_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00426_),
    .Q(net457));
 sky130_fd_sc_hd__dfxtp_4 _19511_ (.CLK(clknet_leaf_146_wb_clk_i),
    .D(_00427_),
    .Q(net458));
 sky130_fd_sc_hd__dfxtp_4 _19512_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_00428_),
    .Q(net459));
 sky130_fd_sc_hd__dfxtp_4 _19513_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_00429_),
    .Q(net460));
 sky130_fd_sc_hd__dfxtp_4 _19514_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_00430_),
    .Q(net462));
 sky130_fd_sc_hd__dfxtp_4 _19515_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_00431_),
    .Q(net463));
 sky130_fd_sc_hd__dfxtp_4 _19516_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_00432_),
    .Q(net464));
 sky130_fd_sc_hd__dfxtp_4 _19517_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00433_),
    .Q(net465));
 sky130_fd_sc_hd__dfxtp_4 _19518_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_00434_),
    .Q(net466));
 sky130_fd_sc_hd__dfxtp_4 _19519_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_00435_),
    .Q(net467));
 sky130_fd_sc_hd__dfxtp_4 _19520_ (.CLK(clknet_leaf_177_wb_clk_i),
    .D(_00436_),
    .Q(net468));
 sky130_fd_sc_hd__dfxtp_4 _19521_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_00437_),
    .Q(net469));
 sky130_fd_sc_hd__dfxtp_4 _19522_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00438_),
    .Q(net470));
 sky130_fd_sc_hd__dfxtp_4 _19523_ (.CLK(clknet_leaf_189_wb_clk_i),
    .D(_00439_),
    .Q(net471));
 sky130_fd_sc_hd__dfxtp_4 _19524_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_00440_),
    .Q(net473));
 sky130_fd_sc_hd__dfxtp_4 _19525_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_00441_),
    .Q(net474));
 sky130_fd_sc_hd__dfxtp_1 _19526_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00442_),
    .Q(\core.cancelStall ));
 sky130_fd_sc_hd__dfxtp_4 _19527_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00443_),
    .Q(\core.pipe1_resultRegister[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19528_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00444_),
    .Q(\core.pipe1_resultRegister[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19529_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00445_),
    .Q(\core.pipe1_resultRegister[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19530_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00446_),
    .Q(\core.pipe1_resultRegister[3] ));
 sky130_fd_sc_hd__dfxtp_2 _19531_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00447_),
    .Q(\core.pipe1_resultRegister[4] ));
 sky130_fd_sc_hd__dfxtp_2 _19532_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00448_),
    .Q(\core.pipe1_resultRegister[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19533_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00449_),
    .Q(\core.pipe1_resultRegister[6] ));
 sky130_fd_sc_hd__dfxtp_2 _19534_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00450_),
    .Q(\core.pipe1_resultRegister[7] ));
 sky130_fd_sc_hd__dfxtp_2 _19535_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00451_),
    .Q(\core.pipe1_resultRegister[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19536_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00452_),
    .Q(\core.pipe1_resultRegister[9] ));
 sky130_fd_sc_hd__dfxtp_4 _19537_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00453_),
    .Q(\core.pipe1_resultRegister[10] ));
 sky130_fd_sc_hd__dfxtp_2 _19538_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00454_),
    .Q(\core.pipe1_resultRegister[11] ));
 sky130_fd_sc_hd__dfxtp_4 _19539_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00455_),
    .Q(\core.pipe1_resultRegister[12] ));
 sky130_fd_sc_hd__dfxtp_4 _19540_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00456_),
    .Q(\core.pipe1_resultRegister[13] ));
 sky130_fd_sc_hd__dfxtp_4 _19541_ (.CLK(clknet_leaf_193_wb_clk_i),
    .D(_00457_),
    .Q(\core.pipe1_resultRegister[14] ));
 sky130_fd_sc_hd__dfxtp_4 _19542_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_00458_),
    .Q(\core.pipe1_resultRegister[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19543_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_00459_),
    .Q(\core.pipe1_resultRegister[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19544_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00460_),
    .Q(\core.pipe1_resultRegister[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19545_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_00461_),
    .Q(\core.pipe1_resultRegister[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19546_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_00462_),
    .Q(\core.pipe1_resultRegister[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19547_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00463_),
    .Q(\core.pipe1_resultRegister[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19548_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00464_),
    .Q(\core.pipe1_resultRegister[21] ));
 sky130_fd_sc_hd__dfxtp_4 _19549_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_00465_),
    .Q(\core.pipe1_resultRegister[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19550_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_00466_),
    .Q(\core.pipe1_resultRegister[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19551_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_00467_),
    .Q(\core.pipe1_resultRegister[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19552_ (.CLK(clknet_4_1__leaf_wb_clk_i),
    .D(_00468_),
    .Q(\core.pipe1_resultRegister[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19553_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_00469_),
    .Q(\core.pipe1_resultRegister[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19554_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_00470_),
    .Q(\core.pipe1_resultRegister[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19555_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00471_),
    .Q(\core.pipe1_resultRegister[28] ));
 sky130_fd_sc_hd__dfxtp_4 _19556_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_00472_),
    .Q(\core.pipe1_resultRegister[29] ));
 sky130_fd_sc_hd__dfxtp_4 _19557_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00473_),
    .Q(\core.pipe1_resultRegister[30] ));
 sky130_fd_sc_hd__dfxtp_4 _19558_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_00474_),
    .Q(\core.pipe1_resultRegister[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19559_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00475_),
    .Q(\core.pipe1_loadResult[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19560_ (.CLK(clknet_leaf_79_wb_clk_i),
    .D(_00476_),
    .Q(\core.pipe1_loadResult[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19561_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00477_),
    .Q(\core.pipe1_loadResult[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19562_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00478_),
    .Q(\core.pipe1_loadResult[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19563_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00479_),
    .Q(\core.pipe1_loadResult[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19564_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00480_),
    .Q(\core.pipe1_loadResult[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19565_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00481_),
    .Q(\core.pipe1_loadResult[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19566_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00482_),
    .Q(\core.pipe1_loadResult[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19567_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00483_),
    .Q(\core.pipe1_loadResult[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19568_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00484_),
    .Q(\core.pipe1_loadResult[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19569_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00485_),
    .Q(\core.pipe1_loadResult[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19570_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00486_),
    .Q(\core.pipe1_loadResult[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19571_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00487_),
    .Q(\core.pipe1_loadResult[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19572_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00488_),
    .Q(\core.pipe1_loadResult[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19573_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00489_),
    .Q(\core.pipe1_loadResult[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19574_ (.CLK(clknet_leaf_89_wb_clk_i),
    .D(_00490_),
    .Q(\core.pipe1_loadResult[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19575_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00491_),
    .Q(\core.pipe1_loadResult[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19576_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00492_),
    .Q(\core.pipe1_loadResult[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19577_ (.CLK(clknet_leaf_78_wb_clk_i),
    .D(_00493_),
    .Q(\core.pipe1_loadResult[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19578_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00494_),
    .Q(\core.pipe1_loadResult[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19579_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00495_),
    .Q(\core.pipe1_loadResult[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19580_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00496_),
    .Q(\core.pipe1_loadResult[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19581_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00497_),
    .Q(\core.pipe1_loadResult[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19582_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00498_),
    .Q(\core.pipe1_loadResult[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19583_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00499_),
    .Q(\core.pipe1_loadResult[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19584_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00500_),
    .Q(\core.pipe1_loadResult[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19585_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00501_),
    .Q(\core.pipe1_loadResult[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19586_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00502_),
    .Q(\core.pipe1_loadResult[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19587_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00503_),
    .Q(\core.pipe1_loadResult[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19588_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00504_),
    .Q(\core.pipe1_loadResult[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19589_ (.CLK(clknet_leaf_91_wb_clk_i),
    .D(_00505_),
    .Q(\core.pipe1_loadResult[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19590_ (.CLK(clknet_leaf_90_wb_clk_i),
    .D(_00506_),
    .Q(\core.pipe1_loadResult[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19591_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00507_),
    .Q(\core.pipe1_csrData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19592_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00508_),
    .Q(\core.pipe1_csrData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19593_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00509_),
    .Q(\core.pipe1_csrData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19594_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00510_),
    .Q(\core.pipe1_csrData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19595_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00511_),
    .Q(\core.pipe1_csrData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19596_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00512_),
    .Q(\core.pipe1_csrData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19597_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00513_),
    .Q(\core.pipe1_csrData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _19598_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00514_),
    .Q(\core.pipe1_csrData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19599_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00515_),
    .Q(\core.pipe1_csrData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19600_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00516_),
    .Q(\core.pipe1_csrData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _19601_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00517_),
    .Q(\core.pipe1_csrData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19602_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00518_),
    .Q(\core.pipe1_csrData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19603_ (.CLK(clknet_leaf_80_wb_clk_i),
    .D(_00519_),
    .Q(\core.pipe1_csrData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _19604_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00520_),
    .Q(\core.pipe1_csrData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19605_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00521_),
    .Q(\core.pipe1_csrData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19606_ (.CLK(clknet_leaf_82_wb_clk_i),
    .D(_00522_),
    .Q(\core.pipe1_csrData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _19607_ (.CLK(clknet_leaf_192_wb_clk_i),
    .D(_00523_),
    .Q(\core.pipe1_csrData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19608_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00524_),
    .Q(\core.pipe1_csrData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19609_ (.CLK(clknet_leaf_190_wb_clk_i),
    .D(_00525_),
    .Q(\core.pipe1_csrData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _19610_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_00526_),
    .Q(\core.pipe1_csrData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19611_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00527_),
    .Q(\core.pipe1_csrData[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19612_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00528_),
    .Q(\core.pipe1_csrData[21] ));
 sky130_fd_sc_hd__dfxtp_1 _19613_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00529_),
    .Q(\core.pipe1_csrData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19614_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_00530_),
    .Q(\core.pipe1_csrData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19615_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_00531_),
    .Q(\core.pipe1_csrData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _19616_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00532_),
    .Q(\core.pipe1_csrData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19617_ (.CLK(clknet_leaf_188_wb_clk_i),
    .D(_00533_),
    .Q(\core.pipe1_csrData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19618_ (.CLK(clknet_leaf_191_wb_clk_i),
    .D(_00534_),
    .Q(\core.pipe1_csrData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _19619_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_00535_),
    .Q(\core.pipe1_csrData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19620_ (.CLK(clknet_leaf_81_wb_clk_i),
    .D(_00536_),
    .Q(\core.pipe1_csrData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19621_ (.CLK(clknet_leaf_83_wb_clk_i),
    .D(_00537_),
    .Q(\core.pipe1_csrData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _19622_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00538_),
    .Q(\core.pipe1_csrData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _19623_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00539_),
    .Q(\core.registers[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19624_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00540_),
    .Q(\core.registers[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19625_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00541_),
    .Q(\core.registers[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19626_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00542_),
    .Q(\core.registers[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19627_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00543_),
    .Q(\core.registers[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19628_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00544_),
    .Q(\core.registers[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19629_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00545_),
    .Q(\core.registers[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19630_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00546_),
    .Q(\core.registers[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19631_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_00547_),
    .Q(\core.registers[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19632_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00548_),
    .Q(\core.registers[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19633_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00549_),
    .Q(\core.registers[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19634_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00550_),
    .Q(\core.registers[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19635_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00551_),
    .Q(\core.registers[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19636_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_00552_),
    .Q(\core.registers[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19637_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00553_),
    .Q(\core.registers[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19638_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00554_),
    .Q(\core.registers[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19639_ (.CLK(clknet_leaf_206_wb_clk_i),
    .D(_00555_),
    .Q(\core.registers[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19640_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00556_),
    .Q(\core.registers[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19641_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00557_),
    .Q(\core.registers[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19642_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00558_),
    .Q(\core.registers[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19643_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_00559_),
    .Q(\core.registers[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19644_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00560_),
    .Q(\core.registers[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19645_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00561_),
    .Q(\core.registers[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19646_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00562_),
    .Q(\core.registers[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19647_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00563_),
    .Q(\core.registers[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19648_ (.CLK(clknet_leaf_211_wb_clk_i),
    .D(_00564_),
    .Q(\core.registers[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19649_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00565_),
    .Q(\core.registers[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19650_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00566_),
    .Q(\core.registers[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19651_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00567_),
    .Q(\core.registers[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19652_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00568_),
    .Q(\core.registers[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19653_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00569_),
    .Q(\core.registers[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19654_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_00570_),
    .Q(\core.registers[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19655_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00571_),
    .Q(\localMemoryInterface.lastCoreByteSelect[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19656_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00572_),
    .Q(\localMemoryInterface.lastCoreByteSelect[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19657_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00573_),
    .Q(\localMemoryInterface.lastCoreByteSelect[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19658_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_00574_),
    .Q(\localMemoryInterface.lastCoreByteSelect[3] ));
 sky130_fd_sc_hd__dfxtp_4 _19659_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00575_),
    .Q(\memoryController.last_instruction_enableLocalMemory ));
 sky130_fd_sc_hd__dfxtp_4 _19660_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00576_),
    .Q(\memoryController.last_data_enableLocalMemory ));
 sky130_fd_sc_hd__dfxtp_4 _19661_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(net728),
    .Q(\memoryController.last_instruction_enableWB ));
 sky130_fd_sc_hd__dfxtp_1 _19662_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00578_),
    .Q(\core.registers[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19663_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00579_),
    .Q(\core.registers[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19664_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00580_),
    .Q(\core.registers[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19665_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00581_),
    .Q(\core.registers[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19666_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_00582_),
    .Q(\core.registers[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19667_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00583_),
    .Q(\core.registers[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19668_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_00584_),
    .Q(\core.registers[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19669_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00585_),
    .Q(\core.registers[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19670_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_00586_),
    .Q(\core.registers[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19671_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00587_),
    .Q(\core.registers[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19672_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_00588_),
    .Q(\core.registers[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19673_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00589_),
    .Q(\core.registers[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19674_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_00590_),
    .Q(\core.registers[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19675_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_00591_),
    .Q(\core.registers[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19676_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00592_),
    .Q(\core.registers[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19677_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00593_),
    .Q(\core.registers[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19678_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_00594_),
    .Q(\core.registers[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19679_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_00595_),
    .Q(\core.registers[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19680_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_00596_),
    .Q(\core.registers[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19681_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00597_),
    .Q(\core.registers[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19682_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_00598_),
    .Q(\core.registers[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19683_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_00599_),
    .Q(\core.registers[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19684_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_00600_),
    .Q(\core.registers[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19685_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00601_),
    .Q(\core.registers[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19686_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_00602_),
    .Q(\core.registers[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19687_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_00603_),
    .Q(\core.registers[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19688_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_00604_),
    .Q(\core.registers[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19689_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_00605_),
    .Q(\core.registers[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19690_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_00606_),
    .Q(\core.registers[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19691_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00607_),
    .Q(\core.registers[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19692_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_00608_),
    .Q(\core.registers[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19693_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00609_),
    .Q(\core.registers[12][31] ));
 sky130_fd_sc_hd__dfxtp_2 _19694_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00610_),
    .Q(\localMemoryInterface.lastRBankSelect ));
 sky130_fd_sc_hd__dfxtp_4 _19695_ (.CLK(clknet_leaf_144_wb_clk_i),
    .D(_00611_),
    .Q(\localMemoryInterface.coreReadReady ));
 sky130_fd_sc_hd__dfxtp_1 _19696_ (.CLK(clknet_leaf_141_wb_clk_i),
    .D(_00612_),
    .Q(\localMemoryInterface.lastWBByteSelect[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19697_ (.CLK(clknet_leaf_140_wb_clk_i),
    .D(_00613_),
    .Q(\localMemoryInterface.lastWBByteSelect[1] ));
 sky130_fd_sc_hd__dfxtp_2 _19698_ (.CLK(clknet_leaf_138_wb_clk_i),
    .D(_00614_),
    .Q(\localMemoryInterface.lastWBByteSelect[2] ));
 sky130_fd_sc_hd__dfxtp_2 _19699_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00615_),
    .Q(\localMemoryInterface.lastWBByteSelect[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19700_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00616_),
    .Q(\localMemoryInterface.lastRWBankSelect ));
 sky130_fd_sc_hd__dfxtp_4 _19701_ (.CLK(clknet_leaf_139_wb_clk_i),
    .D(_00617_),
    .Q(\localMemoryInterface.wbReadReady ));
 sky130_fd_sc_hd__dfxtp_4 _19702_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00618_),
    .Q(\core.csr.cycleTimer.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_2 _19703_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00619_),
    .Q(\core.csr.cycleTimer.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19704_ (.CLK(clknet_leaf_88_wb_clk_i),
    .D(_00620_),
    .Q(\core.csr.cycleTimer.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _19705_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00621_),
    .Q(\core.csr.cycleTimer.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_1 _19706_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00622_),
    .Q(\core.csr.cycleTimer.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _19707_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00623_),
    .Q(\core.csr.cycleTimer.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _19708_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00624_),
    .Q(\core.csr.cycleTimer.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_2 _19709_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00625_),
    .Q(\core.csr.cycleTimer.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_1 _19710_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00626_),
    .Q(\core.csr.cycleTimer.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_1 _19711_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00627_),
    .Q(\core.csr.cycleTimer.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_2 _19712_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00628_),
    .Q(\core.csr.cycleTimer.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_1 _19713_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00629_),
    .Q(\core.csr.cycleTimer.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_1 _19714_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00630_),
    .Q(\core.csr.cycleTimer.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_2 _19715_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00631_),
    .Q(\core.csr.cycleTimer.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _19716_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00632_),
    .Q(\core.csr.cycleTimer.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _19717_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00633_),
    .Q(\core.csr.cycleTimer.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_2 _19718_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00634_),
    .Q(\core.csr.cycleTimer.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_1 _19719_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00635_),
    .Q(\core.csr.cycleTimer.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_1 _19720_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_00636_),
    .Q(\core.csr.cycleTimer.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_2 _19721_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_00637_),
    .Q(\core.csr.cycleTimer.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _19722_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_00638_),
    .Q(\core.csr.cycleTimer.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_1 _19723_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_00639_),
    .Q(\core.csr.cycleTimer.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_2 _19724_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00640_),
    .Q(\core.csr.cycleTimer.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _19725_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00641_),
    .Q(\core.csr.cycleTimer.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_1 _19726_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00642_),
    .Q(\core.csr.cycleTimer.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_2 _19727_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00643_),
    .Q(\core.csr.cycleTimer.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _19728_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00644_),
    .Q(\core.csr.cycleTimer.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_1 _19729_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00645_),
    .Q(\core.csr.cycleTimer.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_2 _19730_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00646_),
    .Q(\core.csr.cycleTimer.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_1 _19731_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_00647_),
    .Q(\core.csr.cycleTimer.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_1 _19732_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00648_),
    .Q(\core.csr.cycleTimer.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_2 _19733_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00649_),
    .Q(\core.csr.cycleTimer.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_2 _19734_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_00650_),
    .Q(\core.csr.cycleTimer.currentValue[32] ));
 sky130_fd_sc_hd__dfxtp_1 _19735_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_00651_),
    .Q(\core.csr.cycleTimer.currentValue[33] ));
 sky130_fd_sc_hd__dfxtp_2 _19736_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00652_),
    .Q(\core.csr.cycleTimer.currentValue[34] ));
 sky130_fd_sc_hd__dfxtp_1 _19737_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_00653_),
    .Q(\core.csr.cycleTimer.currentValue[35] ));
 sky130_fd_sc_hd__dfxtp_1 _19738_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00654_),
    .Q(\core.csr.cycleTimer.currentValue[36] ));
 sky130_fd_sc_hd__dfxtp_2 _19739_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_00655_),
    .Q(\core.csr.cycleTimer.currentValue[37] ));
 sky130_fd_sc_hd__dfxtp_1 _19740_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00656_),
    .Q(\core.csr.cycleTimer.currentValue[38] ));
 sky130_fd_sc_hd__dfxtp_1 _19741_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_00657_),
    .Q(\core.csr.cycleTimer.currentValue[39] ));
 sky130_fd_sc_hd__dfxtp_2 _19742_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00658_),
    .Q(\core.csr.cycleTimer.currentValue[40] ));
 sky130_fd_sc_hd__dfxtp_1 _19743_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_00659_),
    .Q(\core.csr.cycleTimer.currentValue[41] ));
 sky130_fd_sc_hd__dfxtp_1 _19744_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00660_),
    .Q(\core.csr.cycleTimer.currentValue[42] ));
 sky130_fd_sc_hd__dfxtp_2 _19745_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_00661_),
    .Q(\core.csr.cycleTimer.currentValue[43] ));
 sky130_fd_sc_hd__dfxtp_1 _19746_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_00662_),
    .Q(\core.csr.cycleTimer.currentValue[44] ));
 sky130_fd_sc_hd__dfxtp_1 _19747_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_00663_),
    .Q(\core.csr.cycleTimer.currentValue[45] ));
 sky130_fd_sc_hd__dfxtp_2 _19748_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_00664_),
    .Q(\core.csr.cycleTimer.currentValue[46] ));
 sky130_fd_sc_hd__dfxtp_1 _19749_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00665_),
    .Q(\core.csr.cycleTimer.currentValue[47] ));
 sky130_fd_sc_hd__dfxtp_1 _19750_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00666_),
    .Q(\core.csr.cycleTimer.currentValue[48] ));
 sky130_fd_sc_hd__dfxtp_2 _19751_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_00667_),
    .Q(\core.csr.cycleTimer.currentValue[49] ));
 sky130_fd_sc_hd__dfxtp_2 _19752_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00668_),
    .Q(\core.csr.cycleTimer.currentValue[50] ));
 sky130_fd_sc_hd__dfxtp_1 _19753_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_00669_),
    .Q(\core.csr.cycleTimer.currentValue[51] ));
 sky130_fd_sc_hd__dfxtp_2 _19754_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_00670_),
    .Q(\core.csr.cycleTimer.currentValue[52] ));
 sky130_fd_sc_hd__dfxtp_1 _19755_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_00671_),
    .Q(\core.csr.cycleTimer.currentValue[53] ));
 sky130_fd_sc_hd__dfxtp_1 _19756_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_00672_),
    .Q(\core.csr.cycleTimer.currentValue[54] ));
 sky130_fd_sc_hd__dfxtp_2 _19757_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_00673_),
    .Q(\core.csr.cycleTimer.currentValue[55] ));
 sky130_fd_sc_hd__dfxtp_1 _19758_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_00674_),
    .Q(\core.csr.cycleTimer.currentValue[56] ));
 sky130_fd_sc_hd__dfxtp_1 _19759_ (.CLK(clknet_leaf_155_wb_clk_i),
    .D(_00675_),
    .Q(\core.csr.cycleTimer.currentValue[57] ));
 sky130_fd_sc_hd__dfxtp_2 _19760_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00676_),
    .Q(\core.csr.cycleTimer.currentValue[58] ));
 sky130_fd_sc_hd__dfxtp_1 _19761_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00677_),
    .Q(\core.csr.cycleTimer.currentValue[59] ));
 sky130_fd_sc_hd__dfxtp_1 _19762_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00678_),
    .Q(\core.csr.cycleTimer.currentValue[60] ));
 sky130_fd_sc_hd__dfxtp_2 _19763_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00679_),
    .Q(\core.csr.cycleTimer.currentValue[61] ));
 sky130_fd_sc_hd__dfxtp_2 _19764_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00680_),
    .Q(\core.csr.cycleTimer.currentValue[62] ));
 sky130_fd_sc_hd__dfxtp_1 _19765_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00681_),
    .Q(\core.csr.cycleTimer.currentValue[63] ));
 sky130_fd_sc_hd__dfxtp_1 _19766_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00682_),
    .Q(\core.registers[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19767_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00683_),
    .Q(\core.registers[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19768_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00684_),
    .Q(\core.registers[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19769_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00685_),
    .Q(\core.registers[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19770_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00686_),
    .Q(\core.registers[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19771_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_00687_),
    .Q(\core.registers[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19772_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00688_),
    .Q(\core.registers[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19773_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00689_),
    .Q(\core.registers[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19774_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00690_),
    .Q(\core.registers[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19775_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_00691_),
    .Q(\core.registers[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19776_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00692_),
    .Q(\core.registers[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19777_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00693_),
    .Q(\core.registers[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19778_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00694_),
    .Q(\core.registers[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19779_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00695_),
    .Q(\core.registers[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19780_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00696_),
    .Q(\core.registers[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19781_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_00697_),
    .Q(\core.registers[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19782_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00698_),
    .Q(\core.registers[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19783_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00699_),
    .Q(\core.registers[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19784_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00700_),
    .Q(\core.registers[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19785_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00701_),
    .Q(\core.registers[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19786_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00702_),
    .Q(\core.registers[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19787_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_00703_),
    .Q(\core.registers[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19788_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00704_),
    .Q(\core.registers[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19789_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00705_),
    .Q(\core.registers[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19790_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00706_),
    .Q(\core.registers[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19791_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00707_),
    .Q(\core.registers[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19792_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00708_),
    .Q(\core.registers[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19793_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00709_),
    .Q(\core.registers[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19794_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00710_),
    .Q(\core.registers[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19795_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00711_),
    .Q(\core.registers[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19796_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00712_),
    .Q(\core.registers[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19797_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00713_),
    .Q(\core.registers[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19798_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00714_),
    .Q(\core.registers[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19799_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00715_),
    .Q(\core.registers[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19800_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00716_),
    .Q(\core.registers[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19801_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00717_),
    .Q(\core.registers[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19802_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00718_),
    .Q(\core.registers[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19803_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00719_),
    .Q(\core.registers[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19804_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00720_),
    .Q(\core.registers[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19805_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00721_),
    .Q(\core.registers[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19806_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_00722_),
    .Q(\core.registers[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19807_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00723_),
    .Q(\core.registers[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19808_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00724_),
    .Q(\core.registers[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19809_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00725_),
    .Q(\core.registers[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19810_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00726_),
    .Q(\core.registers[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19811_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00727_),
    .Q(\core.registers[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19812_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00728_),
    .Q(\core.registers[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19813_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00729_),
    .Q(\core.registers[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19814_ (.CLK(clknet_leaf_206_wb_clk_i),
    .D(_00730_),
    .Q(\core.registers[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19815_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_00731_),
    .Q(\core.registers[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19816_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00732_),
    .Q(\core.registers[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19817_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00733_),
    .Q(\core.registers[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19818_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00734_),
    .Q(\core.registers[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19819_ (.CLK(clknet_leaf_204_wb_clk_i),
    .D(_00735_),
    .Q(\core.registers[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19820_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00736_),
    .Q(\core.registers[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19821_ (.CLK(clknet_leaf_212_wb_clk_i),
    .D(_00737_),
    .Q(\core.registers[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19822_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00738_),
    .Q(\core.registers[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19823_ (.CLK(clknet_leaf_212_wb_clk_i),
    .D(_00739_),
    .Q(\core.registers[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19824_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00740_),
    .Q(\core.registers[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19825_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00741_),
    .Q(\core.registers[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19826_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00742_),
    .Q(\core.registers[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19827_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00743_),
    .Q(\core.registers[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19828_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00744_),
    .Q(\core.registers[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19829_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00745_),
    .Q(\core.registers[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19830_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_00746_),
    .Q(\coreWBInterface.stb ));
 sky130_fd_sc_hd__dfxtp_4 _19831_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00747_),
    .Q(\coreWBInterface.readDataBuffered[0] ));
 sky130_fd_sc_hd__dfxtp_4 _19832_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00748_),
    .Q(\coreWBInterface.readDataBuffered[1] ));
 sky130_fd_sc_hd__dfxtp_4 _19833_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00749_),
    .Q(\coreWBInterface.readDataBuffered[2] ));
 sky130_fd_sc_hd__dfxtp_4 _19834_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00750_),
    .Q(\coreWBInterface.readDataBuffered[3] ));
 sky130_fd_sc_hd__dfxtp_4 _19835_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00751_),
    .Q(\coreWBInterface.readDataBuffered[4] ));
 sky130_fd_sc_hd__dfxtp_4 _19836_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00752_),
    .Q(\coreWBInterface.readDataBuffered[5] ));
 sky130_fd_sc_hd__dfxtp_4 _19837_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00753_),
    .Q(\coreWBInterface.readDataBuffered[6] ));
 sky130_fd_sc_hd__dfxtp_4 _19838_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00754_),
    .Q(\coreWBInterface.readDataBuffered[7] ));
 sky130_fd_sc_hd__dfxtp_4 _19839_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00755_),
    .Q(\coreWBInterface.readDataBuffered[8] ));
 sky130_fd_sc_hd__dfxtp_4 _19840_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_00756_),
    .Q(\coreWBInterface.readDataBuffered[9] ));
 sky130_fd_sc_hd__dfxtp_4 _19841_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00757_),
    .Q(\coreWBInterface.readDataBuffered[10] ));
 sky130_fd_sc_hd__dfxtp_4 _19842_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00758_),
    .Q(\coreWBInterface.readDataBuffered[11] ));
 sky130_fd_sc_hd__dfxtp_4 _19843_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00759_),
    .Q(\coreWBInterface.readDataBuffered[12] ));
 sky130_fd_sc_hd__dfxtp_4 _19844_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00760_),
    .Q(\coreWBInterface.readDataBuffered[13] ));
 sky130_fd_sc_hd__dfxtp_4 _19845_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00761_),
    .Q(\coreWBInterface.readDataBuffered[14] ));
 sky130_fd_sc_hd__dfxtp_4 _19846_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00762_),
    .Q(\coreWBInterface.readDataBuffered[15] ));
 sky130_fd_sc_hd__dfxtp_4 _19847_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00763_),
    .Q(\coreWBInterface.readDataBuffered[16] ));
 sky130_fd_sc_hd__dfxtp_4 _19848_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00764_),
    .Q(\coreWBInterface.readDataBuffered[17] ));
 sky130_fd_sc_hd__dfxtp_4 _19849_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00765_),
    .Q(\coreWBInterface.readDataBuffered[18] ));
 sky130_fd_sc_hd__dfxtp_4 _19850_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00766_),
    .Q(\coreWBInterface.readDataBuffered[19] ));
 sky130_fd_sc_hd__dfxtp_4 _19851_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00767_),
    .Q(\coreWBInterface.readDataBuffered[20] ));
 sky130_fd_sc_hd__dfxtp_4 _19852_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00768_),
    .Q(\coreWBInterface.readDataBuffered[21] ));
 sky130_fd_sc_hd__dfxtp_4 _19853_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00769_),
    .Q(\coreWBInterface.readDataBuffered[22] ));
 sky130_fd_sc_hd__dfxtp_4 _19854_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00770_),
    .Q(\coreWBInterface.readDataBuffered[23] ));
 sky130_fd_sc_hd__dfxtp_4 _19855_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00771_),
    .Q(\coreWBInterface.readDataBuffered[24] ));
 sky130_fd_sc_hd__dfxtp_4 _19856_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00772_),
    .Q(\coreWBInterface.readDataBuffered[25] ));
 sky130_fd_sc_hd__dfxtp_4 _19857_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00773_),
    .Q(\coreWBInterface.readDataBuffered[26] ));
 sky130_fd_sc_hd__dfxtp_4 _19858_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00774_),
    .Q(\coreWBInterface.readDataBuffered[27] ));
 sky130_fd_sc_hd__dfxtp_4 _19859_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00775_),
    .Q(\coreWBInterface.readDataBuffered[28] ));
 sky130_fd_sc_hd__dfxtp_4 _19860_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00776_),
    .Q(\coreWBInterface.readDataBuffered[29] ));
 sky130_fd_sc_hd__dfxtp_2 _19861_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00777_),
    .Q(\coreWBInterface.readDataBuffered[30] ));
 sky130_fd_sc_hd__dfxtp_4 _19862_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00778_),
    .Q(\coreWBInterface.readDataBuffered[31] ));
 sky130_fd_sc_hd__dfxtp_2 _19863_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_00779_),
    .Q(\coreWBInterface.state[0] ));
 sky130_fd_sc_hd__dfxtp_4 _19864_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_00780_),
    .Q(\coreWBInterface.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _19865_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_00781_),
    .Q(\core.registers[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19866_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_00782_),
    .Q(\core.registers[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19867_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_00783_),
    .Q(\core.registers[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19868_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_00784_),
    .Q(\core.registers[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19869_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_00785_),
    .Q(\core.registers[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19870_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_00786_),
    .Q(\core.registers[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19871_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00787_),
    .Q(\core.registers[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19872_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_00788_),
    .Q(\core.registers[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19873_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_00789_),
    .Q(\core.registers[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19874_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_00790_),
    .Q(\core.registers[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19875_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_00791_),
    .Q(\core.registers[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19876_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00792_),
    .Q(\core.registers[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19877_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00793_),
    .Q(\core.registers[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19878_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_00794_),
    .Q(\core.registers[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19879_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_00795_),
    .Q(\core.registers[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19880_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_00796_),
    .Q(\core.registers[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19881_ (.CLK(clknet_leaf_206_wb_clk_i),
    .D(_00797_),
    .Q(\core.registers[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19882_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_00798_),
    .Q(\core.registers[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19883_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00799_),
    .Q(\core.registers[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19884_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00800_),
    .Q(\core.registers[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19885_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_00801_),
    .Q(\core.registers[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19886_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_00802_),
    .Q(\core.registers[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19887_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_00803_),
    .Q(\core.registers[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19888_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_00804_),
    .Q(\core.registers[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19889_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_00805_),
    .Q(\core.registers[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19890_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00806_),
    .Q(\core.registers[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19891_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_00807_),
    .Q(\core.registers[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19892_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_00808_),
    .Q(\core.registers[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19893_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00809_),
    .Q(\core.registers[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19894_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_00810_),
    .Q(\core.registers[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19895_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_00811_),
    .Q(\core.registers[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19896_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_00812_),
    .Q(\core.registers[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19897_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00813_),
    .Q(\core.registers[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19898_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00814_),
    .Q(\core.registers[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19899_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00815_),
    .Q(\core.registers[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19900_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00816_),
    .Q(\core.registers[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19901_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00817_),
    .Q(\core.registers[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19902_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00818_),
    .Q(\core.registers[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19903_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00819_),
    .Q(\core.registers[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19904_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00820_),
    .Q(\core.registers[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19905_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00821_),
    .Q(\core.registers[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19906_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00822_),
    .Q(\core.registers[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19907_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00823_),
    .Q(\core.registers[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19908_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00824_),
    .Q(\core.registers[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19909_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00825_),
    .Q(\core.registers[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19910_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00826_),
    .Q(\core.registers[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19911_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00827_),
    .Q(\core.registers[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19912_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00828_),
    .Q(\core.registers[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19913_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_00829_),
    .Q(\core.registers[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19914_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00830_),
    .Q(\core.registers[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19915_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00831_),
    .Q(\core.registers[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19916_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00832_),
    .Q(\core.registers[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19917_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00833_),
    .Q(\core.registers[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19918_ (.CLK(clknet_leaf_203_wb_clk_i),
    .D(_00834_),
    .Q(\core.registers[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19919_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00835_),
    .Q(\core.registers[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19920_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00836_),
    .Q(\core.registers[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19921_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00837_),
    .Q(\core.registers[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19922_ (.CLK(clknet_leaf_211_wb_clk_i),
    .D(_00838_),
    .Q(\core.registers[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19923_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00839_),
    .Q(\core.registers[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19924_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00840_),
    .Q(\core.registers[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19925_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00841_),
    .Q(\core.registers[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19926_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00842_),
    .Q(\core.registers[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19927_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00843_),
    .Q(\core.registers[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19928_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00844_),
    .Q(\core.registers[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19929_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00845_),
    .Q(\core.registers[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _19930_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_00846_),
    .Q(\core.registers[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _19931_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00847_),
    .Q(\core.registers[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _19932_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00848_),
    .Q(\core.registers[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _19933_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00849_),
    .Q(\core.registers[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _19934_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00850_),
    .Q(\core.registers[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _19935_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00851_),
    .Q(\core.registers[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _19936_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00852_),
    .Q(\core.registers[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _19937_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_00853_),
    .Q(\core.registers[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _19938_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00854_),
    .Q(\core.registers[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _19939_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_00855_),
    .Q(\core.registers[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _19940_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00856_),
    .Q(\core.registers[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _19941_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00857_),
    .Q(\core.registers[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _19942_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_00858_),
    .Q(\core.registers[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _19943_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00859_),
    .Q(\core.registers[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _19944_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00860_),
    .Q(\core.registers[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _19945_ (.CLK(clknet_leaf_206_wb_clk_i),
    .D(_00861_),
    .Q(\core.registers[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _19946_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00862_),
    .Q(\core.registers[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _19947_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00863_),
    .Q(\core.registers[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _19948_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00864_),
    .Q(\core.registers[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _19949_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_00865_),
    .Q(\core.registers[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _19950_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00866_),
    .Q(\core.registers[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _19951_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00867_),
    .Q(\core.registers[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _19952_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00868_),
    .Q(\core.registers[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _19953_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_00869_),
    .Q(\core.registers[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _19954_ (.CLK(clknet_leaf_212_wb_clk_i),
    .D(_00870_),
    .Q(\core.registers[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _19955_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00871_),
    .Q(\core.registers[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _19956_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_00872_),
    .Q(\core.registers[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _19957_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00873_),
    .Q(\core.registers[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _19958_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00874_),
    .Q(\core.registers[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _19959_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_00875_),
    .Q(\core.registers[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _19960_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_00876_),
    .Q(\core.registers[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _19961_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00877_),
    .Q(net410));
 sky130_fd_sc_hd__dfxtp_1 _19962_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00878_),
    .Q(net421));
 sky130_fd_sc_hd__dfxtp_1 _19963_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00879_),
    .Q(net432));
 sky130_fd_sc_hd__dfxtp_1 _19964_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00880_),
    .Q(net435));
 sky130_fd_sc_hd__dfxtp_1 _19965_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00881_),
    .Q(net436));
 sky130_fd_sc_hd__dfxtp_1 _19966_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00882_),
    .Q(net437));
 sky130_fd_sc_hd__dfxtp_1 _19967_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00883_),
    .Q(net438));
 sky130_fd_sc_hd__dfxtp_1 _19968_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00884_),
    .Q(net439));
 sky130_fd_sc_hd__dfxtp_1 _19969_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00885_),
    .Q(net440));
 sky130_fd_sc_hd__dfxtp_2 _19970_ (.CLK(clknet_leaf_154_wb_clk_i),
    .D(_00886_),
    .Q(net441));
 sky130_fd_sc_hd__dfxtp_1 _19971_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_00887_),
    .Q(net411));
 sky130_fd_sc_hd__dfxtp_1 _19972_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00888_),
    .Q(net412));
 sky130_fd_sc_hd__dfxtp_1 _19973_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00889_),
    .Q(net413));
 sky130_fd_sc_hd__dfxtp_1 _19974_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_00890_),
    .Q(net414));
 sky130_fd_sc_hd__dfxtp_1 _19975_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00891_),
    .Q(net415));
 sky130_fd_sc_hd__dfxtp_1 _19976_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00892_),
    .Q(net416));
 sky130_fd_sc_hd__dfxtp_1 _19977_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00893_),
    .Q(net417));
 sky130_fd_sc_hd__dfxtp_2 _19978_ (.CLK(clknet_leaf_123_wb_clk_i),
    .D(_00894_),
    .Q(net418));
 sky130_fd_sc_hd__dfxtp_1 _19979_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00895_),
    .Q(net419));
 sky130_fd_sc_hd__dfxtp_2 _19980_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_00896_),
    .Q(net420));
 sky130_fd_sc_hd__dfxtp_1 _19981_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00897_),
    .Q(net422));
 sky130_fd_sc_hd__dfxtp_1 _19982_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00898_),
    .Q(net423));
 sky130_fd_sc_hd__dfxtp_1 _19983_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00899_),
    .Q(net424));
 sky130_fd_sc_hd__dfxtp_1 _19984_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00900_),
    .Q(net425));
 sky130_fd_sc_hd__dfxtp_1 _19985_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00901_),
    .Q(net426));
 sky130_fd_sc_hd__dfxtp_1 _19986_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00902_),
    .Q(net427));
 sky130_fd_sc_hd__dfxtp_1 _19987_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00903_),
    .Q(net428));
 sky130_fd_sc_hd__dfxtp_1 _19988_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00904_),
    .Q(net429));
 sky130_fd_sc_hd__dfxtp_1 _19989_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00905_),
    .Q(net430));
 sky130_fd_sc_hd__dfxtp_1 _19990_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_00906_),
    .Q(net431));
 sky130_fd_sc_hd__dfxtp_1 _19991_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00907_),
    .Q(net433));
 sky130_fd_sc_hd__dfxtp_1 _19992_ (.CLK(clknet_leaf_110_wb_clk_i),
    .D(_00908_),
    .Q(net434));
 sky130_fd_sc_hd__dfxtp_1 _19993_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00909_),
    .Q(net409));
 sky130_fd_sc_hd__dfxtp_1 _19994_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00910_),
    .Q(net442));
 sky130_fd_sc_hd__dfxtp_1 _19995_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00911_),
    .Q(\wbSRAMInterface.currentAddress[0] ));
 sky130_fd_sc_hd__dfxtp_1 _19996_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00912_),
    .Q(\wbSRAMInterface.currentAddress[1] ));
 sky130_fd_sc_hd__dfxtp_4 _19997_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00913_),
    .Q(\wbSRAMInterface.currentAddress[2] ));
 sky130_fd_sc_hd__dfxtp_4 _19998_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00914_),
    .Q(\wbSRAMInterface.currentAddress[3] ));
 sky130_fd_sc_hd__dfxtp_4 _19999_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00915_),
    .Q(\wbSRAMInterface.currentAddress[4] ));
 sky130_fd_sc_hd__dfxtp_4 _20000_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_00916_),
    .Q(\wbSRAMInterface.currentAddress[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20001_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00917_),
    .Q(\wbSRAMInterface.currentAddress[6] ));
 sky130_fd_sc_hd__dfxtp_4 _20002_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00918_),
    .Q(\wbSRAMInterface.currentAddress[7] ));
 sky130_fd_sc_hd__dfxtp_4 _20003_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00919_),
    .Q(\wbSRAMInterface.currentAddress[8] ));
 sky130_fd_sc_hd__dfxtp_4 _20004_ (.CLK(clknet_leaf_122_wb_clk_i),
    .D(_00920_),
    .Q(\wbSRAMInterface.currentAddress[9] ));
 sky130_fd_sc_hd__dfxtp_4 _20005_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00921_),
    .Q(\wbSRAMInterface.currentAddress[10] ));
 sky130_fd_sc_hd__dfxtp_4 _20006_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00922_),
    .Q(\wbSRAMInterface.currentAddress[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20007_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00923_),
    .Q(\wbSRAMInterface.currentAddress[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20008_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00924_),
    .Q(\wbSRAMInterface.currentAddress[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20009_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00925_),
    .Q(\wbSRAMInterface.currentAddress[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20010_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_00926_),
    .Q(\wbSRAMInterface.currentAddress[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20011_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00927_),
    .Q(\wbSRAMInterface.currentAddress[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20012_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00928_),
    .Q(\wbSRAMInterface.currentAddress[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20013_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00929_),
    .Q(\wbSRAMInterface.currentAddress[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20014_ (.CLK(clknet_leaf_113_wb_clk_i),
    .D(_00930_),
    .Q(\wbSRAMInterface.currentAddress[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20015_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00931_),
    .Q(\wbSRAMInterface.currentAddress[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20016_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00932_),
    .Q(\wbSRAMInterface.currentAddress[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20017_ (.CLK(clknet_leaf_112_wb_clk_i),
    .D(_00933_),
    .Q(\wbSRAMInterface.currentAddress[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20018_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_00934_),
    .Q(\wbSRAMInterface.currentAddress[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20019_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_00935_),
    .Q(\memoryController.last_data_enableWB ));
 sky130_fd_sc_hd__dfxtp_4 _20020_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00936_),
    .Q(\wbSRAMInterface.state[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20021_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_00937_),
    .Q(\wbSRAMInterface.state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20022_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00938_),
    .Q(\core.registers[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20023_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_00939_),
    .Q(\core.registers[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20024_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_00940_),
    .Q(\core.registers[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20025_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_00941_),
    .Q(\core.registers[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20026_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00942_),
    .Q(\core.registers[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20027_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00943_),
    .Q(\core.registers[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20028_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00944_),
    .Q(\core.registers[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20029_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00945_),
    .Q(\core.registers[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20030_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_00946_),
    .Q(\core.registers[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20031_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00947_),
    .Q(\core.registers[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20032_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_00948_),
    .Q(\core.registers[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20033_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_00949_),
    .Q(\core.registers[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20034_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00950_),
    .Q(\core.registers[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20035_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00951_),
    .Q(\core.registers[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20036_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00952_),
    .Q(\core.registers[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20037_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00953_),
    .Q(\core.registers[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20038_ (.CLK(clknet_leaf_206_wb_clk_i),
    .D(_00954_),
    .Q(\core.registers[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20039_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00955_),
    .Q(\core.registers[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20040_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00956_),
    .Q(\core.registers[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20041_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00957_),
    .Q(\core.registers[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20042_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_00958_),
    .Q(\core.registers[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20043_ (.CLK(clknet_leaf_204_wb_clk_i),
    .D(_00959_),
    .Q(\core.registers[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20044_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00960_),
    .Q(\core.registers[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20045_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00961_),
    .Q(\core.registers[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20046_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00962_),
    .Q(\core.registers[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20047_ (.CLK(clknet_leaf_212_wb_clk_i),
    .D(_00963_),
    .Q(\core.registers[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20048_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00964_),
    .Q(\core.registers[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20049_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_00965_),
    .Q(\core.registers[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20050_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_00966_),
    .Q(\core.registers[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20051_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00967_),
    .Q(\core.registers[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20052_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_00968_),
    .Q(\core.registers[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20053_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00969_),
    .Q(\core.registers[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20054_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00970_),
    .Q(\core.registers[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20055_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00971_),
    .Q(\core.registers[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20056_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00972_),
    .Q(\core.registers[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20057_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_00973_),
    .Q(\core.registers[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20058_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_00974_),
    .Q(\core.registers[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20059_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_00975_),
    .Q(\core.registers[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20060_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_00976_),
    .Q(\core.registers[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20061_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_00977_),
    .Q(\core.registers[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20062_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_00978_),
    .Q(\core.registers[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20063_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_00979_),
    .Q(\core.registers[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20064_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_00980_),
    .Q(\core.registers[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20065_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_00981_),
    .Q(\core.registers[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20066_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_00982_),
    .Q(\core.registers[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20067_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_00983_),
    .Q(\core.registers[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20068_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_00984_),
    .Q(\core.registers[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20069_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_00985_),
    .Q(\core.registers[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20070_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_00986_),
    .Q(\core.registers[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20071_ (.CLK(clknet_leaf_203_wb_clk_i),
    .D(_00987_),
    .Q(\core.registers[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20072_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_00988_),
    .Q(\core.registers[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20073_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_00989_),
    .Q(\core.registers[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20074_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_00990_),
    .Q(\core.registers[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20075_ (.CLK(clknet_leaf_202_wb_clk_i),
    .D(_00991_),
    .Q(\core.registers[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20076_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_00992_),
    .Q(\core.registers[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20077_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_00993_),
    .Q(\core.registers[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20078_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_00994_),
    .Q(\core.registers[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20079_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_00995_),
    .Q(\core.registers[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20080_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_00996_),
    .Q(\core.registers[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20081_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_00997_),
    .Q(\core.registers[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20082_ (.CLK(clknet_leaf_203_wb_clk_i),
    .D(_00998_),
    .Q(\core.registers[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20083_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_00999_),
    .Q(\core.registers[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20084_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_01000_),
    .Q(\core.registers[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20085_ (.CLK(clknet_leaf_64_wb_clk_i),
    .D(_01001_),
    .Q(\core.registers[21][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20086_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01002_),
    .Q(\core.registers[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20087_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01003_),
    .Q(\core.registers[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20088_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01004_),
    .Q(\core.registers[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20089_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01005_),
    .Q(\core.registers[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20090_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01006_),
    .Q(\core.registers[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20091_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01007_),
    .Q(\core.registers[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20092_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01008_),
    .Q(\core.registers[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20093_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01009_),
    .Q(\core.registers[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20094_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01010_),
    .Q(\core.registers[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20095_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01011_),
    .Q(\core.registers[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20096_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01012_),
    .Q(\core.registers[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20097_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01013_),
    .Q(\core.registers[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20098_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01014_),
    .Q(\core.registers[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20099_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01015_),
    .Q(\core.registers[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20100_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01016_),
    .Q(\core.registers[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20101_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01017_),
    .Q(\core.registers[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20102_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_01018_),
    .Q(\core.registers[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20103_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01019_),
    .Q(\core.registers[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20104_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01020_),
    .Q(\core.registers[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20105_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_01021_),
    .Q(\core.registers[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20106_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01022_),
    .Q(\core.registers[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20107_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_01023_),
    .Q(\core.registers[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20108_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01024_),
    .Q(\core.registers[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20109_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01025_),
    .Q(\core.registers[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20110_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01026_),
    .Q(\core.registers[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20111_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_01027_),
    .Q(\core.registers[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20112_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01028_),
    .Q(\core.registers[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20113_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01029_),
    .Q(\core.registers[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20114_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01030_),
    .Q(\core.registers[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20115_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01031_),
    .Q(\core.registers[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20116_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01032_),
    .Q(\core.registers[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20117_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01033_),
    .Q(\core.registers[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20118_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01034_),
    .Q(\core.registers[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20119_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01035_),
    .Q(\core.registers[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20120_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01036_),
    .Q(\core.registers[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20121_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01037_),
    .Q(\core.registers[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20122_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01038_),
    .Q(\core.registers[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20123_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01039_),
    .Q(\core.registers[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20124_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01040_),
    .Q(\core.registers[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20125_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01041_),
    .Q(\core.registers[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20126_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01042_),
    .Q(\core.registers[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20127_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01043_),
    .Q(\core.registers[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20128_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01044_),
    .Q(\core.registers[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20129_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01045_),
    .Q(\core.registers[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20130_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01046_),
    .Q(\core.registers[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20131_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01047_),
    .Q(\core.registers[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20132_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01048_),
    .Q(\core.registers[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20133_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01049_),
    .Q(\core.registers[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20134_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_01050_),
    .Q(\core.registers[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20135_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01051_),
    .Q(\core.registers[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20136_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01052_),
    .Q(\core.registers[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20137_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_01053_),
    .Q(\core.registers[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20138_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01054_),
    .Q(\core.registers[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20139_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_01055_),
    .Q(\core.registers[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20140_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01056_),
    .Q(\core.registers[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20141_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01057_),
    .Q(\core.registers[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20142_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01058_),
    .Q(\core.registers[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20143_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_01059_),
    .Q(\core.registers[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20144_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01060_),
    .Q(\core.registers[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20145_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01061_),
    .Q(\core.registers[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20146_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01062_),
    .Q(\core.registers[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20147_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01063_),
    .Q(\core.registers[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20148_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01064_),
    .Q(\core.registers[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20149_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01065_),
    .Q(\core.registers[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20150_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01066_),
    .Q(\core.registers[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20151_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01067_),
    .Q(\core.registers[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20152_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01068_),
    .Q(\core.registers[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20153_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01069_),
    .Q(\core.registers[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20154_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01070_),
    .Q(\core.registers[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20155_ (.CLK(clknet_leaf_60_wb_clk_i),
    .D(_01071_),
    .Q(\core.registers[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20156_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01072_),
    .Q(\core.registers[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20157_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01073_),
    .Q(\core.registers[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20158_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01074_),
    .Q(\core.registers[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20159_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01075_),
    .Q(\core.registers[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20160_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01076_),
    .Q(\core.registers[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20161_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01077_),
    .Q(\core.registers[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20162_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01078_),
    .Q(\core.registers[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20163_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01079_),
    .Q(\core.registers[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20164_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01080_),
    .Q(\core.registers[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20165_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01081_),
    .Q(\core.registers[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20166_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_01082_),
    .Q(\core.registers[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20167_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01083_),
    .Q(\core.registers[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20168_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01084_),
    .Q(\core.registers[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20169_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_01085_),
    .Q(\core.registers[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20170_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01086_),
    .Q(\core.registers[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20171_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_01087_),
    .Q(\core.registers[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20172_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01088_),
    .Q(\core.registers[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20173_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_01089_),
    .Q(\core.registers[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20174_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01090_),
    .Q(\core.registers[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20175_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_01091_),
    .Q(\core.registers[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20176_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01092_),
    .Q(\core.registers[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20177_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01093_),
    .Q(\core.registers[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20178_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01094_),
    .Q(\core.registers[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20179_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_01095_),
    .Q(\core.registers[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20180_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_01096_),
    .Q(\core.registers[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20181_ (.CLK(clknet_leaf_73_wb_clk_i),
    .D(_01097_),
    .Q(\core.registers[13][31] ));
 sky130_fd_sc_hd__dfxtp_4 _20182_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01098_),
    .Q(\core.management_interruptEnable ));
 sky130_fd_sc_hd__dfxtp_1 _20183_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01099_),
    .Q(\coreManagement.control[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20184_ (.CLK(clknet_leaf_134_wb_clk_i),
    .D(_01100_),
    .Q(\core.management_run ));
 sky130_fd_sc_hd__dfxtp_1 _20185_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01101_),
    .Q(\jtag.dataIDRegister.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20186_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01102_),
    .Q(\jtag.dataIDRegister.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20187_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01103_),
    .Q(\jtag.dataIDRegister.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20188_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01104_),
    .Q(\jtag.dataIDRegister.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20189_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01105_),
    .Q(\jtag.dataIDRegister.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20190_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01106_),
    .Q(\jtag.dataIDRegister.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20191_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01107_),
    .Q(\jtag.dataIDRegister.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20192_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01108_),
    .Q(\jtag.dataIDRegister.data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20193_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01109_),
    .Q(\jtag.dataIDRegister.data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20194_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01110_),
    .Q(\jtag.dataIDRegister.data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20195_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01111_),
    .Q(\jtag.dataIDRegister.data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20196_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01112_),
    .Q(\jtag.dataIDRegister.data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20197_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01113_),
    .Q(\jtag.dataIDRegister.data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20198_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01114_),
    .Q(\jtag.dataIDRegister.data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20199_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01115_),
    .Q(\jtag.dataIDRegister.data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20200_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01116_),
    .Q(\jtag.dataIDRegister.data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20201_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01117_),
    .Q(\jtag.dataIDRegister.data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20202_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_01118_),
    .Q(\jtag.dataIDRegister.data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20203_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_01119_),
    .Q(\jtag.dataIDRegister.data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20204_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_01120_),
    .Q(\jtag.dataIDRegister.data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20205_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_01121_),
    .Q(\jtag.dataIDRegister.data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20206_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01122_),
    .Q(\jtag.dataIDRegister.data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20207_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01123_),
    .Q(\jtag.dataIDRegister.data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20208_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01124_),
    .Q(\jtag.dataIDRegister.data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20209_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01125_),
    .Q(\jtag.dataIDRegister.data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20210_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01126_),
    .Q(\jtag.dataIDRegister.data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20211_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01127_),
    .Q(\jtag.dataIDRegister.data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20212_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01128_),
    .Q(\jtag.dataIDRegister.data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20213_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01129_),
    .Q(\jtag.dataIDRegister.data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20214_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01130_),
    .Q(\jtag.dataIDRegister.data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20215_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01131_),
    .Q(\jtag.dataIDRegister.data[30] ));
 sky130_fd_sc_hd__dfxtp_4 _20216_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01132_),
    .Q(\jtag.dataIDRegister.data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20217_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01133_),
    .Q(\jtag.dataBypassRegister.data ));
 sky130_fd_sc_hd__dfxtp_1 _20218_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01134_),
    .Q(\jtag.dataBSRRegister.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20219_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_01135_),
    .Q(\jtag.dataBSRRegister.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20220_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_01136_),
    .Q(\jtag.dataBSRRegister.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20221_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_01137_),
    .Q(\jtag.dataBSRRegister.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20222_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01138_),
    .Q(\jtag.dataBSRRegister.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20223_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_01139_),
    .Q(\jtag.dataBSRRegister.data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20224_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_01140_),
    .Q(\jtag.dataBSRRegister.data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20225_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_01141_),
    .Q(\jtag.dataBSRRegister.data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20226_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_01142_),
    .Q(\jtag.dataBSRRegister.data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20227_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01143_),
    .Q(\jtag.dataBSRRegister.data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20228_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01144_),
    .Q(\jtag.dataBSRRegister.data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20229_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01145_),
    .Q(\jtag.dataBSRRegister.data[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20230_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01146_),
    .Q(\jtag.dataBSRRegister.data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20231_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_01147_),
    .Q(\jtag.dataBSRRegister.data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20232_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01148_),
    .Q(\jtag.dataBSRRegister.data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20233_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01149_),
    .Q(\jtag.dataBSRRegister.data[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20234_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_01150_),
    .Q(\jtag.dataBSRRegister.data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20235_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01151_),
    .Q(\jtag.dataBSRRegister.data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20236_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01152_),
    .Q(\jtag.dataBSRRegister.data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20237_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01153_),
    .Q(\jtag.dataBSRRegister.data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20238_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_01154_),
    .Q(\jtag.dataBSRRegister.data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20239_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01155_),
    .Q(\jtag.dataBSRRegister.data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20240_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01156_),
    .Q(\jtag.dataBSRRegister.data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20241_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01157_),
    .Q(\jtag.dataBSRRegister.data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20242_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01158_),
    .Q(\jtag.dataBSRRegister.data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20243_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01159_),
    .Q(\jtag.dataBSRRegister.data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20244_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01160_),
    .Q(\jtag.dataBSRRegister.data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20245_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01161_),
    .Q(\jtag.dataBSRRegister.data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20246_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01162_),
    .Q(\jtag.dataBSRRegister.data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20247_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01163_),
    .Q(\jtag.dataBSRRegister.data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20248_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01164_),
    .Q(\jtag.dataBSRRegister.data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20249_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_01165_),
    .Q(\jtag.dataBSRRegister.data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20250_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01166_),
    .Q(\jtag.instructionRegister.data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20251_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01167_),
    .Q(\jtag.instructionRegister.data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20252_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01168_),
    .Q(\jtag.instructionRegister.data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20253_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01169_),
    .Q(\jtag.instructionRegister.data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20254_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01170_),
    .Q(\jtag.instructionRegister.data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20255_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01171_),
    .Q(\jtag.tckRisingEdge ));
 sky130_fd_sc_hd__dfxtp_1 _20256_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01172_),
    .Q(\jtag.tckState ));
 sky130_fd_sc_hd__dfxtp_4 _20257_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01173_),
    .Q(net445));
 sky130_fd_sc_hd__dfxtp_4 _20258_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01174_),
    .Q(net446));
 sky130_fd_sc_hd__dfxtp_4 _20259_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_01175_),
    .Q(net447));
 sky130_fd_sc_hd__dfxtp_4 _20260_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01176_),
    .Q(net448));
 sky130_fd_sc_hd__dfxtp_4 _20261_ (.CLK(clknet_leaf_183_wb_clk_i),
    .D(_01177_),
    .Q(net449));
 sky130_fd_sc_hd__dfxtp_1 _20262_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_01178_),
    .Q(\jtag.state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20263_ (.CLK(clknet_leaf_186_wb_clk_i),
    .D(_01179_),
    .Q(\jtag.state[1] ));
 sky130_fd_sc_hd__dfxtp_4 _20264_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_01180_),
    .Q(\jtag.state[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20265_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_01181_),
    .Q(\jtag.state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20266_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01182_),
    .Q(\jtag.managementReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20267_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01183_),
    .Q(\jtag.managementReadData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20268_ (.CLK(clknet_leaf_124_wb_clk_i),
    .D(_01184_),
    .Q(\jtag.managementReadData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20269_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01185_),
    .Q(\jtag.managementReadData[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20270_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01186_),
    .Q(\jtag.managementReadData[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20271_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_01187_),
    .Q(\jtag.managementReadData[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20272_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01188_),
    .Q(\jtag.managementReadData[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20273_ (.CLK(clknet_leaf_86_wb_clk_i),
    .D(_01189_),
    .Q(\jtag.managementReadData[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20274_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_01190_),
    .Q(\jtag.managementReadData[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20275_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01191_),
    .Q(\jtag.managementReadData[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20276_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01192_),
    .Q(\jtag.managementReadData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20277_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01193_),
    .Q(\jtag.managementReadData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20278_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01194_),
    .Q(\jtag.managementReadData[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20279_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01195_),
    .Q(\jtag.managementReadData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20280_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01196_),
    .Q(\jtag.managementReadData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20281_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01197_),
    .Q(\jtag.managementReadData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20282_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_01198_),
    .Q(\jtag.managementReadData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20283_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01199_),
    .Q(\jtag.managementReadData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20284_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01200_),
    .Q(\jtag.managementReadData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20285_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01201_),
    .Q(\jtag.managementReadData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20286_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01202_),
    .Q(\jtag.managementReadData[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20287_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01203_),
    .Q(\jtag.managementReadData[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20288_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01204_),
    .Q(\jtag.managementReadData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20289_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01205_),
    .Q(\jtag.managementReadData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20290_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01206_),
    .Q(\jtag.managementReadData[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20291_ (.CLK(clknet_leaf_179_wb_clk_i),
    .D(_01207_),
    .Q(\jtag.managementReadData[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20292_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01208_),
    .Q(\jtag.managementReadData[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20293_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01209_),
    .Q(\jtag.managementReadData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20294_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01210_),
    .Q(\jtag.managementReadData[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20295_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01211_),
    .Q(\jtag.managementReadData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20296_ (.CLK(clknet_leaf_180_wb_clk_i),
    .D(_01212_),
    .Q(\jtag.managementReadData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20297_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_01213_),
    .Q(\jtag.managementReadData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20298_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_01214_),
    .Q(\jtag.managementState[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20299_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_01215_),
    .Q(\jtag.managementState[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20300_ (.CLK(clknet_leaf_181_wb_clk_i),
    .D(_01216_),
    .Q(\jtag.managementState[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20301_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01217_),
    .Q(\core.registers[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20302_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01218_),
    .Q(\core.registers[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20303_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01219_),
    .Q(\core.registers[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20304_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01220_),
    .Q(\core.registers[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20305_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_01221_),
    .Q(\core.registers[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20306_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01222_),
    .Q(\core.registers[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20307_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_01223_),
    .Q(\core.registers[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20308_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01224_),
    .Q(\core.registers[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20309_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01225_),
    .Q(\core.registers[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20310_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01226_),
    .Q(\core.registers[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20311_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01227_),
    .Q(\core.registers[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20312_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01228_),
    .Q(\core.registers[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20313_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01229_),
    .Q(\core.registers[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20314_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01230_),
    .Q(\core.registers[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20315_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_01231_),
    .Q(\core.registers[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20316_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01232_),
    .Q(\core.registers[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20317_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_01233_),
    .Q(\core.registers[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20318_ (.CLK(clknet_leaf_204_wb_clk_i),
    .D(_01234_),
    .Q(\core.registers[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20319_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_01235_),
    .Q(\core.registers[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20320_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01236_),
    .Q(\core.registers[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20321_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01237_),
    .Q(\core.registers[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20322_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_01238_),
    .Q(\core.registers[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20323_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01239_),
    .Q(\core.registers[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20324_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_01240_),
    .Q(\core.registers[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20325_ (.CLK(clknet_leaf_218_wb_clk_i),
    .D(_01241_),
    .Q(\core.registers[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20326_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_01242_),
    .Q(\core.registers[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20327_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01243_),
    .Q(\core.registers[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20328_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01244_),
    .Q(\core.registers[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20329_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01245_),
    .Q(\core.registers[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20330_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01246_),
    .Q(\core.registers[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20331_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01247_),
    .Q(\core.registers[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20332_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01248_),
    .Q(\core.registers[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20333_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01249_),
    .Q(\core.registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20334_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01250_),
    .Q(\core.registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20335_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01251_),
    .Q(\core.registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20336_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01252_),
    .Q(\core.registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20337_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01253_),
    .Q(\core.registers[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20338_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01254_),
    .Q(\core.registers[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20339_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_01255_),
    .Q(\core.registers[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20340_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01256_),
    .Q(\core.registers[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20341_ (.CLK(clknet_leaf_71_wb_clk_i),
    .D(_01257_),
    .Q(\core.registers[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20342_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01258_),
    .Q(\core.registers[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20343_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01259_),
    .Q(\core.registers[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20344_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01260_),
    .Q(\core.registers[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20345_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01261_),
    .Q(\core.registers[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20346_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01262_),
    .Q(\core.registers[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20347_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01263_),
    .Q(\core.registers[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20348_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_01264_),
    .Q(\core.registers[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20349_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01265_),
    .Q(\core.registers[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20350_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01266_),
    .Q(\core.registers[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20351_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01267_),
    .Q(\core.registers[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20352_ (.CLK(clknet_leaf_210_wb_clk_i),
    .D(_01268_),
    .Q(\core.registers[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20353_ (.CLK(clknet_leaf_197_wb_clk_i),
    .D(_01269_),
    .Q(\core.registers[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20354_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01270_),
    .Q(\core.registers[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20355_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01271_),
    .Q(\core.registers[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20356_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01272_),
    .Q(\core.registers[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20357_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01273_),
    .Q(\core.registers[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20358_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_01274_),
    .Q(\core.registers[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20359_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01275_),
    .Q(\core.registers[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20360_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01276_),
    .Q(\core.registers[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20361_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01277_),
    .Q(\core.registers[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20362_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01278_),
    .Q(\core.registers[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20363_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01279_),
    .Q(\core.registers[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20364_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01280_),
    .Q(\core.registers[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20365_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01281_),
    .Q(\core.registers[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20366_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01282_),
    .Q(\core.registers[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20367_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01283_),
    .Q(\core.registers[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20368_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01284_),
    .Q(\core.registers[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20369_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_01285_),
    .Q(\core.registers[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20370_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01286_),
    .Q(\core.registers[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20371_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_01287_),
    .Q(\core.registers[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20372_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01288_),
    .Q(\core.registers[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20373_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01289_),
    .Q(\core.registers[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20374_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01290_),
    .Q(\core.registers[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20375_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01291_),
    .Q(\core.registers[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20376_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01292_),
    .Q(\core.registers[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20377_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_01293_),
    .Q(\core.registers[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20378_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01294_),
    .Q(\core.registers[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20379_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_01295_),
    .Q(\core.registers[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20380_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01296_),
    .Q(\core.registers[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20381_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_01297_),
    .Q(\core.registers[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20382_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_01298_),
    .Q(\core.registers[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20383_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01299_),
    .Q(\core.registers[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20384_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01300_),
    .Q(\core.registers[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20385_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01301_),
    .Q(\core.registers[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20386_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_01302_),
    .Q(\core.registers[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20387_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_01303_),
    .Q(\core.registers[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20388_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01304_),
    .Q(\core.registers[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20389_ (.CLK(clknet_leaf_218_wb_clk_i),
    .D(_01305_),
    .Q(\core.registers[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20390_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01306_),
    .Q(\core.registers[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20391_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01307_),
    .Q(\core.registers[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20392_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_01308_),
    .Q(\core.registers[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20393_ (.CLK(clknet_leaf_204_wb_clk_i),
    .D(_01309_),
    .Q(\core.registers[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20394_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01310_),
    .Q(\core.registers[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20395_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01311_),
    .Q(\core.registers[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20396_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01312_),
    .Q(\core.registers[10][31] ));
 sky130_fd_sc_hd__dfxtp_4 _20397_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01313_),
    .Q(\core.registers[0][0] ));
 sky130_fd_sc_hd__dfxtp_4 _20398_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01314_),
    .Q(\core.registers[0][1] ));
 sky130_fd_sc_hd__dfxtp_4 _20399_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01315_),
    .Q(\core.registers[0][2] ));
 sky130_fd_sc_hd__dfxtp_4 _20400_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01316_),
    .Q(\core.registers[0][3] ));
 sky130_fd_sc_hd__dfxtp_2 _20401_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01317_),
    .Q(\core.registers[0][4] ));
 sky130_fd_sc_hd__dfxtp_4 _20402_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01318_),
    .Q(\core.registers[0][5] ));
 sky130_fd_sc_hd__dfxtp_4 _20403_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01319_),
    .Q(\core.registers[0][6] ));
 sky130_fd_sc_hd__dfxtp_4 _20404_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01320_),
    .Q(\core.registers[0][7] ));
 sky130_fd_sc_hd__dfxtp_2 _20405_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01321_),
    .Q(\core.registers[0][8] ));
 sky130_fd_sc_hd__dfxtp_2 _20406_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01322_),
    .Q(\core.registers[0][9] ));
 sky130_fd_sc_hd__dfxtp_4 _20407_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01323_),
    .Q(\core.registers[0][10] ));
 sky130_fd_sc_hd__dfxtp_4 _20408_ (.CLK(clknet_4_3__leaf_wb_clk_i),
    .D(_01324_),
    .Q(\core.registers[0][11] ));
 sky130_fd_sc_hd__dfxtp_4 _20409_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01325_),
    .Q(\core.registers[0][12] ));
 sky130_fd_sc_hd__dfxtp_2 _20410_ (.CLK(clknet_leaf_84_wb_clk_i),
    .D(_01326_),
    .Q(\core.registers[0][13] ));
 sky130_fd_sc_hd__dfxtp_4 _20411_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01327_),
    .Q(\core.registers[0][14] ));
 sky130_fd_sc_hd__dfxtp_4 _20412_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_01328_),
    .Q(\core.registers[0][15] ));
 sky130_fd_sc_hd__dfxtp_4 _20413_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_01329_),
    .Q(\core.registers[0][16] ));
 sky130_fd_sc_hd__dfxtp_2 _20414_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_01330_),
    .Q(\core.registers[0][17] ));
 sky130_fd_sc_hd__dfxtp_4 _20415_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01331_),
    .Q(\core.registers[0][18] ));
 sky130_fd_sc_hd__dfxtp_4 _20416_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01332_),
    .Q(\core.registers[0][19] ));
 sky130_fd_sc_hd__dfxtp_2 _20417_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_01333_),
    .Q(\core.registers[0][20] ));
 sky130_fd_sc_hd__dfxtp_2 _20418_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_01334_),
    .Q(\core.registers[0][21] ));
 sky130_fd_sc_hd__dfxtp_4 _20419_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01335_),
    .Q(\core.registers[0][22] ));
 sky130_fd_sc_hd__dfxtp_4 _20420_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_01336_),
    .Q(\core.registers[0][23] ));
 sky130_fd_sc_hd__dfxtp_2 _20421_ (.CLK(clknet_leaf_182_wb_clk_i),
    .D(_01337_),
    .Q(\core.registers[0][24] ));
 sky130_fd_sc_hd__dfxtp_4 _20422_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01338_),
    .Q(\core.registers[0][25] ));
 sky130_fd_sc_hd__dfxtp_4 _20423_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01339_),
    .Q(\core.registers[0][26] ));
 sky130_fd_sc_hd__dfxtp_2 _20424_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01340_),
    .Q(\core.registers[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20425_ (.CLK(clknet_leaf_185_wb_clk_i),
    .D(_01341_),
    .Q(\core.registers[0][28] ));
 sky130_fd_sc_hd__dfxtp_4 _20426_ (.CLK(clknet_leaf_92_wb_clk_i),
    .D(_01342_),
    .Q(\core.registers[0][29] ));
 sky130_fd_sc_hd__dfxtp_4 _20427_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01343_),
    .Q(\core.registers[0][30] ));
 sky130_fd_sc_hd__dfxtp_4 _20428_ (.CLK(clknet_leaf_95_wb_clk_i),
    .D(_01344_),
    .Q(\core.registers[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20429_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01345_),
    .Q(\core.registers[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20430_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01346_),
    .Q(\core.registers[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20431_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01347_),
    .Q(\core.registers[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20432_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01348_),
    .Q(\core.registers[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20433_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_01349_),
    .Q(\core.registers[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20434_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01350_),
    .Q(\core.registers[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20435_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_01351_),
    .Q(\core.registers[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20436_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01352_),
    .Q(\core.registers[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20437_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01353_),
    .Q(\core.registers[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20438_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_01354_),
    .Q(\core.registers[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20439_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01355_),
    .Q(\core.registers[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20440_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01356_),
    .Q(\core.registers[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20441_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_01357_),
    .Q(\core.registers[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20442_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01358_),
    .Q(\core.registers[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20443_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01359_),
    .Q(\core.registers[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20444_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01360_),
    .Q(\core.registers[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20445_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_01361_),
    .Q(\core.registers[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20446_ (.CLK(clknet_leaf_203_wb_clk_i),
    .D(_01362_),
    .Q(\core.registers[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20447_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01363_),
    .Q(\core.registers[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20448_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01364_),
    .Q(\core.registers[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20449_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01365_),
    .Q(\core.registers[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20450_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_01366_),
    .Q(\core.registers[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20451_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_01367_),
    .Q(\core.registers[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20452_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01368_),
    .Q(\core.registers[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20453_ (.CLK(clknet_leaf_218_wb_clk_i),
    .D(_01369_),
    .Q(\core.registers[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20454_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01370_),
    .Q(\core.registers[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20455_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01371_),
    .Q(\core.registers[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20456_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_01372_),
    .Q(\core.registers[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20457_ (.CLK(clknet_leaf_204_wb_clk_i),
    .D(_01373_),
    .Q(\core.registers[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20458_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01374_),
    .Q(\core.registers[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20459_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01375_),
    .Q(\core.registers[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20460_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01376_),
    .Q(\core.registers[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20461_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01377_),
    .Q(\core.registers[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20462_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01378_),
    .Q(\core.registers[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20463_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_01379_),
    .Q(\core.registers[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20464_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01380_),
    .Q(\core.registers[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20465_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_01381_),
    .Q(\core.registers[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20466_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01382_),
    .Q(\core.registers[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20467_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_01383_),
    .Q(\core.registers[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20468_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_01384_),
    .Q(\core.registers[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20469_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01385_),
    .Q(\core.registers[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20470_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01386_),
    .Q(\core.registers[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20471_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_01387_),
    .Q(\core.registers[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20472_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_01388_),
    .Q(\core.registers[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20473_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01389_),
    .Q(\core.registers[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20474_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01390_),
    .Q(\core.registers[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20475_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01391_),
    .Q(\core.registers[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20476_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01392_),
    .Q(\core.registers[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20477_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_01393_),
    .Q(\core.registers[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20478_ (.CLK(clknet_leaf_204_wb_clk_i),
    .D(_01394_),
    .Q(\core.registers[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20479_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_01395_),
    .Q(\core.registers[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20480_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_01396_),
    .Q(\core.registers[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20481_ (.CLK(clknet_leaf_217_wb_clk_i),
    .D(_01397_),
    .Q(\core.registers[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20482_ (.CLK(clknet_leaf_215_wb_clk_i),
    .D(_01398_),
    .Q(\core.registers[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20483_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01399_),
    .Q(\core.registers[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20484_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_01400_),
    .Q(\core.registers[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20485_ (.CLK(clknet_leaf_218_wb_clk_i),
    .D(_01401_),
    .Q(\core.registers[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20486_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_01402_),
    .Q(\core.registers[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20487_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01403_),
    .Q(\core.registers[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20488_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01404_),
    .Q(\core.registers[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20489_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01405_),
    .Q(\core.registers[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20490_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01406_),
    .Q(\core.registers[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20491_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_01407_),
    .Q(\core.registers[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20492_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01408_),
    .Q(\core.registers[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20493_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01409_),
    .Q(\core.registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20494_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01410_),
    .Q(\core.registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20495_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01411_),
    .Q(\core.registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20496_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01412_),
    .Q(\core.registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20497_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01413_),
    .Q(\core.registers[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20498_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01414_),
    .Q(\core.registers[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20499_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01415_),
    .Q(\core.registers[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20500_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01416_),
    .Q(\core.registers[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20501_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01417_),
    .Q(\core.registers[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20502_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01418_),
    .Q(\core.registers[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20503_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01419_),
    .Q(\core.registers[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20504_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01420_),
    .Q(\core.registers[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20505_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_01421_),
    .Q(\core.registers[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20506_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01422_),
    .Q(\core.registers[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20507_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01423_),
    .Q(\core.registers[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20508_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01424_),
    .Q(\core.registers[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20509_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01425_),
    .Q(\core.registers[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20510_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01426_),
    .Q(\core.registers[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20511_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01427_),
    .Q(\core.registers[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20512_ (.CLK(clknet_leaf_210_wb_clk_i),
    .D(_01428_),
    .Q(\core.registers[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20513_ (.CLK(clknet_leaf_208_wb_clk_i),
    .D(_01429_),
    .Q(\core.registers[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20514_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01430_),
    .Q(\core.registers[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20515_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01431_),
    .Q(\core.registers[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20516_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_01432_),
    .Q(\core.registers[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20517_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01433_),
    .Q(\core.registers[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20518_ (.CLK(clknet_leaf_211_wb_clk_i),
    .D(_01434_),
    .Q(\core.registers[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20519_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01435_),
    .Q(\core.registers[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20520_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01436_),
    .Q(\core.registers[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20521_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01437_),
    .Q(\core.registers[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20522_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01438_),
    .Q(\core.registers[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20523_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01439_),
    .Q(\core.registers[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20524_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01440_),
    .Q(\core.registers[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20525_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01441_),
    .Q(\core.registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20526_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01442_),
    .Q(\core.registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20527_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01443_),
    .Q(\core.registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20528_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01444_),
    .Q(\core.registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20529_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01445_),
    .Q(\core.registers[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20530_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01446_),
    .Q(\core.registers[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20531_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01447_),
    .Q(\core.registers[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20532_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01448_),
    .Q(\core.registers[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20533_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01449_),
    .Q(\core.registers[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20534_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01450_),
    .Q(\core.registers[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20535_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01451_),
    .Q(\core.registers[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20536_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01452_),
    .Q(\core.registers[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20537_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_01453_),
    .Q(\core.registers[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20538_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01454_),
    .Q(\core.registers[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20539_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_01455_),
    .Q(\core.registers[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20540_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01456_),
    .Q(\core.registers[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20541_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01457_),
    .Q(\core.registers[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20542_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01458_),
    .Q(\core.registers[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20543_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01459_),
    .Q(\core.registers[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20544_ (.CLK(clknet_leaf_210_wb_clk_i),
    .D(_01460_),
    .Q(\core.registers[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20545_ (.CLK(clknet_leaf_208_wb_clk_i),
    .D(_01461_),
    .Q(\core.registers[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20546_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01462_),
    .Q(\core.registers[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20547_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01463_),
    .Q(\core.registers[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20548_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_01464_),
    .Q(\core.registers[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20549_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01465_),
    .Q(\core.registers[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20550_ (.CLK(clknet_leaf_211_wb_clk_i),
    .D(_01466_),
    .Q(\core.registers[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20551_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01467_),
    .Q(\core.registers[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20552_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01468_),
    .Q(\core.registers[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20553_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01469_),
    .Q(\core.registers[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20554_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01470_),
    .Q(\core.registers[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20555_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01471_),
    .Q(\core.registers[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20556_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01472_),
    .Q(\core.registers[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20557_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_01473_),
    .Q(\core.registers[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20558_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01474_),
    .Q(\core.registers[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20559_ (.CLK(clknet_leaf_58_wb_clk_i),
    .D(_01475_),
    .Q(\core.registers[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20560_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01476_),
    .Q(\core.registers[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20561_ (.CLK(clknet_leaf_75_wb_clk_i),
    .D(_01477_),
    .Q(\core.registers[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20562_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01478_),
    .Q(\core.registers[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20563_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(_01479_),
    .Q(\core.registers[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20564_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01480_),
    .Q(\core.registers[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20565_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_01481_),
    .Q(\core.registers[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20566_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01482_),
    .Q(\core.registers[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20567_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01483_),
    .Q(\core.registers[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20568_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_01484_),
    .Q(\core.registers[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20569_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01485_),
    .Q(\core.registers[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20570_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_01486_),
    .Q(\core.registers[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20571_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01487_),
    .Q(\core.registers[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20572_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01488_),
    .Q(\core.registers[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20573_ (.CLK(clknet_leaf_214_wb_clk_i),
    .D(_01489_),
    .Q(\core.registers[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20574_ (.CLK(clknet_leaf_196_wb_clk_i),
    .D(_01490_),
    .Q(\core.registers[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20575_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01491_),
    .Q(\core.registers[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20576_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01492_),
    .Q(\core.registers[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20577_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_01493_),
    .Q(\core.registers[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20578_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_01494_),
    .Q(\core.registers[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20579_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_01495_),
    .Q(\core.registers[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20580_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_01496_),
    .Q(\core.registers[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20581_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01497_),
    .Q(\core.registers[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20582_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_01498_),
    .Q(\core.registers[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20583_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_01499_),
    .Q(\core.registers[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20584_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01500_),
    .Q(\core.registers[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20585_ (.CLK(clknet_leaf_208_wb_clk_i),
    .D(_01501_),
    .Q(\core.registers[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20586_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_01502_),
    .Q(\core.registers[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20587_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01503_),
    .Q(\core.registers[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20588_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01504_),
    .Q(\core.registers[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20589_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01505_),
    .Q(\core.registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20590_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01506_),
    .Q(\core.registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20591_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01507_),
    .Q(\core.registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20592_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01508_),
    .Q(\core.registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20593_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01509_),
    .Q(\core.registers[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20594_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01510_),
    .Q(\core.registers[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20595_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01511_),
    .Q(\core.registers[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20596_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01512_),
    .Q(\core.registers[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20597_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01513_),
    .Q(\core.registers[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20598_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01514_),
    .Q(\core.registers[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20599_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01515_),
    .Q(\core.registers[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20600_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01516_),
    .Q(\core.registers[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20601_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01517_),
    .Q(\core.registers[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20602_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01518_),
    .Q(\core.registers[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20603_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01519_),
    .Q(\core.registers[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20604_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01520_),
    .Q(\core.registers[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20605_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01521_),
    .Q(\core.registers[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20606_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01522_),
    .Q(\core.registers[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20607_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01523_),
    .Q(\core.registers[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20608_ (.CLK(clknet_leaf_210_wb_clk_i),
    .D(_01524_),
    .Q(\core.registers[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20609_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01525_),
    .Q(\core.registers[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20610_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01526_),
    .Q(\core.registers[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20611_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01527_),
    .Q(\core.registers[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20612_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_01528_),
    .Q(\core.registers[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20613_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01529_),
    .Q(\core.registers[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20614_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_01530_),
    .Q(\core.registers[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20615_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01531_),
    .Q(\core.registers[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20616_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01532_),
    .Q(\core.registers[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20617_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01533_),
    .Q(\core.registers[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20618_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01534_),
    .Q(\core.registers[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20619_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01535_),
    .Q(\core.registers[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20620_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01536_),
    .Q(\core.registers[5][31] ));
 sky130_fd_sc_hd__dfxtp_4 _20621_ (.CLK(clknet_leaf_126_wb_clk_i),
    .D(_01537_),
    .Q(\wbSRAMInterface.currentByteSelect[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20622_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_01538_),
    .Q(\wbSRAMInterface.currentByteSelect[1] ));
 sky130_fd_sc_hd__dfxtp_4 _20623_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_01539_),
    .Q(\wbSRAMInterface.currentByteSelect[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20624_ (.CLK(clknet_leaf_125_wb_clk_i),
    .D(_01540_),
    .Q(\wbSRAMInterface.currentByteSelect[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20625_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01541_),
    .Q(\core.registers[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20626_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01542_),
    .Q(\core.registers[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20627_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01543_),
    .Q(\core.registers[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20628_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01544_),
    .Q(\core.registers[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20629_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01545_),
    .Q(\core.registers[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20630_ (.CLK(clknet_leaf_65_wb_clk_i),
    .D(_01546_),
    .Q(\core.registers[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20631_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01547_),
    .Q(\core.registers[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20632_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01548_),
    .Q(\core.registers[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20633_ (.CLK(clknet_leaf_72_wb_clk_i),
    .D(_01549_),
    .Q(\core.registers[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20634_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01550_),
    .Q(\core.registers[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20635_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_01551_),
    .Q(\core.registers[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20636_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01552_),
    .Q(\core.registers[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20637_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01553_),
    .Q(\core.registers[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20638_ (.CLK(clknet_leaf_76_wb_clk_i),
    .D(_01554_),
    .Q(\core.registers[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20639_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01555_),
    .Q(\core.registers[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20640_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01556_),
    .Q(\core.registers[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20641_ (.CLK(clknet_leaf_205_wb_clk_i),
    .D(_01557_),
    .Q(\core.registers[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20642_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01558_),
    .Q(\core.registers[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20643_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01559_),
    .Q(\core.registers[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20644_ (.CLK(clknet_leaf_210_wb_clk_i),
    .D(_01560_),
    .Q(\core.registers[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20645_ (.CLK(clknet_leaf_204_wb_clk_i),
    .D(_01561_),
    .Q(\core.registers[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20646_ (.CLK(clknet_leaf_201_wb_clk_i),
    .D(_01562_),
    .Q(\core.registers[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20647_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_01563_),
    .Q(\core.registers[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20648_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_01564_),
    .Q(\core.registers[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20649_ (.CLK(clknet_leaf_198_wb_clk_i),
    .D(_01565_),
    .Q(\core.registers[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20650_ (.CLK(clknet_leaf_211_wb_clk_i),
    .D(_01566_),
    .Q(\core.registers[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20651_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01567_),
    .Q(\core.registers[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20652_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01568_),
    .Q(\core.registers[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20653_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01569_),
    .Q(\core.registers[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20654_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01570_),
    .Q(\core.registers[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20655_ (.CLK(clknet_leaf_62_wb_clk_i),
    .D(_01571_),
    .Q(\core.registers[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20656_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01572_),
    .Q(\core.registers[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20657_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_01573_),
    .Q(\core.registers[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20658_ (.CLK(clknet_leaf_69_wb_clk_i),
    .D(_01574_),
    .Q(\core.registers[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20659_ (.CLK(clknet_leaf_68_wb_clk_i),
    .D(_01575_),
    .Q(\core.registers[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20660_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_01576_),
    .Q(\core.registers[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20661_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01577_),
    .Q(\core.registers[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20662_ (.CLK(clknet_leaf_66_wb_clk_i),
    .D(_01578_),
    .Q(\core.registers[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20663_ (.CLK(clknet_leaf_93_wb_clk_i),
    .D(_01579_),
    .Q(\core.registers[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20664_ (.CLK(clknet_leaf_63_wb_clk_i),
    .D(_01580_),
    .Q(\core.registers[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20665_ (.CLK(clknet_leaf_70_wb_clk_i),
    .D(_01581_),
    .Q(\core.registers[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20666_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_01582_),
    .Q(\core.registers[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20667_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_01583_),
    .Q(\core.registers[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20668_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_01584_),
    .Q(\core.registers[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20669_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_01585_),
    .Q(\core.registers[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20670_ (.CLK(clknet_leaf_77_wb_clk_i),
    .D(_01586_),
    .Q(\core.registers[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20671_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_01587_),
    .Q(\core.registers[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20672_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_01588_),
    .Q(\core.registers[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20673_ (.CLK(clknet_leaf_206_wb_clk_i),
    .D(_01589_),
    .Q(\core.registers[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20674_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01590_),
    .Q(\core.registers[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20675_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_01591_),
    .Q(\core.registers[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20676_ (.CLK(clknet_leaf_210_wb_clk_i),
    .D(_01592_),
    .Q(\core.registers[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20677_ (.CLK(clknet_leaf_207_wb_clk_i),
    .D(_01593_),
    .Q(\core.registers[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20678_ (.CLK(clknet_leaf_200_wb_clk_i),
    .D(_01594_),
    .Q(\core.registers[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20679_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_01595_),
    .Q(\core.registers[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20680_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01596_),
    .Q(\core.registers[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20681_ (.CLK(clknet_leaf_199_wb_clk_i),
    .D(_01597_),
    .Q(\core.registers[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20682_ (.CLK(clknet_leaf_211_wb_clk_i),
    .D(_01598_),
    .Q(\core.registers[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20683_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_01599_),
    .Q(\core.registers[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20684_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01600_),
    .Q(\core.registers[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20685_ (.CLK(clknet_leaf_184_wb_clk_i),
    .D(_01601_),
    .Q(\core.registers[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20686_ (.CLK(clknet_leaf_67_wb_clk_i),
    .D(_01602_),
    .Q(\core.registers[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20687_ (.CLK(clknet_leaf_61_wb_clk_i),
    .D(_01603_),
    .Q(\core.registers[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20688_ (.CLK(clknet_leaf_94_wb_clk_i),
    .D(_01604_),
    .Q(\core.registers[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20689_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01605_),
    .Q(\core.registers[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20690_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_01606_),
    .Q(\core.registers[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20691_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01607_),
    .Q(\core.registers[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20692_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_01608_),
    .Q(\core.registers[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20693_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01609_),
    .Q(\core.registers[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20694_ (.CLK(clknet_leaf_74_wb_clk_i),
    .D(_01610_),
    .Q(\core.registers[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20695_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01611_),
    .Q(\core.registers[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20696_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01612_),
    .Q(\core.registers[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20697_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01613_),
    .Q(\core.registers[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20698_ (.CLK(clknet_leaf_194_wb_clk_i),
    .D(_01614_),
    .Q(\core.registers[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20699_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01615_),
    .Q(\core.registers[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20700_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01616_),
    .Q(\core.registers[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20701_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_01617_),
    .Q(\core.registers[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20702_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_01618_),
    .Q(\core.registers[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20703_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_01619_),
    .Q(\core.registers[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20704_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_01620_),
    .Q(\core.registers[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20705_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_01621_),
    .Q(\core.registers[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _20706_ (.CLK(clknet_leaf_195_wb_clk_i),
    .D(_01622_),
    .Q(\core.registers[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _20707_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01623_),
    .Q(\core.registers[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _20708_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_01624_),
    .Q(\core.registers[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _20709_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01625_),
    .Q(\core.registers[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _20710_ (.CLK(clknet_leaf_213_wb_clk_i),
    .D(_01626_),
    .Q(\core.registers[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _20711_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_01627_),
    .Q(\core.registers[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _20712_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_01628_),
    .Q(\core.registers[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _20713_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_01629_),
    .Q(\core.registers[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _20714_ (.CLK(clknet_leaf_216_wb_clk_i),
    .D(_01630_),
    .Q(\core.registers[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _20715_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_01631_),
    .Q(\core.registers[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _20716_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_01632_),
    .Q(\core.registers[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _20717_ (.CLK(clknet_leaf_209_wb_clk_i),
    .D(_01633_),
    .Q(\core.registers[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _20718_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_01634_),
    .Q(\core.registers[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _20719_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_01635_),
    .Q(\core.registers[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _20720_ (.CLK(clknet_leaf_59_wb_clk_i),
    .D(_01636_),
    .Q(\core.registers[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _20721_ (.CLK(clknet_leaf_85_wb_clk_i),
    .D(_01637_),
    .Q(net482));
 sky130_fd_sc_hd__dfxtp_1 _20722_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_01638_),
    .Q(\core.csr.instretTimer.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20723_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_01639_),
    .Q(\core.csr.instretTimer.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20724_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_01640_),
    .Q(\core.csr.instretTimer.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20725_ (.CLK(clknet_leaf_101_wb_clk_i),
    .D(_01641_),
    .Q(\core.csr.instretTimer.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20726_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01642_),
    .Q(\core.csr.instretTimer.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20727_ (.CLK(clknet_leaf_97_wb_clk_i),
    .D(_01643_),
    .Q(\core.csr.instretTimer.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20728_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_01644_),
    .Q(\core.csr.instretTimer.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20729_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01645_),
    .Q(\core.csr.instretTimer.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20730_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01646_),
    .Q(\core.csr.instretTimer.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20731_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01647_),
    .Q(\core.csr.instretTimer.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20732_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01648_),
    .Q(\core.csr.instretTimer.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20733_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01649_),
    .Q(\core.csr.instretTimer.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20734_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01650_),
    .Q(\core.csr.instretTimer.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20735_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01651_),
    .Q(\core.csr.instretTimer.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20736_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01652_),
    .Q(\core.csr.instretTimer.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20737_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01653_),
    .Q(\core.csr.instretTimer.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20738_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01654_),
    .Q(\core.csr.instretTimer.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20739_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01655_),
    .Q(\core.csr.instretTimer.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20740_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01656_),
    .Q(\core.csr.instretTimer.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20741_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_01657_),
    .Q(\core.csr.instretTimer.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20742_ (.CLK(clknet_leaf_158_wb_clk_i),
    .D(_01658_),
    .Q(\core.csr.instretTimer.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20743_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01659_),
    .Q(\core.csr.instretTimer.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20744_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01660_),
    .Q(\core.csr.instretTimer.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20745_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01661_),
    .Q(\core.csr.instretTimer.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20746_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01662_),
    .Q(\core.csr.instretTimer.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20747_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01663_),
    .Q(\core.csr.instretTimer.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20748_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01664_),
    .Q(\core.csr.instretTimer.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20749_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01665_),
    .Q(\core.csr.instretTimer.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20750_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_01666_),
    .Q(\core.csr.instretTimer.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20751_ (.CLK(clknet_leaf_121_wb_clk_i),
    .D(_01667_),
    .Q(\core.csr.instretTimer.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20752_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01668_),
    .Q(\core.csr.instretTimer.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20753_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01669_),
    .Q(\core.csr.instretTimer.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20754_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_01670_),
    .Q(\core.csr.instretTimer.currentValue[32] ));
 sky130_fd_sc_hd__dfxtp_1 _20755_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_01671_),
    .Q(\core.csr.instretTimer.currentValue[33] ));
 sky130_fd_sc_hd__dfxtp_1 _20756_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_01672_),
    .Q(\core.csr.instretTimer.currentValue[34] ));
 sky130_fd_sc_hd__dfxtp_1 _20757_ (.CLK(clknet_leaf_100_wb_clk_i),
    .D(_01673_),
    .Q(\core.csr.instretTimer.currentValue[35] ));
 sky130_fd_sc_hd__dfxtp_1 _20758_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01674_),
    .Q(\core.csr.instretTimer.currentValue[36] ));
 sky130_fd_sc_hd__dfxtp_1 _20759_ (.CLK(clknet_leaf_96_wb_clk_i),
    .D(_01675_),
    .Q(\core.csr.instretTimer.currentValue[37] ));
 sky130_fd_sc_hd__dfxtp_1 _20760_ (.CLK(clknet_leaf_98_wb_clk_i),
    .D(_01676_),
    .Q(\core.csr.instretTimer.currentValue[38] ));
 sky130_fd_sc_hd__dfxtp_1 _20761_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01677_),
    .Q(\core.csr.instretTimer.currentValue[39] ));
 sky130_fd_sc_hd__dfxtp_1 _20762_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01678_),
    .Q(\core.csr.instretTimer.currentValue[40] ));
 sky130_fd_sc_hd__dfxtp_1 _20763_ (.CLK(clknet_leaf_99_wb_clk_i),
    .D(_01679_),
    .Q(\core.csr.instretTimer.currentValue[41] ));
 sky130_fd_sc_hd__dfxtp_1 _20764_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01680_),
    .Q(\core.csr.instretTimer.currentValue[42] ));
 sky130_fd_sc_hd__dfxtp_1 _20765_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01681_),
    .Q(\core.csr.instretTimer.currentValue[43] ));
 sky130_fd_sc_hd__dfxtp_1 _20766_ (.CLK(clknet_leaf_107_wb_clk_i),
    .D(_01682_),
    .Q(\core.csr.instretTimer.currentValue[44] ));
 sky130_fd_sc_hd__dfxtp_1 _20767_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01683_),
    .Q(\core.csr.instretTimer.currentValue[45] ));
 sky130_fd_sc_hd__dfxtp_1 _20768_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01684_),
    .Q(\core.csr.instretTimer.currentValue[46] ));
 sky130_fd_sc_hd__dfxtp_1 _20769_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01685_),
    .Q(\core.csr.instretTimer.currentValue[47] ));
 sky130_fd_sc_hd__dfxtp_1 _20770_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01686_),
    .Q(\core.csr.instretTimer.currentValue[48] ));
 sky130_fd_sc_hd__dfxtp_2 _20771_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01687_),
    .Q(\core.csr.instretTimer.currentValue[49] ));
 sky130_fd_sc_hd__dfxtp_1 _20772_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01688_),
    .Q(\core.csr.instretTimer.currentValue[50] ));
 sky130_fd_sc_hd__dfxtp_1 _20773_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01689_),
    .Q(\core.csr.instretTimer.currentValue[51] ));
 sky130_fd_sc_hd__dfxtp_1 _20774_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01690_),
    .Q(\core.csr.instretTimer.currentValue[52] ));
 sky130_fd_sc_hd__dfxtp_1 _20775_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01691_),
    .Q(\core.csr.instretTimer.currentValue[53] ));
 sky130_fd_sc_hd__dfxtp_1 _20776_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01692_),
    .Q(\core.csr.instretTimer.currentValue[54] ));
 sky130_fd_sc_hd__dfxtp_1 _20777_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01693_),
    .Q(\core.csr.instretTimer.currentValue[55] ));
 sky130_fd_sc_hd__dfxtp_1 _20778_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01694_),
    .Q(\core.csr.instretTimer.currentValue[56] ));
 sky130_fd_sc_hd__dfxtp_1 _20779_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01695_),
    .Q(\core.csr.instretTimer.currentValue[57] ));
 sky130_fd_sc_hd__dfxtp_1 _20780_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01696_),
    .Q(\core.csr.instretTimer.currentValue[58] ));
 sky130_fd_sc_hd__dfxtp_1 _20781_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01697_),
    .Q(\core.csr.instretTimer.currentValue[59] ));
 sky130_fd_sc_hd__dfxtp_1 _20782_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_01698_),
    .Q(\core.csr.instretTimer.currentValue[60] ));
 sky130_fd_sc_hd__dfxtp_1 _20783_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_01699_),
    .Q(\core.csr.instretTimer.currentValue[61] ));
 sky130_fd_sc_hd__dfxtp_1 _20784_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01700_),
    .Q(\core.csr.instretTimer.currentValue[62] ));
 sky130_fd_sc_hd__dfxtp_1 _20785_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01701_),
    .Q(\core.csr.instretTimer.currentValue[63] ));
 sky130_fd_sc_hd__dfxtp_1 _20786_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_01702_),
    .Q(\core.csr.mconfigptr.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20787_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01703_),
    .Q(\core.csr.mconfigptr.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20788_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01704_),
    .Q(\core.csr.mconfigptr.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20789_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_01705_),
    .Q(\core.csr.mconfigptr.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20790_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01706_),
    .Q(\core.csr.mconfigptr.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20791_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01707_),
    .Q(\core.csr.mconfigptr.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20792_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_01708_),
    .Q(\core.csr.mconfigptr.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20793_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01709_),
    .Q(\core.csr.mconfigptr.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20794_ (.CLK(clknet_leaf_102_wb_clk_i),
    .D(_01710_),
    .Q(\core.csr.mconfigptr.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20795_ (.CLK(clknet_leaf_106_wb_clk_i),
    .D(_01711_),
    .Q(\core.csr.mconfigptr.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20796_ (.CLK(clknet_leaf_108_wb_clk_i),
    .D(_01712_),
    .Q(\core.csr.mconfigptr.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20797_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01713_),
    .Q(\core.csr.mconfigptr.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20798_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01714_),
    .Q(\core.csr.mconfigptr.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20799_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_01715_),
    .Q(\core.csr.mconfigptr.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20800_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01716_),
    .Q(\core.csr.mconfigptr.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20801_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01717_),
    .Q(\core.csr.mconfigptr.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20802_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01718_),
    .Q(\core.csr.mconfigptr.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20803_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01719_),
    .Q(\core.csr.mconfigptr.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20804_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_01720_),
    .Q(\core.csr.mconfigptr.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20805_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01721_),
    .Q(\core.csr.mconfigptr.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20806_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01722_),
    .Q(\core.csr.mconfigptr.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20807_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01723_),
    .Q(\core.csr.mconfigptr.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20808_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01724_),
    .Q(\core.csr.mconfigptr.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20809_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01725_),
    .Q(\core.csr.mconfigptr.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20810_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01726_),
    .Q(\core.csr.mconfigptr.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20811_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01727_),
    .Q(\core.csr.mconfigptr.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20812_ (.CLK(clknet_leaf_167_wb_clk_i),
    .D(_01728_),
    .Q(\core.csr.mconfigptr.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20813_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01729_),
    .Q(\core.csr.mconfigptr.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20814_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_01730_),
    .Q(\core.csr.mconfigptr.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20815_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01731_),
    .Q(\core.csr.mconfigptr.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20816_ (.CLK(clknet_leaf_120_wb_clk_i),
    .D(_01732_),
    .Q(\core.csr.mconfigptr.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20817_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01733_),
    .Q(\core.csr.mconfigptr.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20818_ (.CLK(clknet_leaf_103_wb_clk_i),
    .D(_01734_),
    .Q(\core.csr.traps.mscratch.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20819_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01735_),
    .Q(\core.csr.traps.mscratch.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20820_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01736_),
    .Q(\core.csr.traps.mscratch.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20821_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01737_),
    .Q(\core.csr.traps.mscratch.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20822_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01738_),
    .Q(\core.csr.traps.mscratch.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20823_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_01739_),
    .Q(\core.csr.traps.mscratch.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20824_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01740_),
    .Q(\core.csr.traps.mscratch.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20825_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01741_),
    .Q(\core.csr.traps.mscratch.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20826_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01742_),
    .Q(\core.csr.traps.mscratch.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20827_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01743_),
    .Q(\core.csr.traps.mscratch.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20828_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01744_),
    .Q(\core.csr.traps.mscratch.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20829_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01745_),
    .Q(\core.csr.traps.mscratch.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20830_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01746_),
    .Q(\core.csr.traps.mscratch.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20831_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01747_),
    .Q(\core.csr.traps.mscratch.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20832_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01748_),
    .Q(\core.csr.traps.mscratch.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20833_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_01749_),
    .Q(\core.csr.traps.mscratch.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20834_ (.CLK(clknet_leaf_161_wb_clk_i),
    .D(_01750_),
    .Q(\core.csr.traps.mscratch.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20835_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01751_),
    .Q(\core.csr.traps.mscratch.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20836_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01752_),
    .Q(\core.csr.traps.mscratch.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20837_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01753_),
    .Q(\core.csr.traps.mscratch.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20838_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01754_),
    .Q(\core.csr.traps.mscratch.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20839_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_01755_),
    .Q(\core.csr.traps.mscratch.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20840_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_01756_),
    .Q(\core.csr.traps.mscratch.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20841_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_01757_),
    .Q(\core.csr.traps.mscratch.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20842_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01758_),
    .Q(\core.csr.traps.mscratch.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20843_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01759_),
    .Q(\core.csr.traps.mscratch.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20844_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01760_),
    .Q(\core.csr.traps.mscratch.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20845_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01761_),
    .Q(\core.csr.traps.mscratch.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20846_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01762_),
    .Q(\core.csr.traps.mscratch.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20847_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01763_),
    .Q(\core.csr.traps.mscratch.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20848_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01764_),
    .Q(\core.csr.traps.mscratch.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20849_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01765_),
    .Q(\core.csr.traps.mscratch.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20850_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_01766_),
    .Q(\core.csr.traps.mie.currentValue[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20851_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01767_),
    .Q(\core.csr.traps.mie.currentValue[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20852_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01768_),
    .Q(\core.csr.traps.mie.currentValue[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20853_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_01769_),
    .Q(\core.csr.traps.mie.currentValue[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20854_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01770_),
    .Q(\core.csr.traps.mie.currentValue[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20855_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01771_),
    .Q(\core.csr.traps.mie.currentValue[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20856_ (.CLK(clknet_leaf_104_wb_clk_i),
    .D(_01772_),
    .Q(\core.csr.traps.mie.currentValue[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20857_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01773_),
    .Q(\core.csr.traps.mie.currentValue[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20858_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01774_),
    .Q(\core.csr.traps.mie.currentValue[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20859_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01775_),
    .Q(\core.csr.traps.mie.currentValue[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20860_ (.CLK(clknet_leaf_109_wb_clk_i),
    .D(_01776_),
    .Q(\core.csr.traps.mie.currentValue[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20861_ (.CLK(clknet_leaf_105_wb_clk_i),
    .D(_01777_),
    .Q(\core.csr.traps.mie.currentValue[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20862_ (.CLK(clknet_leaf_111_wb_clk_i),
    .D(_01778_),
    .Q(\core.csr.traps.mie.currentValue[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20863_ (.CLK(clknet_leaf_115_wb_clk_i),
    .D(_01779_),
    .Q(\core.csr.traps.mie.currentValue[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20864_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01780_),
    .Q(\core.csr.traps.mie.currentValue[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20865_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01781_),
    .Q(\core.csr.traps.mie.currentValue[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20866_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_01782_),
    .Q(\core.csr.traps.mie.currentValue[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20867_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01783_),
    .Q(\core.csr.traps.mie.currentValue[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20868_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01784_),
    .Q(\core.csr.traps.mie.currentValue[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20869_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01785_),
    .Q(\core.csr.traps.mie.currentValue[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20870_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01786_),
    .Q(\core.csr.traps.mie.currentValue[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20871_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_01787_),
    .Q(\core.csr.traps.mie.currentValue[21] ));
 sky130_fd_sc_hd__dfxtp_1 _20872_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_01788_),
    .Q(\core.csr.traps.mie.currentValue[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20873_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_01789_),
    .Q(\core.csr.traps.mie.currentValue[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20874_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_01790_),
    .Q(\core.csr.traps.mie.currentValue[24] ));
 sky130_fd_sc_hd__dfxtp_1 _20875_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01791_),
    .Q(\core.csr.traps.mie.currentValue[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20876_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01792_),
    .Q(\core.csr.traps.mie.currentValue[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20877_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01793_),
    .Q(\core.csr.traps.mie.currentValue[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20878_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01794_),
    .Q(\core.csr.traps.mie.currentValue[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20879_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01795_),
    .Q(\core.csr.traps.mie.currentValue[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20880_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01796_),
    .Q(\core.csr.traps.mie.currentValue[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20881_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01797_),
    .Q(\core.csr.traps.mie.currentValue[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20882_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01798_),
    .Q(\core.csr.traps.mcause.csrReadData[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20883_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01799_),
    .Q(\core.csr.traps.mcause.csrReadData[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20884_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01800_),
    .Q(\core.csr.traps.mcause.csrReadData[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20885_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01801_),
    .Q(\core.csr.traps.mcause.csrReadData[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20886_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01802_),
    .Q(\core.csr.traps.mcause.csrReadData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20887_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01803_),
    .Q(\core.csr.traps.mcause.csrReadData[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20888_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01804_),
    .Q(\core.csr.traps.mcause.csrReadData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20889_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01805_),
    .Q(\core.csr.traps.mcause.csrReadData[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20890_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01806_),
    .Q(\core.csr.traps.mcause.csrReadData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20891_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01807_),
    .Q(\core.csr.traps.mcause.csrReadData[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20892_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01808_),
    .Q(\core.csr.traps.mcause.csrReadData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20893_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01809_),
    .Q(\core.csr.traps.mcause.csrReadData[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20894_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01810_),
    .Q(\core.csr.traps.mcause.csrReadData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20895_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01811_),
    .Q(\core.csr.traps.mcause.csrReadData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20896_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01812_),
    .Q(\core.csr.traps.mcause.csrReadData[14] ));
 sky130_fd_sc_hd__dfxtp_4 _20897_ (.CLK(clknet_leaf_161_wb_clk_i),
    .D(_01813_),
    .Q(\core.csr.traps.mcause.csrReadData[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20898_ (.CLK(clknet_leaf_161_wb_clk_i),
    .D(_01814_),
    .Q(\core.csr.traps.mcause.csrReadData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20899_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01815_),
    .Q(\core.csr.traps.mcause.csrReadData[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20900_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01816_),
    .Q(\core.csr.traps.mcause.csrReadData[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20901_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01817_),
    .Q(\core.csr.traps.mcause.csrReadData[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20902_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01818_),
    .Q(\core.csr.traps.mcause.csrReadData[20] ));
 sky130_fd_sc_hd__dfxtp_1 _20903_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01819_),
    .Q(\core.csr.traps.mcause.csrReadData[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20904_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01820_),
    .Q(\core.csr.traps.mcause.csrReadData[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20905_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01821_),
    .Q(\core.csr.traps.mcause.csrReadData[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20906_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01822_),
    .Q(\core.csr.traps.mcause.csrReadData[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20907_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_01823_),
    .Q(\core.csr.traps.mcause.csrReadData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _20908_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01824_),
    .Q(\core.csr.traps.mcause.csrReadData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _20909_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01825_),
    .Q(\core.csr.traps.mcause.csrReadData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _20910_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01826_),
    .Q(\core.csr.traps.mcause.csrReadData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20911_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_01827_),
    .Q(\core.csr.traps.mcause.csrReadData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _20912_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01828_),
    .Q(\core.csr.traps.mcause.csrReadData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _20913_ (.CLK(clknet_leaf_163_wb_clk_i),
    .D(_01829_),
    .Q(\core.csr.traps.mcause.csrReadData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20914_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01830_),
    .Q(\core.csr.trapReturnVector[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20915_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01831_),
    .Q(\core.csr.trapReturnVector[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20916_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01832_),
    .Q(\core.csr.trapReturnVector[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20917_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01833_),
    .Q(\core.csr.trapReturnVector[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20918_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01834_),
    .Q(\core.csr.trapReturnVector[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20919_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_01835_),
    .Q(\core.csr.trapReturnVector[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20920_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01836_),
    .Q(\core.csr.trapReturnVector[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20921_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01837_),
    .Q(\core.csr.trapReturnVector[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20922_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01838_),
    .Q(\core.csr.trapReturnVector[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20923_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01839_),
    .Q(\core.csr.trapReturnVector[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20924_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01840_),
    .Q(\core.csr.trapReturnVector[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20925_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01841_),
    .Q(\core.csr.trapReturnVector[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20926_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01842_),
    .Q(\core.csr.trapReturnVector[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20927_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01843_),
    .Q(\core.csr.trapReturnVector[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20928_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01844_),
    .Q(\core.csr.trapReturnVector[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20929_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01845_),
    .Q(\core.csr.trapReturnVector[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20930_ (.CLK(clknet_leaf_147_wb_clk_i),
    .D(_01846_),
    .Q(\core.csr.trapReturnVector[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20931_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01847_),
    .Q(\core.csr.trapReturnVector[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20932_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01848_),
    .Q(\core.csr.trapReturnVector[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20933_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01849_),
    .Q(\core.csr.trapReturnVector[19] ));
 sky130_fd_sc_hd__dfxtp_1 _20934_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01850_),
    .Q(\core.csr.trapReturnVector[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20935_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01851_),
    .Q(\core.csr.trapReturnVector[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20936_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01852_),
    .Q(\core.csr.trapReturnVector[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20937_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01853_),
    .Q(\core.csr.trapReturnVector[23] ));
 sky130_fd_sc_hd__dfxtp_1 _20938_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01854_),
    .Q(\core.csr.trapReturnVector[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20939_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_01855_),
    .Q(\core.csr.trapReturnVector[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20940_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01856_),
    .Q(\core.csr.trapReturnVector[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20941_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01857_),
    .Q(\core.csr.trapReturnVector[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20942_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01858_),
    .Q(\core.csr.trapReturnVector[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20943_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_01859_),
    .Q(\core.csr.trapReturnVector[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20944_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01860_),
    .Q(\core.csr.trapReturnVector[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20945_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_01861_),
    .Q(\core.csr.trapReturnVector[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20946_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01862_),
    .Q(\core.csr.traps.mtvec.csrReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20947_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01863_),
    .Q(\core.csr.traps.mtvec.csrReadData[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20948_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01864_),
    .Q(\core.csr.traps.mtvec.csrReadData[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20949_ (.CLK(clknet_leaf_118_wb_clk_i),
    .D(_01865_),
    .Q(\core.csr.traps.mtvec.csrReadData[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20950_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01866_),
    .Q(\core.csr.traps.mtvec.csrReadData[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20951_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_01867_),
    .Q(\core.csr.traps.mtvec.csrReadData[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20952_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01868_),
    .Q(\core.csr.traps.mtvec.csrReadData[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20953_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01869_),
    .Q(\core.csr.traps.mtvec.csrReadData[7] ));
 sky130_fd_sc_hd__dfxtp_4 _20954_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01870_),
    .Q(\core.csr.traps.mtvec.csrReadData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20955_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01871_),
    .Q(\core.csr.traps.mtvec.csrReadData[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20956_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01872_),
    .Q(\core.csr.traps.mtvec.csrReadData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20957_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01873_),
    .Q(\core.csr.traps.mtvec.csrReadData[11] ));
 sky130_fd_sc_hd__dfxtp_4 _20958_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01874_),
    .Q(\core.csr.traps.mtvec.csrReadData[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20959_ (.CLK(clknet_leaf_151_wb_clk_i),
    .D(_01875_),
    .Q(\core.csr.traps.mtvec.csrReadData[13] ));
 sky130_fd_sc_hd__dfxtp_4 _20960_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01876_),
    .Q(\core.csr.traps.mtvec.csrReadData[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20961_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_01877_),
    .Q(\core.csr.traps.mtvec.csrReadData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20962_ (.CLK(clknet_leaf_157_wb_clk_i),
    .D(_01878_),
    .Q(\core.csr.traps.mtvec.csrReadData[16] ));
 sky130_fd_sc_hd__dfxtp_4 _20963_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01879_),
    .Q(\core.csr.traps.mtvec.csrReadData[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20964_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01880_),
    .Q(\core.csr.traps.mtvec.csrReadData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20965_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01881_),
    .Q(\core.csr.traps.mtvec.csrReadData[19] ));
 sky130_fd_sc_hd__dfxtp_4 _20966_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01882_),
    .Q(\core.csr.traps.mtvec.csrReadData[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20967_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01883_),
    .Q(\core.csr.traps.mtvec.csrReadData[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20968_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01884_),
    .Q(\core.csr.traps.mtvec.csrReadData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20969_ (.CLK(clknet_leaf_171_wb_clk_i),
    .D(_01885_),
    .Q(\core.csr.traps.mtvec.csrReadData[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20970_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01886_),
    .Q(\core.csr.traps.mtvec.csrReadData[24] ));
 sky130_fd_sc_hd__dfxtp_4 _20971_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01887_),
    .Q(\core.csr.traps.mtvec.csrReadData[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20972_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01888_),
    .Q(\core.csr.traps.mtvec.csrReadData[26] ));
 sky130_fd_sc_hd__dfxtp_4 _20973_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01889_),
    .Q(\core.csr.traps.mtvec.csrReadData[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20974_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01890_),
    .Q(\core.csr.traps.mtvec.csrReadData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _20975_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01891_),
    .Q(\core.csr.traps.mtvec.csrReadData[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20976_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01892_),
    .Q(\core.csr.traps.mtvec.csrReadData[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20977_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01893_),
    .Q(\core.csr.traps.mtvec.csrReadData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _20978_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01894_),
    .Q(\core.csr.traps.machineInterruptEnable ));
 sky130_fd_sc_hd__dfxtp_2 _20979_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01895_),
    .Q(\core.csr.traps.machinePreviousInterruptEnable ));
 sky130_fd_sc_hd__dfxtp_1 _20980_ (.CLK(clknet_leaf_133_wb_clk_i),
    .D(_01896_),
    .Q(\core.csr.traps.mtval.csrReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20981_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01897_),
    .Q(\core.csr.traps.mtval.csrReadData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20982_ (.CLK(clknet_leaf_132_wb_clk_i),
    .D(_01898_),
    .Q(\core.csr.traps.mtval.csrReadData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20983_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01899_),
    .Q(\core.csr.traps.mtval.csrReadData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20984_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01900_),
    .Q(\core.csr.traps.mtval.csrReadData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20985_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_01901_),
    .Q(\core.csr.traps.mtval.csrReadData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20986_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01902_),
    .Q(\core.csr.traps.mtval.csrReadData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20987_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01903_),
    .Q(\core.csr.traps.mtval.csrReadData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20988_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01904_),
    .Q(\core.csr.traps.mtval.csrReadData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20989_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01905_),
    .Q(\core.csr.traps.mtval.csrReadData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20990_ (.CLK(clknet_leaf_153_wb_clk_i),
    .D(_01906_),
    .Q(\core.csr.traps.mtval.csrReadData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20991_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01907_),
    .Q(\core.csr.traps.mtval.csrReadData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _20992_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01908_),
    .Q(\core.csr.traps.mtval.csrReadData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _20993_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01909_),
    .Q(\core.csr.traps.mtval.csrReadData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _20994_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01910_),
    .Q(\core.csr.traps.mtval.csrReadData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20995_ (.CLK(clknet_leaf_161_wb_clk_i),
    .D(_01911_),
    .Q(\core.csr.traps.mtval.csrReadData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20996_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01912_),
    .Q(\core.csr.traps.mtval.csrReadData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _20997_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01913_),
    .Q(\core.csr.traps.mtval.csrReadData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _20998_ (.CLK(clknet_leaf_162_wb_clk_i),
    .D(_01914_),
    .Q(\core.csr.traps.mtval.csrReadData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _20999_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01915_),
    .Q(\core.csr.traps.mtval.csrReadData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21000_ (.CLK(clknet_leaf_172_wb_clk_i),
    .D(_01916_),
    .Q(\core.csr.traps.mtval.csrReadData[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21001_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01917_),
    .Q(\core.csr.traps.mtval.csrReadData[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21002_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01918_),
    .Q(\core.csr.traps.mtval.csrReadData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21003_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01919_),
    .Q(\core.csr.traps.mtval.csrReadData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21004_ (.CLK(clknet_leaf_174_wb_clk_i),
    .D(_01920_),
    .Q(\core.csr.traps.mtval.csrReadData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21005_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_01921_),
    .Q(\core.csr.traps.mtval.csrReadData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21006_ (.CLK(clknet_leaf_165_wb_clk_i),
    .D(_01922_),
    .Q(\core.csr.traps.mtval.csrReadData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21007_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01923_),
    .Q(\core.csr.traps.mtval.csrReadData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21008_ (.CLK(clknet_leaf_175_wb_clk_i),
    .D(_01924_),
    .Q(\core.csr.traps.mtval.csrReadData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21009_ (.CLK(clknet_leaf_176_wb_clk_i),
    .D(_01925_),
    .Q(\core.csr.traps.mtval.csrReadData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21010_ (.CLK(clknet_leaf_173_wb_clk_i),
    .D(_01926_),
    .Q(\core.csr.traps.mtval.csrReadData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21011_ (.CLK(clknet_leaf_164_wb_clk_i),
    .D(_01927_),
    .Q(\core.csr.traps.mtval.csrReadData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21012_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01928_),
    .Q(\core.csr.traps.mip.csrReadData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21013_ (.CLK(clknet_leaf_117_wb_clk_i),
    .D(_01929_),
    .Q(\core.csr.traps.mip.csrReadData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21014_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01930_),
    .Q(\core.csr.traps.mip.csrReadData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21015_ (.CLK(clknet_leaf_131_wb_clk_i),
    .D(_01931_),
    .Q(\core.csr.traps.mip.csrReadData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21016_ (.CLK(clknet_leaf_119_wb_clk_i),
    .D(_01932_),
    .Q(\core.csr.traps.mip.csrReadData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21017_ (.CLK(clknet_leaf_128_wb_clk_i),
    .D(_01933_),
    .Q(\core.csr.traps.mip.csrReadData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21018_ (.CLK(clknet_leaf_116_wb_clk_i),
    .D(_01934_),
    .Q(\core.csr.traps.mip.csrReadData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21019_ (.CLK(clknet_leaf_129_wb_clk_i),
    .D(_01935_),
    .Q(\core.csr.traps.mip.csrReadData[7] ));
 sky130_fd_sc_hd__dfxtp_2 _21020_ (.CLK(clknet_leaf_114_wb_clk_i),
    .D(_01936_),
    .Q(\core.csr.traps.mip.csrReadData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21021_ (.CLK(clknet_leaf_130_wb_clk_i),
    .D(_01937_),
    .Q(\core.csr.traps.mip.csrReadData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21022_ (.CLK(clknet_leaf_127_wb_clk_i),
    .D(_01938_),
    .Q(\core.csr.traps.mip.csrReadData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21023_ (.CLK(clknet_leaf_150_wb_clk_i),
    .D(_01939_),
    .Q(\core.csr.traps.mip.csrReadData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21024_ (.CLK(clknet_leaf_152_wb_clk_i),
    .D(_01940_),
    .Q(\core.csr.traps.mip.csrReadData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21025_ (.CLK(clknet_leaf_148_wb_clk_i),
    .D(_01941_),
    .Q(\core.csr.traps.mip.csrReadData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21026_ (.CLK(clknet_leaf_156_wb_clk_i),
    .D(_01942_),
    .Q(\core.csr.traps.mip.csrReadData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21027_ (.CLK(clknet_leaf_161_wb_clk_i),
    .D(_01943_),
    .Q(\core.csr.traps.mip.csrReadData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21028_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01944_),
    .Q(\core.csr.traps.mip.csrReadData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21029_ (.CLK(clknet_leaf_159_wb_clk_i),
    .D(_01945_),
    .Q(\core.csr.traps.mip.csrReadData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21030_ (.CLK(clknet_leaf_160_wb_clk_i),
    .D(_01946_),
    .Q(\core.csr.traps.mip.csrReadData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21031_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01947_),
    .Q(\core.csr.traps.mip.csrReadData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21032_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01948_),
    .Q(\core.csr.traps.mip.csrReadData[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21033_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_01949_),
    .Q(\core.csr.traps.mip.csrReadData[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21034_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_01950_),
    .Q(\core.csr.traps.mip.csrReadData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21035_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_01951_),
    .Q(\core.csr.traps.mip.csrReadData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21036_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_01952_),
    .Q(\core.csr.traps.mip.csrReadData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21037_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01953_),
    .Q(\core.csr.traps.mip.csrReadData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21038_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01954_),
    .Q(\core.csr.traps.mip.csrReadData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21039_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01955_),
    .Q(\core.csr.traps.mip.csrReadData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21040_ (.CLK(clknet_leaf_169_wb_clk_i),
    .D(_01956_),
    .Q(\core.csr.traps.mip.csrReadData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21041_ (.CLK(clknet_leaf_168_wb_clk_i),
    .D(_01957_),
    .Q(\core.csr.traps.mip.csrReadData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21042_ (.CLK(clknet_leaf_170_wb_clk_i),
    .D(_01958_),
    .Q(\core.csr.traps.mip.csrReadData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21043_ (.CLK(clknet_leaf_166_wb_clk_i),
    .D(_01959_),
    .Q(\core.csr.traps.mip.csrReadData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21044_ (.CLK(clknet_leaf_87_wb_clk_i),
    .D(_01960_),
    .Q(\core.pipe2_stall ));
 sky130_fd_sc_hd__buf_2 _21046_ (.A(clknet_leaf_218_wb_clk_i),
    .X(net303));
 sky130_fd_sc_hd__buf_2 _21047_ (.A(clknet_leaf_39_wb_clk_i),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.A(clknet_3_0_0_wb_clk_i),
    .X(clknet_4_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.A(clknet_3_5_0_wb_clk_i),
    .X(clknet_4_10__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.A(clknet_3_5_0_wb_clk_i),
    .X(clknet_4_11__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.A(clknet_3_6_0_wb_clk_i),
    .X(clknet_4_12__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.A(clknet_3_6_0_wb_clk_i),
    .X(clknet_4_13__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.A(clknet_3_7_0_wb_clk_i),
    .X(clknet_4_14__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.A(clknet_3_7_0_wb_clk_i),
    .X(clknet_4_15__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.A(clknet_3_0_0_wb_clk_i),
    .X(clknet_4_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.A(clknet_3_1_0_wb_clk_i),
    .X(clknet_4_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.A(clknet_3_1_0_wb_clk_i),
    .X(clknet_4_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.A(clknet_3_2_0_wb_clk_i),
    .X(clknet_4_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.A(clknet_3_2_0_wb_clk_i),
    .X(clknet_4_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.A(clknet_3_3_0_wb_clk_i),
    .X(clknet_4_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.A(clknet_3_3_0_wb_clk_i),
    .X(clknet_4_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.A(clknet_3_4_0_wb_clk_i),
    .X(clknet_4_8__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.A(clknet_3_4_0_wb_clk_i),
    .X(clknet_4_9__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_100_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_101_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_102_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_103_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_104_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_105_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_106_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_107_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_108_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_109_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_110_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_111_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_112_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_113_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_114_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.A(clknet_4_15__leaf_wb_clk_i),
    .X(clknet_leaf_115_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_116_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_117_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_118_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_119_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_120_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_121_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_122_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_123_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_124_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_125_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_126_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_127_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_128_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_129_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_130_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_131_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.A(clknet_4_13__leaf_wb_clk_i),
    .X(clknet_leaf_132_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_133_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_134_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_135_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_137_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_138_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_139_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_140_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_141_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_142_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_143_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_144_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_145_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_146_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_147_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_148_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_149_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_150_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_151_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_152_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_153_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_154_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_155_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_156_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_157_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_158_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_159_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_160_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_161_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_wb_clk_i (.A(clknet_4_7__leaf_wb_clk_i),
    .X(clknet_leaf_162_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_163_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_164_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_165_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_166_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_167_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_168_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_169_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_170_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_171_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_172_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_173_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_174_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_175_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_wb_clk_i (.A(clknet_4_5__leaf_wb_clk_i),
    .X(clknet_leaf_176_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_177_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_178_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_179_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_180_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_181_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_182_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_183_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_184_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_185_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_186_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_188_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_wb_clk_i (.A(clknet_4_4__leaf_wb_clk_i),
    .X(clknet_leaf_189_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_190_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_191_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_192_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_wb_clk_i (.A(clknet_4_6__leaf_wb_clk_i),
    .X(clknet_leaf_193_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_194_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_195_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_196_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_197_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_198_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_199_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_200_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_201_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_202_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_203_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_204_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_205_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_206_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_207_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_wb_clk_i (.A(clknet_4_1__leaf_wb_clk_i),
    .X(clknet_leaf_208_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_209_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_210_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_211_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_212_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_213_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_214_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_215_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_216_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_217_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_218_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_4_3__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_4_8__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_4_0__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_51_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_53_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_54_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_55_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_56_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_57_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_58_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.A(clknet_4_10__leaf_wb_clk_i),
    .X(clknet_leaf_59_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_60_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_61_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_62_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_63_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_64_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_65_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_66_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_67_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_68_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_69_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_70_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_71_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_72_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_73_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.A(clknet_4_11__leaf_wb_clk_i),
    .X(clknet_leaf_74_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_75_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_76_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_77_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_78_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_79_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.A(clknet_4_9__leaf_wb_clk_i),
    .X(clknet_leaf_80_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_81_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_82_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_83_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_84_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.A(clknet_4_12__leaf_wb_clk_i),
    .X(clknet_leaf_85_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_86_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_87_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_88_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_89_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_90_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_91_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_92_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_93_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_94_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_95_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_96_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_97_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_98_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.A(clknet_4_14__leaf_wb_clk_i),
    .X(clknet_leaf_99_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_4_2__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout1000 (.A(net1001),
    .X(net1000));
 sky130_fd_sc_hd__buf_8 fanout1001 (.A(_09244_),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_16 fanout1002 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_16 fanout1003 (.A(net1004),
    .X(net1003));
 sky130_fd_sc_hd__buf_8 fanout1004 (.A(net1005),
    .X(net1004));
 sky130_fd_sc_hd__buf_12 fanout1005 (.A(net1006),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_16 fanout1006 (.A(_09244_),
    .X(net1006));
 sky130_fd_sc_hd__buf_4 fanout1007 (.A(_09243_),
    .X(net1007));
 sky130_fd_sc_hd__buf_4 fanout1008 (.A(net1009),
    .X(net1008));
 sky130_fd_sc_hd__buf_4 fanout1009 (.A(net1011),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_8 fanout1010 (.A(net1011),
    .X(net1010));
 sky130_fd_sc_hd__buf_4 fanout1011 (.A(_09221_),
    .X(net1011));
 sky130_fd_sc_hd__buf_4 fanout1012 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 fanout1013 (.A(net1015),
    .X(net1013));
 sky130_fd_sc_hd__buf_6 fanout1014 (.A(net1015),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 fanout1015 (.A(_09220_),
    .X(net1015));
 sky130_fd_sc_hd__buf_4 fanout1016 (.A(net1017),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_4 fanout1017 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__buf_2 fanout1018 (.A(net1020),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_8 fanout1019 (.A(net1020),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_4 fanout1020 (.A(_07496_),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 fanout1021 (.A(net1024),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout1022 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__buf_6 fanout1023 (.A(net1024),
    .X(net1023));
 sky130_fd_sc_hd__buf_6 fanout1024 (.A(_03111_),
    .X(net1024));
 sky130_fd_sc_hd__buf_4 fanout1025 (.A(net1028),
    .X(net1025));
 sky130_fd_sc_hd__buf_4 fanout1026 (.A(net1027),
    .X(net1026));
 sky130_fd_sc_hd__buf_6 fanout1027 (.A(net1028),
    .X(net1027));
 sky130_fd_sc_hd__buf_6 fanout1028 (.A(_03102_),
    .X(net1028));
 sky130_fd_sc_hd__buf_4 fanout1029 (.A(_02338_),
    .X(net1029));
 sky130_fd_sc_hd__buf_2 fanout1030 (.A(_02338_),
    .X(net1030));
 sky130_fd_sc_hd__buf_4 fanout1031 (.A(net1032),
    .X(net1031));
 sky130_fd_sc_hd__buf_4 fanout1032 (.A(_09242_),
    .X(net1032));
 sky130_fd_sc_hd__buf_4 fanout1033 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__buf_6 fanout1034 (.A(_09241_),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_4 fanout1035 (.A(net1037),
    .X(net1035));
 sky130_fd_sc_hd__clkbuf_2 fanout1036 (.A(net1037),
    .X(net1036));
 sky130_fd_sc_hd__buf_4 fanout1037 (.A(net1038),
    .X(net1037));
 sky130_fd_sc_hd__buf_4 fanout1038 (.A(_06160_),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_4 fanout1039 (.A(net1040),
    .X(net1039));
 sky130_fd_sc_hd__buf_2 fanout1040 (.A(net1042),
    .X(net1040));
 sky130_fd_sc_hd__buf_8 fanout1041 (.A(net1042),
    .X(net1041));
 sky130_fd_sc_hd__buf_6 fanout1042 (.A(_06065_),
    .X(net1042));
 sky130_fd_sc_hd__buf_4 fanout1043 (.A(net1046),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_4 fanout1044 (.A(net1046),
    .X(net1044));
 sky130_fd_sc_hd__buf_2 fanout1045 (.A(net1046),
    .X(net1045));
 sky130_fd_sc_hd__clkbuf_4 fanout1046 (.A(net1047),
    .X(net1046));
 sky130_fd_sc_hd__buf_8 fanout1047 (.A(_05976_),
    .X(net1047));
 sky130_fd_sc_hd__buf_4 fanout1048 (.A(net1052),
    .X(net1048));
 sky130_fd_sc_hd__clkbuf_2 fanout1049 (.A(net1052),
    .X(net1049));
 sky130_fd_sc_hd__buf_4 fanout1050 (.A(net1051),
    .X(net1050));
 sky130_fd_sc_hd__buf_2 fanout1051 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__buf_4 fanout1052 (.A(_05891_),
    .X(net1052));
 sky130_fd_sc_hd__buf_4 fanout1053 (.A(_05807_),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_4 fanout1054 (.A(_05807_),
    .X(net1054));
 sky130_fd_sc_hd__clkbuf_4 fanout1055 (.A(net1056),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_2 fanout1056 (.A(_05807_),
    .X(net1056));
 sky130_fd_sc_hd__clkbuf_4 fanout1057 (.A(net1060),
    .X(net1057));
 sky130_fd_sc_hd__clkbuf_4 fanout1058 (.A(net1060),
    .X(net1058));
 sky130_fd_sc_hd__buf_6 fanout1059 (.A(_05726_),
    .X(net1059));
 sky130_fd_sc_hd__buf_2 fanout1060 (.A(_05726_),
    .X(net1060));
 sky130_fd_sc_hd__buf_4 fanout1061 (.A(net1063),
    .X(net1061));
 sky130_fd_sc_hd__buf_2 fanout1062 (.A(net1063),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_8 fanout1063 (.A(_05641_),
    .X(net1063));
 sky130_fd_sc_hd__buf_6 fanout1064 (.A(_05641_),
    .X(net1064));
 sky130_fd_sc_hd__buf_6 fanout1065 (.A(net1067),
    .X(net1065));
 sky130_fd_sc_hd__buf_12 fanout1066 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__buf_6 fanout1067 (.A(_04662_),
    .X(net1067));
 sky130_fd_sc_hd__buf_4 fanout1068 (.A(net1069),
    .X(net1068));
 sky130_fd_sc_hd__buf_4 fanout1069 (.A(_04661_),
    .X(net1069));
 sky130_fd_sc_hd__buf_8 fanout1070 (.A(net1071),
    .X(net1070));
 sky130_fd_sc_hd__buf_6 fanout1071 (.A(_04661_),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_4 fanout1072 (.A(net1074),
    .X(net1072));
 sky130_fd_sc_hd__clkbuf_2 fanout1073 (.A(net1074),
    .X(net1073));
 sky130_fd_sc_hd__buf_2 fanout1074 (.A(_09085_),
    .X(net1074));
 sky130_fd_sc_hd__clkbuf_4 fanout1075 (.A(_09085_),
    .X(net1075));
 sky130_fd_sc_hd__buf_6 fanout1076 (.A(net1078),
    .X(net1076));
 sky130_fd_sc_hd__buf_6 fanout1077 (.A(net1078),
    .X(net1077));
 sky130_fd_sc_hd__buf_12 fanout1078 (.A(net443),
    .X(net1078));
 sky130_fd_sc_hd__buf_6 fanout1079 (.A(_07490_),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_4 fanout1080 (.A(_07490_),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_8 fanout1081 (.A(net1083),
    .X(net1081));
 sky130_fd_sc_hd__buf_2 fanout1082 (.A(net1083),
    .X(net1082));
 sky130_fd_sc_hd__buf_6 fanout1083 (.A(_07489_),
    .X(net1083));
 sky130_fd_sc_hd__buf_4 fanout1084 (.A(net1086),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_2 fanout1085 (.A(net1086),
    .X(net1085));
 sky130_fd_sc_hd__buf_4 fanout1086 (.A(net1087),
    .X(net1086));
 sky130_fd_sc_hd__buf_8 fanout1087 (.A(_07280_),
    .X(net1087));
 sky130_fd_sc_hd__clkbuf_4 fanout1088 (.A(net1089),
    .X(net1088));
 sky130_fd_sc_hd__buf_4 fanout1089 (.A(net1090),
    .X(net1089));
 sky130_fd_sc_hd__buf_6 fanout1090 (.A(net1091),
    .X(net1090));
 sky130_fd_sc_hd__buf_8 fanout1091 (.A(_07206_),
    .X(net1091));
 sky130_fd_sc_hd__clkbuf_4 fanout1092 (.A(net1094),
    .X(net1092));
 sky130_fd_sc_hd__clkbuf_2 fanout1093 (.A(net1094),
    .X(net1093));
 sky130_fd_sc_hd__buf_6 fanout1094 (.A(_07123_),
    .X(net1094));
 sky130_fd_sc_hd__buf_6 fanout1095 (.A(_07123_),
    .X(net1095));
 sky130_fd_sc_hd__buf_4 fanout1096 (.A(net1097),
    .X(net1096));
 sky130_fd_sc_hd__buf_4 fanout1097 (.A(_07069_),
    .X(net1097));
 sky130_fd_sc_hd__buf_4 fanout1098 (.A(net1099),
    .X(net1098));
 sky130_fd_sc_hd__buf_4 fanout1099 (.A(_07069_),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_4 fanout1100 (.A(net1101),
    .X(net1100));
 sky130_fd_sc_hd__clkbuf_2 fanout1101 (.A(net1102),
    .X(net1101));
 sky130_fd_sc_hd__buf_4 fanout1102 (.A(net1103),
    .X(net1102));
 sky130_fd_sc_hd__buf_6 fanout1103 (.A(_06953_),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_4 fanout1104 (.A(net1106),
    .X(net1104));
 sky130_fd_sc_hd__clkbuf_2 fanout1105 (.A(net1106),
    .X(net1105));
 sky130_fd_sc_hd__buf_4 fanout1106 (.A(net1107),
    .X(net1106));
 sky130_fd_sc_hd__buf_4 fanout1107 (.A(_06877_),
    .X(net1107));
 sky130_fd_sc_hd__buf_4 fanout1108 (.A(net1109),
    .X(net1108));
 sky130_fd_sc_hd__buf_4 fanout1109 (.A(net1111),
    .X(net1109));
 sky130_fd_sc_hd__clkbuf_4 fanout1110 (.A(net1111),
    .X(net1110));
 sky130_fd_sc_hd__buf_6 fanout1111 (.A(_06799_),
    .X(net1111));
 sky130_fd_sc_hd__clkbuf_4 fanout1112 (.A(net1113),
    .X(net1112));
 sky130_fd_sc_hd__buf_2 fanout1113 (.A(_06720_),
    .X(net1113));
 sky130_fd_sc_hd__buf_4 fanout1114 (.A(net1115),
    .X(net1114));
 sky130_fd_sc_hd__buf_4 fanout1115 (.A(_06720_),
    .X(net1115));
 sky130_fd_sc_hd__clkbuf_4 fanout1116 (.A(net1118),
    .X(net1116));
 sky130_fd_sc_hd__clkbuf_4 fanout1117 (.A(net1118),
    .X(net1117));
 sky130_fd_sc_hd__buf_4 fanout1118 (.A(net1119),
    .X(net1118));
 sky130_fd_sc_hd__clkbuf_4 fanout1119 (.A(_06602_),
    .X(net1119));
 sky130_fd_sc_hd__clkbuf_4 fanout1120 (.A(net1121),
    .X(net1120));
 sky130_fd_sc_hd__buf_4 fanout1121 (.A(net1122),
    .X(net1121));
 sky130_fd_sc_hd__buf_4 fanout1122 (.A(net1123),
    .X(net1122));
 sky130_fd_sc_hd__clkbuf_4 fanout1123 (.A(_06525_),
    .X(net1123));
 sky130_fd_sc_hd__clkbuf_4 fanout1124 (.A(net1126),
    .X(net1124));
 sky130_fd_sc_hd__clkbuf_2 fanout1125 (.A(net1126),
    .X(net1125));
 sky130_fd_sc_hd__clkbuf_4 fanout1126 (.A(net1127),
    .X(net1126));
 sky130_fd_sc_hd__clkbuf_4 fanout1127 (.A(_06447_),
    .X(net1127));
 sky130_fd_sc_hd__buf_4 fanout1128 (.A(net1130),
    .X(net1128));
 sky130_fd_sc_hd__buf_4 fanout1129 (.A(net1130),
    .X(net1129));
 sky130_fd_sc_hd__buf_2 fanout1130 (.A(net1131),
    .X(net1130));
 sky130_fd_sc_hd__buf_4 fanout1131 (.A(_06367_),
    .X(net1131));
 sky130_fd_sc_hd__buf_4 fanout1132 (.A(net1133),
    .X(net1132));
 sky130_fd_sc_hd__buf_4 fanout1133 (.A(net1134),
    .X(net1133));
 sky130_fd_sc_hd__buf_4 fanout1134 (.A(net1135),
    .X(net1134));
 sky130_fd_sc_hd__buf_8 fanout1135 (.A(_05594_),
    .X(net1135));
 sky130_fd_sc_hd__clkbuf_4 fanout1136 (.A(_04860_),
    .X(net1136));
 sky130_fd_sc_hd__clkbuf_2 fanout1137 (.A(_04860_),
    .X(net1137));
 sky130_fd_sc_hd__clkbuf_8 fanout1138 (.A(_04860_),
    .X(net1138));
 sky130_fd_sc_hd__clkbuf_4 fanout1139 (.A(_04860_),
    .X(net1139));
 sky130_fd_sc_hd__clkbuf_4 fanout1140 (.A(net1141),
    .X(net1140));
 sky130_fd_sc_hd__buf_2 fanout1141 (.A(net1144),
    .X(net1141));
 sky130_fd_sc_hd__buf_4 fanout1142 (.A(net1144),
    .X(net1142));
 sky130_fd_sc_hd__buf_2 fanout1143 (.A(net1144),
    .X(net1143));
 sky130_fd_sc_hd__clkbuf_8 fanout1144 (.A(_04783_),
    .X(net1144));
 sky130_fd_sc_hd__clkbuf_4 fanout1145 (.A(net1148),
    .X(net1145));
 sky130_fd_sc_hd__buf_2 fanout1146 (.A(net1148),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_4 fanout1147 (.A(net1148),
    .X(net1147));
 sky130_fd_sc_hd__clkbuf_4 fanout1148 (.A(_04703_),
    .X(net1148));
 sky130_fd_sc_hd__clkbuf_4 fanout1149 (.A(net1150),
    .X(net1149));
 sky130_fd_sc_hd__buf_2 fanout1150 (.A(net1151),
    .X(net1150));
 sky130_fd_sc_hd__clkbuf_4 fanout1151 (.A(net1152),
    .X(net1151));
 sky130_fd_sc_hd__buf_6 fanout1152 (.A(_04600_),
    .X(net1152));
 sky130_fd_sc_hd__buf_12 fanout1153 (.A(net1154),
    .X(net1153));
 sky130_fd_sc_hd__buf_8 fanout1154 (.A(_04545_),
    .X(net1154));
 sky130_fd_sc_hd__buf_12 fanout1155 (.A(net1156),
    .X(net1155));
 sky130_fd_sc_hd__buf_12 fanout1156 (.A(_04545_),
    .X(net1156));
 sky130_fd_sc_hd__buf_8 fanout1157 (.A(_04544_),
    .X(net1157));
 sky130_fd_sc_hd__buf_4 fanout1158 (.A(_04544_),
    .X(net1158));
 sky130_fd_sc_hd__clkbuf_16 fanout1159 (.A(_04544_),
    .X(net1159));
 sky130_fd_sc_hd__buf_4 fanout1160 (.A(_04544_),
    .X(net1160));
 sky130_fd_sc_hd__buf_4 fanout1161 (.A(net1162),
    .X(net1161));
 sky130_fd_sc_hd__buf_6 fanout1162 (.A(_04486_),
    .X(net1162));
 sky130_fd_sc_hd__buf_8 fanout1163 (.A(_04169_),
    .X(net1163));
 sky130_fd_sc_hd__buf_4 fanout1164 (.A(net1165),
    .X(net1164));
 sky130_fd_sc_hd__clkbuf_4 fanout1165 (.A(_09435_),
    .X(net1165));
 sky130_fd_sc_hd__buf_6 fanout1166 (.A(_09270_),
    .X(net1166));
 sky130_fd_sc_hd__buf_4 fanout1167 (.A(net1168),
    .X(net1167));
 sky130_fd_sc_hd__buf_4 fanout1168 (.A(_09238_),
    .X(net1168));
 sky130_fd_sc_hd__buf_6 fanout1169 (.A(_09237_),
    .X(net1169));
 sky130_fd_sc_hd__clkbuf_4 fanout1170 (.A(_09237_),
    .X(net1170));
 sky130_fd_sc_hd__buf_4 fanout1171 (.A(net1173),
    .X(net1171));
 sky130_fd_sc_hd__buf_6 fanout1172 (.A(net1173),
    .X(net1172));
 sky130_fd_sc_hd__buf_6 fanout1173 (.A(_09235_),
    .X(net1173));
 sky130_fd_sc_hd__buf_6 fanout1174 (.A(_09148_),
    .X(net1174));
 sky130_fd_sc_hd__buf_4 fanout1175 (.A(net1176),
    .X(net1175));
 sky130_fd_sc_hd__buf_4 fanout1176 (.A(_07471_),
    .X(net1176));
 sky130_fd_sc_hd__clkbuf_8 fanout1177 (.A(net1179),
    .X(net1177));
 sky130_fd_sc_hd__buf_2 fanout1178 (.A(net1179),
    .X(net1178));
 sky130_fd_sc_hd__buf_4 fanout1179 (.A(_07429_),
    .X(net1179));
 sky130_fd_sc_hd__buf_8 fanout1180 (.A(_07429_),
    .X(net1180));
 sky130_fd_sc_hd__clkbuf_4 fanout1181 (.A(_07429_),
    .X(net1181));
 sky130_fd_sc_hd__buf_4 fanout1182 (.A(net1183),
    .X(net1182));
 sky130_fd_sc_hd__clkbuf_16 fanout1183 (.A(_07399_),
    .X(net1183));
 sky130_fd_sc_hd__buf_6 fanout1184 (.A(net1186),
    .X(net1184));
 sky130_fd_sc_hd__buf_2 fanout1185 (.A(net1186),
    .X(net1185));
 sky130_fd_sc_hd__buf_6 fanout1186 (.A(_07398_),
    .X(net1186));
 sky130_fd_sc_hd__buf_6 fanout1187 (.A(_04599_),
    .X(net1187));
 sky130_fd_sc_hd__buf_6 fanout1188 (.A(net1191),
    .X(net1188));
 sky130_fd_sc_hd__buf_6 fanout1189 (.A(net1190),
    .X(net1189));
 sky130_fd_sc_hd__buf_4 fanout1190 (.A(net1191),
    .X(net1190));
 sky130_fd_sc_hd__buf_6 fanout1191 (.A(_04556_),
    .X(net1191));
 sky130_fd_sc_hd__buf_4 fanout1192 (.A(net1193),
    .X(net1192));
 sky130_fd_sc_hd__buf_4 fanout1193 (.A(net1194),
    .X(net1193));
 sky130_fd_sc_hd__clkbuf_8 fanout1194 (.A(_04485_),
    .X(net1194));
 sky130_fd_sc_hd__clkbuf_4 fanout1195 (.A(net1196),
    .X(net1195));
 sky130_fd_sc_hd__buf_2 fanout1196 (.A(net1198),
    .X(net1196));
 sky130_fd_sc_hd__buf_4 fanout1197 (.A(net1198),
    .X(net1197));
 sky130_fd_sc_hd__clkbuf_4 fanout1198 (.A(_03401_),
    .X(net1198));
 sky130_fd_sc_hd__buf_4 fanout1199 (.A(net1200),
    .X(net1199));
 sky130_fd_sc_hd__buf_4 fanout1200 (.A(net1202),
    .X(net1200));
 sky130_fd_sc_hd__buf_4 fanout1201 (.A(net1202),
    .X(net1201));
 sky130_fd_sc_hd__clkbuf_4 fanout1202 (.A(_03400_),
    .X(net1202));
 sky130_fd_sc_hd__buf_4 fanout1203 (.A(net1205),
    .X(net1203));
 sky130_fd_sc_hd__clkbuf_2 fanout1204 (.A(net1205),
    .X(net1204));
 sky130_fd_sc_hd__clkbuf_4 fanout1205 (.A(_03399_),
    .X(net1205));
 sky130_fd_sc_hd__buf_4 fanout1206 (.A(_03399_),
    .X(net1206));
 sky130_fd_sc_hd__buf_6 fanout1207 (.A(_02040_),
    .X(net1207));
 sky130_fd_sc_hd__buf_6 fanout1208 (.A(_09434_),
    .X(net1208));
 sky130_fd_sc_hd__buf_2 fanout1209 (.A(_09434_),
    .X(net1209));
 sky130_fd_sc_hd__buf_4 fanout1210 (.A(_09366_),
    .X(net1210));
 sky130_fd_sc_hd__buf_4 fanout1211 (.A(net1212),
    .X(net1211));
 sky130_fd_sc_hd__buf_6 fanout1212 (.A(_09365_),
    .X(net1212));
 sky130_fd_sc_hd__buf_4 fanout1213 (.A(net1214),
    .X(net1213));
 sky130_fd_sc_hd__buf_4 fanout1214 (.A(net1215),
    .X(net1214));
 sky130_fd_sc_hd__buf_8 fanout1215 (.A(_09147_),
    .X(net1215));
 sky130_fd_sc_hd__buf_6 fanout1216 (.A(net1217),
    .X(net1216));
 sky130_fd_sc_hd__buf_8 fanout1217 (.A(net1218),
    .X(net1217));
 sky130_fd_sc_hd__buf_8 fanout1218 (.A(_09064_),
    .X(net1218));
 sky130_fd_sc_hd__clkbuf_8 fanout1219 (.A(net1221),
    .X(net1219));
 sky130_fd_sc_hd__clkbuf_4 fanout1220 (.A(net1221),
    .X(net1220));
 sky130_fd_sc_hd__clkbuf_4 fanout1221 (.A(net1222),
    .X(net1221));
 sky130_fd_sc_hd__buf_4 fanout1222 (.A(_08005_),
    .X(net1222));
 sky130_fd_sc_hd__buf_6 fanout1223 (.A(net1225),
    .X(net1223));
 sky130_fd_sc_hd__buf_4 fanout1224 (.A(net1225),
    .X(net1224));
 sky130_fd_sc_hd__buf_4 fanout1225 (.A(_08005_),
    .X(net1225));
 sky130_fd_sc_hd__clkbuf_8 fanout1226 (.A(net1227),
    .X(net1226));
 sky130_fd_sc_hd__buf_4 fanout1227 (.A(net1228),
    .X(net1227));
 sky130_fd_sc_hd__buf_4 fanout1228 (.A(_07395_),
    .X(net1228));
 sky130_fd_sc_hd__buf_6 fanout1229 (.A(_07394_),
    .X(net1229));
 sky130_fd_sc_hd__clkbuf_4 fanout1230 (.A(_07394_),
    .X(net1230));
 sky130_fd_sc_hd__buf_4 fanout1231 (.A(net1232),
    .X(net1231));
 sky130_fd_sc_hd__buf_6 fanout1232 (.A(_07394_),
    .X(net1232));
 sky130_fd_sc_hd__buf_4 fanout1233 (.A(_04949_),
    .X(net1233));
 sky130_fd_sc_hd__buf_6 fanout1234 (.A(_04597_),
    .X(net1234));
 sky130_fd_sc_hd__buf_2 fanout1235 (.A(_04597_),
    .X(net1235));
 sky130_fd_sc_hd__buf_12 fanout1236 (.A(_04596_),
    .X(net1236));
 sky130_fd_sc_hd__buf_6 fanout1237 (.A(_04596_),
    .X(net1237));
 sky130_fd_sc_hd__buf_6 fanout1238 (.A(net1240),
    .X(net1238));
 sky130_fd_sc_hd__buf_6 fanout1239 (.A(net1240),
    .X(net1239));
 sky130_fd_sc_hd__buf_8 fanout1240 (.A(_04509_),
    .X(net1240));
 sky130_fd_sc_hd__buf_12 fanout1241 (.A(_04483_),
    .X(net1241));
 sky130_fd_sc_hd__buf_4 fanout1242 (.A(net1243),
    .X(net1242));
 sky130_fd_sc_hd__buf_6 fanout1243 (.A(_03471_),
    .X(net1243));
 sky130_fd_sc_hd__buf_6 fanout1244 (.A(net1245),
    .X(net1244));
 sky130_fd_sc_hd__buf_6 fanout1245 (.A(_03471_),
    .X(net1245));
 sky130_fd_sc_hd__buf_4 fanout1246 (.A(net1247),
    .X(net1246));
 sky130_fd_sc_hd__buf_6 fanout1247 (.A(_03470_),
    .X(net1247));
 sky130_fd_sc_hd__buf_6 fanout1248 (.A(net1249),
    .X(net1248));
 sky130_fd_sc_hd__buf_6 fanout1249 (.A(_03470_),
    .X(net1249));
 sky130_fd_sc_hd__buf_4 fanout1250 (.A(net1251),
    .X(net1250));
 sky130_fd_sc_hd__buf_6 fanout1251 (.A(_03469_),
    .X(net1251));
 sky130_fd_sc_hd__buf_6 fanout1252 (.A(net1253),
    .X(net1252));
 sky130_fd_sc_hd__buf_6 fanout1253 (.A(_03469_),
    .X(net1253));
 sky130_fd_sc_hd__buf_6 fanout1255 (.A(net1256),
    .X(net1255));
 sky130_fd_sc_hd__buf_8 fanout1256 (.A(_07842_),
    .X(net1256));
 sky130_fd_sc_hd__buf_4 fanout1257 (.A(net1258),
    .X(net1257));
 sky130_fd_sc_hd__buf_6 fanout1258 (.A(_07493_),
    .X(net1258));
 sky130_fd_sc_hd__buf_8 fanout1259 (.A(net1262),
    .X(net1259));
 sky130_fd_sc_hd__clkbuf_8 fanout1260 (.A(net1262),
    .X(net1260));
 sky130_fd_sc_hd__buf_2 fanout1261 (.A(net1262),
    .X(net1261));
 sky130_fd_sc_hd__buf_4 fanout1262 (.A(_07390_),
    .X(net1262));
 sky130_fd_sc_hd__clkbuf_16 fanout1263 (.A(net1264),
    .X(net1263));
 sky130_fd_sc_hd__buf_6 fanout1264 (.A(_04602_),
    .X(net1264));
 sky130_fd_sc_hd__buf_6 fanout1265 (.A(net1266),
    .X(net1265));
 sky130_fd_sc_hd__clkbuf_16 fanout1266 (.A(_04602_),
    .X(net1266));
 sky130_fd_sc_hd__buf_6 fanout1267 (.A(_04520_),
    .X(net1267));
 sky130_fd_sc_hd__buf_4 fanout1268 (.A(net1269),
    .X(net1268));
 sky130_fd_sc_hd__clkbuf_4 fanout1269 (.A(net1270),
    .X(net1269));
 sky130_fd_sc_hd__buf_6 fanout1270 (.A(_04520_),
    .X(net1270));
 sky130_fd_sc_hd__buf_6 fanout1271 (.A(_04507_),
    .X(net1271));
 sky130_fd_sc_hd__buf_4 fanout1272 (.A(_04479_),
    .X(net1272));
 sky130_fd_sc_hd__clkbuf_4 fanout1273 (.A(_04479_),
    .X(net1273));
 sky130_fd_sc_hd__buf_6 fanout1274 (.A(_04479_),
    .X(net1274));
 sky130_fd_sc_hd__buf_12 fanout1276 (.A(net1280),
    .X(net1276));
 sky130_fd_sc_hd__buf_4 fanout1277 (.A(net1280),
    .X(net1277));
 sky130_fd_sc_hd__buf_8 fanout1278 (.A(net1280),
    .X(net1278));
 sky130_fd_sc_hd__buf_6 fanout1279 (.A(net1280),
    .X(net1279));
 sky130_fd_sc_hd__buf_8 fanout1280 (.A(_04460_),
    .X(net1280));
 sky130_fd_sc_hd__buf_6 fanout1281 (.A(net1282),
    .X(net1281));
 sky130_fd_sc_hd__buf_6 fanout1282 (.A(_04460_),
    .X(net1282));
 sky130_fd_sc_hd__buf_4 fanout1283 (.A(_04460_),
    .X(net1283));
 sky130_fd_sc_hd__buf_4 fanout1284 (.A(_04460_),
    .X(net1284));
 sky130_fd_sc_hd__buf_6 fanout1285 (.A(net1286),
    .X(net1285));
 sky130_fd_sc_hd__clkbuf_16 fanout1286 (.A(_04459_),
    .X(net1286));
 sky130_fd_sc_hd__buf_8 fanout1287 (.A(net1289),
    .X(net1287));
 sky130_fd_sc_hd__buf_4 fanout1288 (.A(net1289),
    .X(net1288));
 sky130_fd_sc_hd__buf_6 fanout1289 (.A(_04459_),
    .X(net1289));
 sky130_fd_sc_hd__clkbuf_16 fanout1290 (.A(_04454_),
    .X(net1290));
 sky130_fd_sc_hd__buf_4 fanout1291 (.A(net1292),
    .X(net1291));
 sky130_fd_sc_hd__buf_2 fanout1292 (.A(net1293),
    .X(net1292));
 sky130_fd_sc_hd__clkbuf_2 fanout1293 (.A(net1297),
    .X(net1293));
 sky130_fd_sc_hd__buf_8 fanout1294 (.A(net1297),
    .X(net1294));
 sky130_fd_sc_hd__buf_6 fanout1295 (.A(net1296),
    .X(net1295));
 sky130_fd_sc_hd__buf_6 fanout1296 (.A(net1297),
    .X(net1296));
 sky130_fd_sc_hd__buf_6 fanout1297 (.A(_04453_),
    .X(net1297));
 sky130_fd_sc_hd__buf_6 fanout1298 (.A(net1299),
    .X(net1298));
 sky130_fd_sc_hd__buf_6 fanout1299 (.A(_08769_),
    .X(net1299));
 sky130_fd_sc_hd__clkbuf_16 fanout1300 (.A(net1301),
    .X(net1300));
 sky130_fd_sc_hd__buf_8 fanout1301 (.A(_08769_),
    .X(net1301));
 sky130_fd_sc_hd__buf_6 fanout1302 (.A(net1303),
    .X(net1302));
 sky130_fd_sc_hd__buf_6 fanout1303 (.A(net1305),
    .X(net1303));
 sky130_fd_sc_hd__buf_6 fanout1304 (.A(net1305),
    .X(net1304));
 sky130_fd_sc_hd__buf_6 fanout1305 (.A(_08372_),
    .X(net1305));
 sky130_fd_sc_hd__buf_6 fanout1306 (.A(_07836_),
    .X(net1306));
 sky130_fd_sc_hd__buf_4 fanout1307 (.A(_07836_),
    .X(net1307));
 sky130_fd_sc_hd__buf_4 fanout1308 (.A(net1312),
    .X(net1308));
 sky130_fd_sc_hd__clkbuf_4 fanout1309 (.A(net1312),
    .X(net1309));
 sky130_fd_sc_hd__clkbuf_8 fanout1310 (.A(net1311),
    .X(net1310));
 sky130_fd_sc_hd__buf_6 fanout1311 (.A(net1312),
    .X(net1311));
 sky130_fd_sc_hd__buf_4 fanout1312 (.A(_07387_),
    .X(net1312));
 sky130_fd_sc_hd__buf_6 fanout1313 (.A(_07386_),
    .X(net1313));
 sky130_fd_sc_hd__buf_6 fanout1314 (.A(net1315),
    .X(net1314));
 sky130_fd_sc_hd__clkbuf_4 fanout1315 (.A(_07386_),
    .X(net1315));
 sky130_fd_sc_hd__buf_6 fanout1316 (.A(_07383_),
    .X(net1316));
 sky130_fd_sc_hd__buf_6 fanout1317 (.A(net1319),
    .X(net1317));
 sky130_fd_sc_hd__buf_2 fanout1318 (.A(net1319),
    .X(net1318));
 sky130_fd_sc_hd__buf_6 fanout1319 (.A(_07380_),
    .X(net1319));
 sky130_fd_sc_hd__buf_6 fanout1320 (.A(net1322),
    .X(net1320));
 sky130_fd_sc_hd__clkbuf_4 fanout1321 (.A(net1322),
    .X(net1321));
 sky130_fd_sc_hd__buf_6 fanout1322 (.A(_07378_),
    .X(net1322));
 sky130_fd_sc_hd__buf_4 fanout1323 (.A(net1325),
    .X(net1323));
 sky130_fd_sc_hd__buf_4 fanout1324 (.A(net1325),
    .X(net1324));
 sky130_fd_sc_hd__buf_4 fanout1325 (.A(_07375_),
    .X(net1325));
 sky130_fd_sc_hd__buf_8 fanout1326 (.A(net1327),
    .X(net1326));
 sky130_fd_sc_hd__buf_8 fanout1327 (.A(_07372_),
    .X(net1327));
 sky130_fd_sc_hd__buf_6 fanout1328 (.A(net1330),
    .X(net1328));
 sky130_fd_sc_hd__buf_6 fanout1329 (.A(net1330),
    .X(net1329));
 sky130_fd_sc_hd__buf_6 fanout1330 (.A(_07371_),
    .X(net1330));
 sky130_fd_sc_hd__clkbuf_16 fanout1331 (.A(net1333),
    .X(net1331));
 sky130_fd_sc_hd__buf_6 fanout1332 (.A(net1333),
    .X(net1332));
 sky130_fd_sc_hd__buf_8 fanout1333 (.A(_04651_),
    .X(net1333));
 sky130_fd_sc_hd__buf_8 fanout1334 (.A(net1338),
    .X(net1334));
 sky130_fd_sc_hd__buf_8 fanout1335 (.A(net1337),
    .X(net1335));
 sky130_fd_sc_hd__clkbuf_4 fanout1336 (.A(net1337),
    .X(net1336));
 sky130_fd_sc_hd__buf_4 fanout1337 (.A(net1338),
    .X(net1337));
 sky130_fd_sc_hd__buf_8 fanout1338 (.A(_04651_),
    .X(net1338));
 sky130_fd_sc_hd__buf_6 fanout1339 (.A(_04601_),
    .X(net1339));
 sky130_fd_sc_hd__buf_2 fanout1340 (.A(_04601_),
    .X(net1340));
 sky130_fd_sc_hd__buf_6 fanout1341 (.A(_04601_),
    .X(net1341));
 sky130_fd_sc_hd__buf_6 fanout1342 (.A(net1343),
    .X(net1342));
 sky130_fd_sc_hd__clkbuf_4 fanout1343 (.A(net1344),
    .X(net1343));
 sky130_fd_sc_hd__buf_8 fanout1344 (.A(_03397_),
    .X(net1344));
 sky130_fd_sc_hd__buf_4 fanout1345 (.A(net1347),
    .X(net1345));
 sky130_fd_sc_hd__buf_2 fanout1346 (.A(net1347),
    .X(net1346));
 sky130_fd_sc_hd__buf_6 fanout1347 (.A(net1348),
    .X(net1347));
 sky130_fd_sc_hd__buf_6 fanout1348 (.A(net1349),
    .X(net1348));
 sky130_fd_sc_hd__buf_6 fanout1349 (.A(_03397_),
    .X(net1349));
 sky130_fd_sc_hd__buf_6 fanout1350 (.A(net1353),
    .X(net1350));
 sky130_fd_sc_hd__buf_2 fanout1351 (.A(net1353),
    .X(net1351));
 sky130_fd_sc_hd__buf_6 fanout1352 (.A(net1353),
    .X(net1352));
 sky130_fd_sc_hd__buf_6 fanout1353 (.A(_03373_),
    .X(net1353));
 sky130_fd_sc_hd__clkbuf_4 fanout1354 (.A(net1355),
    .X(net1354));
 sky130_fd_sc_hd__clkbuf_4 fanout1355 (.A(net1356),
    .X(net1355));
 sky130_fd_sc_hd__clkbuf_4 fanout1356 (.A(net1357),
    .X(net1356));
 sky130_fd_sc_hd__buf_2 fanout1357 (.A(net1358),
    .X(net1357));
 sky130_fd_sc_hd__clkbuf_8 fanout1358 (.A(_03047_),
    .X(net1358));
 sky130_fd_sc_hd__buf_4 fanout1359 (.A(net1361),
    .X(net1359));
 sky130_fd_sc_hd__buf_4 fanout1360 (.A(net1361),
    .X(net1360));
 sky130_fd_sc_hd__clkbuf_4 fanout1361 (.A(net1362),
    .X(net1361));
 sky130_fd_sc_hd__clkbuf_8 fanout1362 (.A(_08636_),
    .X(net1362));
 sky130_fd_sc_hd__clkbuf_4 fanout1363 (.A(net1364),
    .X(net1363));
 sky130_fd_sc_hd__buf_2 fanout1364 (.A(net1366),
    .X(net1364));
 sky130_fd_sc_hd__buf_4 fanout1365 (.A(net1366),
    .X(net1365));
 sky130_fd_sc_hd__buf_4 fanout1366 (.A(_08623_),
    .X(net1366));
 sky130_fd_sc_hd__buf_6 fanout1367 (.A(net1368),
    .X(net1367));
 sky130_fd_sc_hd__buf_8 fanout1368 (.A(_07833_),
    .X(net1368));
 sky130_fd_sc_hd__buf_8 fanout1369 (.A(net1371),
    .X(net1369));
 sky130_fd_sc_hd__buf_6 fanout1370 (.A(net1371),
    .X(net1370));
 sky130_fd_sc_hd__buf_6 fanout1371 (.A(_07833_),
    .X(net1371));
 sky130_fd_sc_hd__clkbuf_16 fanout1372 (.A(_07368_),
    .X(net1372));
 sky130_fd_sc_hd__buf_6 fanout1373 (.A(net1378),
    .X(net1373));
 sky130_fd_sc_hd__buf_6 fanout1374 (.A(net1375),
    .X(net1374));
 sky130_fd_sc_hd__clkbuf_8 fanout1375 (.A(net1378),
    .X(net1375));
 sky130_fd_sc_hd__buf_8 fanout1376 (.A(net1378),
    .X(net1376));
 sky130_fd_sc_hd__buf_8 fanout1377 (.A(net1378),
    .X(net1377));
 sky130_fd_sc_hd__buf_12 fanout1378 (.A(_04650_),
    .X(net1378));
 sky130_fd_sc_hd__buf_6 fanout1379 (.A(net1380),
    .X(net1379));
 sky130_fd_sc_hd__buf_6 fanout1380 (.A(net1387),
    .X(net1380));
 sky130_fd_sc_hd__buf_4 fanout1381 (.A(net1382),
    .X(net1381));
 sky130_fd_sc_hd__buf_6 fanout1382 (.A(net1387),
    .X(net1382));
 sky130_fd_sc_hd__buf_6 fanout1383 (.A(net1386),
    .X(net1383));
 sky130_fd_sc_hd__clkbuf_8 fanout1384 (.A(net1386),
    .X(net1384));
 sky130_fd_sc_hd__buf_6 fanout1385 (.A(net1386),
    .X(net1385));
 sky130_fd_sc_hd__buf_4 fanout1386 (.A(net1387),
    .X(net1386));
 sky130_fd_sc_hd__buf_4 fanout1387 (.A(_04649_),
    .X(net1387));
 sky130_fd_sc_hd__buf_6 fanout1388 (.A(net1389),
    .X(net1388));
 sky130_fd_sc_hd__buf_6 fanout1389 (.A(net1393),
    .X(net1389));
 sky130_fd_sc_hd__buf_6 fanout1390 (.A(net1391),
    .X(net1390));
 sky130_fd_sc_hd__buf_6 fanout1391 (.A(net1393),
    .X(net1391));
 sky130_fd_sc_hd__buf_6 fanout1392 (.A(net1393),
    .X(net1392));
 sky130_fd_sc_hd__buf_4 fanout1393 (.A(_04649_),
    .X(net1393));
 sky130_fd_sc_hd__clkbuf_8 fanout1394 (.A(net1398),
    .X(net1394));
 sky130_fd_sc_hd__clkbuf_8 fanout1395 (.A(net1398),
    .X(net1395));
 sky130_fd_sc_hd__buf_6 fanout1396 (.A(net1398),
    .X(net1396));
 sky130_fd_sc_hd__buf_4 fanout1397 (.A(net1398),
    .X(net1397));
 sky130_fd_sc_hd__buf_4 fanout1398 (.A(net1403),
    .X(net1398));
 sky130_fd_sc_hd__buf_6 fanout1399 (.A(net1400),
    .X(net1399));
 sky130_fd_sc_hd__buf_6 fanout1400 (.A(net1401),
    .X(net1400));
 sky130_fd_sc_hd__buf_8 fanout1401 (.A(net1403),
    .X(net1401));
 sky130_fd_sc_hd__buf_6 fanout1402 (.A(net1403),
    .X(net1402));
 sky130_fd_sc_hd__buf_6 fanout1403 (.A(_04649_),
    .X(net1403));
 sky130_fd_sc_hd__buf_6 fanout1404 (.A(net1407),
    .X(net1404));
 sky130_fd_sc_hd__buf_6 fanout1405 (.A(net1407),
    .X(net1405));
 sky130_fd_sc_hd__buf_6 fanout1406 (.A(net1407),
    .X(net1406));
 sky130_fd_sc_hd__buf_4 fanout1407 (.A(net1430),
    .X(net1407));
 sky130_fd_sc_hd__clkbuf_8 fanout1408 (.A(net1409),
    .X(net1408));
 sky130_fd_sc_hd__buf_6 fanout1409 (.A(net1412),
    .X(net1409));
 sky130_fd_sc_hd__buf_6 fanout1410 (.A(net1412),
    .X(net1410));
 sky130_fd_sc_hd__buf_2 fanout1411 (.A(net1412),
    .X(net1411));
 sky130_fd_sc_hd__buf_4 fanout1412 (.A(net1430),
    .X(net1412));
 sky130_fd_sc_hd__buf_6 fanout1413 (.A(net1414),
    .X(net1413));
 sky130_fd_sc_hd__buf_6 fanout1414 (.A(net1430),
    .X(net1414));
 sky130_fd_sc_hd__buf_6 fanout1415 (.A(net1422),
    .X(net1415));
 sky130_fd_sc_hd__buf_4 fanout1416 (.A(net1422),
    .X(net1416));
 sky130_fd_sc_hd__buf_6 fanout1417 (.A(net1422),
    .X(net1417));
 sky130_fd_sc_hd__clkbuf_8 fanout1418 (.A(net1422),
    .X(net1418));
 sky130_fd_sc_hd__buf_6 fanout1419 (.A(net1421),
    .X(net1419));
 sky130_fd_sc_hd__buf_6 fanout1420 (.A(net1421),
    .X(net1420));
 sky130_fd_sc_hd__buf_6 fanout1421 (.A(net1422),
    .X(net1421));
 sky130_fd_sc_hd__clkbuf_8 fanout1422 (.A(net1430),
    .X(net1422));
 sky130_fd_sc_hd__buf_6 fanout1423 (.A(net1425),
    .X(net1423));
 sky130_fd_sc_hd__clkbuf_4 fanout1424 (.A(net1425),
    .X(net1424));
 sky130_fd_sc_hd__buf_4 fanout1425 (.A(net1430),
    .X(net1425));
 sky130_fd_sc_hd__buf_6 fanout1426 (.A(net1429),
    .X(net1426));
 sky130_fd_sc_hd__clkbuf_4 fanout1427 (.A(net1429),
    .X(net1427));
 sky130_fd_sc_hd__buf_6 fanout1428 (.A(net1429),
    .X(net1428));
 sky130_fd_sc_hd__buf_4 fanout1429 (.A(net1430),
    .X(net1429));
 sky130_fd_sc_hd__buf_6 fanout1430 (.A(_04649_),
    .X(net1430));
 sky130_fd_sc_hd__buf_6 fanout1431 (.A(net1433),
    .X(net1431));
 sky130_fd_sc_hd__buf_6 fanout1432 (.A(net1433),
    .X(net1432));
 sky130_fd_sc_hd__buf_6 fanout1433 (.A(net1437),
    .X(net1433));
 sky130_fd_sc_hd__buf_6 fanout1434 (.A(net1437),
    .X(net1434));
 sky130_fd_sc_hd__buf_6 fanout1435 (.A(net1436),
    .X(net1435));
 sky130_fd_sc_hd__buf_8 fanout1436 (.A(net1437),
    .X(net1436));
 sky130_fd_sc_hd__buf_8 fanout1437 (.A(_04648_),
    .X(net1437));
 sky130_fd_sc_hd__buf_6 fanout1438 (.A(net1439),
    .X(net1438));
 sky130_fd_sc_hd__buf_6 fanout1439 (.A(_04648_),
    .X(net1439));
 sky130_fd_sc_hd__buf_12 fanout1440 (.A(net1441),
    .X(net1440));
 sky130_fd_sc_hd__buf_12 fanout1441 (.A(_04648_),
    .X(net1441));
 sky130_fd_sc_hd__buf_6 fanout1442 (.A(net1450),
    .X(net1442));
 sky130_fd_sc_hd__clkbuf_4 fanout1443 (.A(net1444),
    .X(net1443));
 sky130_fd_sc_hd__buf_8 fanout1444 (.A(net1450),
    .X(net1444));
 sky130_fd_sc_hd__buf_6 fanout1445 (.A(net1446),
    .X(net1445));
 sky130_fd_sc_hd__buf_6 fanout1446 (.A(net1450),
    .X(net1446));
 sky130_fd_sc_hd__buf_6 fanout1447 (.A(net1449),
    .X(net1447));
 sky130_fd_sc_hd__buf_6 fanout1448 (.A(net1449),
    .X(net1448));
 sky130_fd_sc_hd__buf_6 fanout1449 (.A(net1450),
    .X(net1449));
 sky130_fd_sc_hd__buf_6 fanout1450 (.A(_04647_),
    .X(net1450));
 sky130_fd_sc_hd__buf_6 fanout1451 (.A(net1453),
    .X(net1451));
 sky130_fd_sc_hd__buf_4 fanout1452 (.A(net1453),
    .X(net1452));
 sky130_fd_sc_hd__buf_6 fanout1453 (.A(net1454),
    .X(net1453));
 sky130_fd_sc_hd__clkbuf_4 fanout1454 (.A(_04647_),
    .X(net1454));
 sky130_fd_sc_hd__clkbuf_8 fanout1455 (.A(net1456),
    .X(net1455));
 sky130_fd_sc_hd__clkbuf_4 fanout1456 (.A(_04647_),
    .X(net1456));
 sky130_fd_sc_hd__buf_6 fanout1457 (.A(net1459),
    .X(net1457));
 sky130_fd_sc_hd__clkbuf_4 fanout1458 (.A(net1459),
    .X(net1458));
 sky130_fd_sc_hd__clkbuf_8 fanout1459 (.A(_04647_),
    .X(net1459));
 sky130_fd_sc_hd__buf_8 fanout1460 (.A(_04646_),
    .X(net1460));
 sky130_fd_sc_hd__buf_6 fanout1461 (.A(_04646_),
    .X(net1461));
 sky130_fd_sc_hd__buf_12 fanout1462 (.A(_04646_),
    .X(net1462));
 sky130_fd_sc_hd__buf_6 fanout1463 (.A(_04646_),
    .X(net1463));
 sky130_fd_sc_hd__clkbuf_16 fanout1464 (.A(_04645_),
    .X(net1464));
 sky130_fd_sc_hd__buf_8 fanout1465 (.A(net1477),
    .X(net1465));
 sky130_fd_sc_hd__buf_4 fanout1466 (.A(net1477),
    .X(net1466));
 sky130_fd_sc_hd__buf_6 fanout1467 (.A(net1468),
    .X(net1467));
 sky130_fd_sc_hd__buf_6 fanout1468 (.A(net1477),
    .X(net1468));
 sky130_fd_sc_hd__buf_8 fanout1469 (.A(net1471),
    .X(net1469));
 sky130_fd_sc_hd__buf_4 fanout1470 (.A(net1471),
    .X(net1470));
 sky130_fd_sc_hd__buf_4 fanout1471 (.A(net1477),
    .X(net1471));
 sky130_fd_sc_hd__clkbuf_16 fanout1472 (.A(net1473),
    .X(net1472));
 sky130_fd_sc_hd__buf_12 fanout1473 (.A(net1477),
    .X(net1473));
 sky130_fd_sc_hd__clkbuf_16 fanout1474 (.A(net1476),
    .X(net1474));
 sky130_fd_sc_hd__buf_8 fanout1475 (.A(net1476),
    .X(net1475));
 sky130_fd_sc_hd__buf_12 fanout1476 (.A(net1477),
    .X(net1476));
 sky130_fd_sc_hd__buf_12 fanout1477 (.A(_04644_),
    .X(net1477));
 sky130_fd_sc_hd__buf_6 fanout1478 (.A(net1479),
    .X(net1478));
 sky130_fd_sc_hd__clkbuf_8 fanout1479 (.A(net1480),
    .X(net1479));
 sky130_fd_sc_hd__clkbuf_16 fanout1480 (.A(net1483),
    .X(net1480));
 sky130_fd_sc_hd__buf_6 fanout1481 (.A(net1482),
    .X(net1481));
 sky130_fd_sc_hd__clkbuf_4 fanout1482 (.A(net1483),
    .X(net1482));
 sky130_fd_sc_hd__buf_12 fanout1483 (.A(_04643_),
    .X(net1483));
 sky130_fd_sc_hd__buf_8 fanout1484 (.A(net1486),
    .X(net1484));
 sky130_fd_sc_hd__buf_4 fanout1485 (.A(net1486),
    .X(net1485));
 sky130_fd_sc_hd__clkbuf_16 fanout1486 (.A(_04642_),
    .X(net1486));
 sky130_fd_sc_hd__buf_12 fanout1487 (.A(net1488),
    .X(net1487));
 sky130_fd_sc_hd__buf_12 fanout1488 (.A(_04642_),
    .X(net1488));
 sky130_fd_sc_hd__buf_6 fanout1489 (.A(net1490),
    .X(net1489));
 sky130_fd_sc_hd__buf_12 fanout1490 (.A(_04641_),
    .X(net1490));
 sky130_fd_sc_hd__clkbuf_16 fanout1491 (.A(net1492),
    .X(net1491));
 sky130_fd_sc_hd__buf_12 fanout1492 (.A(_04641_),
    .X(net1492));
 sky130_fd_sc_hd__buf_8 fanout1493 (.A(net1495),
    .X(net1493));
 sky130_fd_sc_hd__buf_6 fanout1494 (.A(net1495),
    .X(net1494));
 sky130_fd_sc_hd__clkbuf_8 fanout1495 (.A(net1503),
    .X(net1495));
 sky130_fd_sc_hd__buf_6 fanout1496 (.A(net1497),
    .X(net1496));
 sky130_fd_sc_hd__buf_6 fanout1497 (.A(net1503),
    .X(net1497));
 sky130_fd_sc_hd__buf_6 fanout1498 (.A(net1499),
    .X(net1498));
 sky130_fd_sc_hd__buf_6 fanout1499 (.A(net1503),
    .X(net1499));
 sky130_fd_sc_hd__buf_2 fanout1500 (.A(net1503),
    .X(net1500));
 sky130_fd_sc_hd__buf_8 fanout1501 (.A(net1502),
    .X(net1501));
 sky130_fd_sc_hd__buf_8 fanout1502 (.A(net1503),
    .X(net1502));
 sky130_fd_sc_hd__buf_8 fanout1503 (.A(_04541_),
    .X(net1503));
 sky130_fd_sc_hd__buf_6 fanout1504 (.A(net1505),
    .X(net1504));
 sky130_fd_sc_hd__clkbuf_8 fanout1505 (.A(net1508),
    .X(net1505));
 sky130_fd_sc_hd__buf_6 fanout1506 (.A(net1507),
    .X(net1506));
 sky130_fd_sc_hd__buf_6 fanout1507 (.A(net1508),
    .X(net1507));
 sky130_fd_sc_hd__clkbuf_4 fanout1508 (.A(net1534),
    .X(net1508));
 sky130_fd_sc_hd__buf_6 fanout1509 (.A(net1510),
    .X(net1509));
 sky130_fd_sc_hd__buf_6 fanout1510 (.A(net1513),
    .X(net1510));
 sky130_fd_sc_hd__clkbuf_8 fanout1511 (.A(net1512),
    .X(net1511));
 sky130_fd_sc_hd__buf_6 fanout1512 (.A(net1513),
    .X(net1512));
 sky130_fd_sc_hd__clkbuf_8 fanout1513 (.A(net1534),
    .X(net1513));
 sky130_fd_sc_hd__buf_6 fanout1514 (.A(net1515),
    .X(net1514));
 sky130_fd_sc_hd__buf_6 fanout1515 (.A(net1522),
    .X(net1515));
 sky130_fd_sc_hd__clkbuf_4 fanout1516 (.A(net1522),
    .X(net1516));
 sky130_fd_sc_hd__buf_6 fanout1517 (.A(net1518),
    .X(net1517));
 sky130_fd_sc_hd__buf_6 fanout1518 (.A(net1522),
    .X(net1518));
 sky130_fd_sc_hd__clkbuf_4 fanout1519 (.A(net1522),
    .X(net1519));
 sky130_fd_sc_hd__buf_6 fanout1520 (.A(net1521),
    .X(net1520));
 sky130_fd_sc_hd__buf_4 fanout1521 (.A(net1522),
    .X(net1521));
 sky130_fd_sc_hd__buf_4 fanout1522 (.A(net1534),
    .X(net1522));
 sky130_fd_sc_hd__buf_6 fanout1523 (.A(net1527),
    .X(net1523));
 sky130_fd_sc_hd__buf_6 fanout1524 (.A(net1527),
    .X(net1524));
 sky130_fd_sc_hd__buf_6 fanout1525 (.A(net1526),
    .X(net1525));
 sky130_fd_sc_hd__buf_6 fanout1526 (.A(net1527),
    .X(net1526));
 sky130_fd_sc_hd__buf_4 fanout1527 (.A(net1534),
    .X(net1527));
 sky130_fd_sc_hd__buf_6 fanout1528 (.A(net1529),
    .X(net1528));
 sky130_fd_sc_hd__buf_6 fanout1529 (.A(net1531),
    .X(net1529));
 sky130_fd_sc_hd__buf_6 fanout1530 (.A(net1531),
    .X(net1530));
 sky130_fd_sc_hd__buf_4 fanout1531 (.A(net1534),
    .X(net1531));
 sky130_fd_sc_hd__buf_6 fanout1532 (.A(net1533),
    .X(net1532));
 sky130_fd_sc_hd__buf_4 fanout1533 (.A(net1534),
    .X(net1533));
 sky130_fd_sc_hd__buf_6 fanout1534 (.A(net1566),
    .X(net1534));
 sky130_fd_sc_hd__buf_6 fanout1535 (.A(net1538),
    .X(net1535));
 sky130_fd_sc_hd__clkbuf_8 fanout1536 (.A(net1538),
    .X(net1536));
 sky130_fd_sc_hd__buf_6 fanout1537 (.A(net1538),
    .X(net1537));
 sky130_fd_sc_hd__buf_6 fanout1538 (.A(net1546),
    .X(net1538));
 sky130_fd_sc_hd__buf_6 fanout1539 (.A(net1543),
    .X(net1539));
 sky130_fd_sc_hd__buf_6 fanout1540 (.A(net1543),
    .X(net1540));
 sky130_fd_sc_hd__buf_6 fanout1541 (.A(net1543),
    .X(net1541));
 sky130_fd_sc_hd__clkbuf_4 fanout1542 (.A(net1543),
    .X(net1542));
 sky130_fd_sc_hd__clkbuf_8 fanout1543 (.A(net1546),
    .X(net1543));
 sky130_fd_sc_hd__buf_6 fanout1544 (.A(net1545),
    .X(net1544));
 sky130_fd_sc_hd__buf_4 fanout1545 (.A(net1546),
    .X(net1545));
 sky130_fd_sc_hd__buf_4 fanout1546 (.A(net1566),
    .X(net1546));
 sky130_fd_sc_hd__buf_6 fanout1547 (.A(net1556),
    .X(net1547));
 sky130_fd_sc_hd__buf_4 fanout1548 (.A(net1556),
    .X(net1548));
 sky130_fd_sc_hd__buf_6 fanout1549 (.A(net1556),
    .X(net1549));
 sky130_fd_sc_hd__buf_4 fanout1550 (.A(net1556),
    .X(net1550));
 sky130_fd_sc_hd__buf_6 fanout1551 (.A(net1552),
    .X(net1551));
 sky130_fd_sc_hd__clkbuf_4 fanout1552 (.A(net1556),
    .X(net1552));
 sky130_fd_sc_hd__buf_6 fanout1553 (.A(net1555),
    .X(net1553));
 sky130_fd_sc_hd__buf_6 fanout1554 (.A(net1555),
    .X(net1554));
 sky130_fd_sc_hd__clkbuf_4 fanout1555 (.A(net1556),
    .X(net1555));
 sky130_fd_sc_hd__clkbuf_8 fanout1556 (.A(net1566),
    .X(net1556));
 sky130_fd_sc_hd__clkbuf_8 fanout1557 (.A(net1559),
    .X(net1557));
 sky130_fd_sc_hd__clkbuf_8 fanout1558 (.A(net1559),
    .X(net1558));
 sky130_fd_sc_hd__buf_6 fanout1559 (.A(net1566),
    .X(net1559));
 sky130_fd_sc_hd__buf_6 fanout1560 (.A(net1565),
    .X(net1560));
 sky130_fd_sc_hd__clkbuf_8 fanout1561 (.A(net1565),
    .X(net1561));
 sky130_fd_sc_hd__buf_6 fanout1562 (.A(net1564),
    .X(net1562));
 sky130_fd_sc_hd__clkbuf_4 fanout1563 (.A(net1564),
    .X(net1563));
 sky130_fd_sc_hd__clkbuf_8 fanout1564 (.A(net1565),
    .X(net1564));
 sky130_fd_sc_hd__buf_4 fanout1565 (.A(net1566),
    .X(net1565));
 sky130_fd_sc_hd__buf_6 fanout1566 (.A(_04540_),
    .X(net1566));
 sky130_fd_sc_hd__buf_8 fanout1567 (.A(_04538_),
    .X(net1567));
 sky130_fd_sc_hd__buf_4 fanout1568 (.A(_04538_),
    .X(net1568));
 sky130_fd_sc_hd__clkbuf_16 fanout1569 (.A(_04538_),
    .X(net1569));
 sky130_fd_sc_hd__buf_4 fanout1570 (.A(_04538_),
    .X(net1570));
 sky130_fd_sc_hd__buf_8 fanout1571 (.A(_04537_),
    .X(net1571));
 sky130_fd_sc_hd__buf_4 fanout1572 (.A(_04537_),
    .X(net1572));
 sky130_fd_sc_hd__buf_8 fanout1573 (.A(_04537_),
    .X(net1573));
 sky130_fd_sc_hd__buf_6 fanout1574 (.A(_04537_),
    .X(net1574));
 sky130_fd_sc_hd__buf_6 fanout1575 (.A(net1576),
    .X(net1575));
 sky130_fd_sc_hd__buf_8 fanout1576 (.A(net1585),
    .X(net1576));
 sky130_fd_sc_hd__buf_6 fanout1577 (.A(net1585),
    .X(net1577));
 sky130_fd_sc_hd__clkbuf_4 fanout1578 (.A(net1585),
    .X(net1578));
 sky130_fd_sc_hd__buf_6 fanout1579 (.A(net1580),
    .X(net1579));
 sky130_fd_sc_hd__buf_6 fanout1580 (.A(net1584),
    .X(net1580));
 sky130_fd_sc_hd__buf_6 fanout1581 (.A(net1583),
    .X(net1581));
 sky130_fd_sc_hd__buf_4 fanout1582 (.A(net1583),
    .X(net1582));
 sky130_fd_sc_hd__clkbuf_8 fanout1583 (.A(net1584),
    .X(net1583));
 sky130_fd_sc_hd__clkbuf_8 fanout1584 (.A(net1585),
    .X(net1584));
 sky130_fd_sc_hd__buf_8 fanout1585 (.A(_04535_),
    .X(net1585));
 sky130_fd_sc_hd__buf_8 fanout1586 (.A(net1587),
    .X(net1586));
 sky130_fd_sc_hd__buf_8 fanout1587 (.A(net1596),
    .X(net1587));
 sky130_fd_sc_hd__buf_6 fanout1588 (.A(net1596),
    .X(net1588));
 sky130_fd_sc_hd__clkbuf_4 fanout1589 (.A(net1596),
    .X(net1589));
 sky130_fd_sc_hd__buf_6 fanout1590 (.A(net1591),
    .X(net1590));
 sky130_fd_sc_hd__buf_8 fanout1591 (.A(net1595),
    .X(net1591));
 sky130_fd_sc_hd__buf_6 fanout1592 (.A(net1594),
    .X(net1592));
 sky130_fd_sc_hd__clkbuf_4 fanout1593 (.A(net1594),
    .X(net1593));
 sky130_fd_sc_hd__clkbuf_8 fanout1594 (.A(net1595),
    .X(net1594));
 sky130_fd_sc_hd__buf_6 fanout1595 (.A(net1596),
    .X(net1595));
 sky130_fd_sc_hd__buf_6 fanout1596 (.A(_04534_),
    .X(net1596));
 sky130_fd_sc_hd__buf_6 fanout1597 (.A(net1598),
    .X(net1597));
 sky130_fd_sc_hd__buf_6 fanout1598 (.A(net1601),
    .X(net1598));
 sky130_fd_sc_hd__buf_6 fanout1599 (.A(net1600),
    .X(net1599));
 sky130_fd_sc_hd__buf_6 fanout1600 (.A(net1601),
    .X(net1600));
 sky130_fd_sc_hd__buf_4 fanout1601 (.A(_04531_),
    .X(net1601));
 sky130_fd_sc_hd__buf_6 fanout1602 (.A(net1603),
    .X(net1602));
 sky130_fd_sc_hd__buf_8 fanout1603 (.A(net1604),
    .X(net1603));
 sky130_fd_sc_hd__buf_4 fanout1604 (.A(_04531_),
    .X(net1604));
 sky130_fd_sc_hd__buf_8 fanout1605 (.A(net1606),
    .X(net1605));
 sky130_fd_sc_hd__buf_8 fanout1606 (.A(_04531_),
    .X(net1606));
 sky130_fd_sc_hd__buf_6 fanout1607 (.A(net1609),
    .X(net1607));
 sky130_fd_sc_hd__clkbuf_4 fanout1608 (.A(net1609),
    .X(net1608));
 sky130_fd_sc_hd__buf_6 fanout1609 (.A(net1610),
    .X(net1609));
 sky130_fd_sc_hd__buf_6 fanout1610 (.A(_04531_),
    .X(net1610));
 sky130_fd_sc_hd__buf_6 fanout1611 (.A(net1613),
    .X(net1611));
 sky130_fd_sc_hd__buf_6 fanout1612 (.A(net1613),
    .X(net1612));
 sky130_fd_sc_hd__buf_6 fanout1613 (.A(net1630),
    .X(net1613));
 sky130_fd_sc_hd__buf_6 fanout1614 (.A(net1616),
    .X(net1614));
 sky130_fd_sc_hd__buf_4 fanout1615 (.A(net1616),
    .X(net1615));
 sky130_fd_sc_hd__buf_4 fanout1616 (.A(net1630),
    .X(net1616));
 sky130_fd_sc_hd__buf_6 fanout1617 (.A(net1618),
    .X(net1617));
 sky130_fd_sc_hd__buf_8 fanout1618 (.A(net1619),
    .X(net1618));
 sky130_fd_sc_hd__buf_6 fanout1619 (.A(net1630),
    .X(net1619));
 sky130_fd_sc_hd__buf_8 fanout1620 (.A(net1622),
    .X(net1620));
 sky130_fd_sc_hd__buf_6 fanout1621 (.A(net1622),
    .X(net1621));
 sky130_fd_sc_hd__buf_6 fanout1622 (.A(net1623),
    .X(net1622));
 sky130_fd_sc_hd__buf_6 fanout1623 (.A(net1630),
    .X(net1623));
 sky130_fd_sc_hd__buf_6 fanout1624 (.A(net1626),
    .X(net1624));
 sky130_fd_sc_hd__clkbuf_4 fanout1625 (.A(net1626),
    .X(net1625));
 sky130_fd_sc_hd__buf_8 fanout1626 (.A(net1630),
    .X(net1626));
 sky130_fd_sc_hd__buf_6 fanout1627 (.A(net1630),
    .X(net1627));
 sky130_fd_sc_hd__buf_4 fanout1628 (.A(net1629),
    .X(net1628));
 sky130_fd_sc_hd__buf_6 fanout1629 (.A(net1630),
    .X(net1629));
 sky130_fd_sc_hd__buf_12 fanout1630 (.A(_04530_),
    .X(net1630));
 sky130_fd_sc_hd__buf_8 fanout1631 (.A(_04528_),
    .X(net1631));
 sky130_fd_sc_hd__buf_6 fanout1632 (.A(_04528_),
    .X(net1632));
 sky130_fd_sc_hd__buf_12 fanout1633 (.A(_04528_),
    .X(net1633));
 sky130_fd_sc_hd__buf_4 fanout1634 (.A(_04528_),
    .X(net1634));
 sky130_fd_sc_hd__buf_8 fanout1635 (.A(_04527_),
    .X(net1635));
 sky130_fd_sc_hd__buf_4 fanout1636 (.A(_04527_),
    .X(net1636));
 sky130_fd_sc_hd__buf_8 fanout1637 (.A(net1638),
    .X(net1637));
 sky130_fd_sc_hd__buf_12 fanout1638 (.A(_04527_),
    .X(net1638));
 sky130_fd_sc_hd__buf_4 fanout1639 (.A(net1640),
    .X(net1639));
 sky130_fd_sc_hd__clkbuf_4 fanout1640 (.A(net1641),
    .X(net1640));
 sky130_fd_sc_hd__clkbuf_8 fanout1641 (.A(_07834_),
    .X(net1641));
 sky130_fd_sc_hd__buf_6 fanout1642 (.A(net1643),
    .X(net1642));
 sky130_fd_sc_hd__buf_6 fanout1643 (.A(_07834_),
    .X(net1643));
 sky130_fd_sc_hd__buf_6 fanout1644 (.A(net1646),
    .X(net1644));
 sky130_fd_sc_hd__buf_6 fanout1645 (.A(net1646),
    .X(net1645));
 sky130_fd_sc_hd__buf_8 fanout1646 (.A(_07445_),
    .X(net1646));
 sky130_fd_sc_hd__buf_6 fanout1647 (.A(net1648),
    .X(net1647));
 sky130_fd_sc_hd__buf_4 fanout1648 (.A(_07444_),
    .X(net1648));
 sky130_fd_sc_hd__buf_8 fanout1649 (.A(_07444_),
    .X(net1649));
 sky130_fd_sc_hd__clkbuf_4 fanout1650 (.A(_07444_),
    .X(net1650));
 sky130_fd_sc_hd__buf_6 fanout1651 (.A(_04583_),
    .X(net1651));
 sky130_fd_sc_hd__buf_2 fanout1652 (.A(_04583_),
    .X(net1652));
 sky130_fd_sc_hd__buf_4 fanout1653 (.A(net1654),
    .X(net1653));
 sky130_fd_sc_hd__clkbuf_8 fanout1654 (.A(_04575_),
    .X(net1654));
 sky130_fd_sc_hd__buf_12 fanout1655 (.A(_04568_),
    .X(net1655));
 sky130_fd_sc_hd__buf_4 fanout1656 (.A(_04568_),
    .X(net1656));
 sky130_fd_sc_hd__buf_4 fanout1657 (.A(net1658),
    .X(net1657));
 sky130_fd_sc_hd__buf_8 fanout1658 (.A(net1659),
    .X(net1658));
 sky130_fd_sc_hd__buf_8 fanout1659 (.A(_04561_),
    .X(net1659));
 sky130_fd_sc_hd__buf_4 fanout1660 (.A(_04559_),
    .X(net1660));
 sky130_fd_sc_hd__buf_4 fanout1661 (.A(_04559_),
    .X(net1661));
 sky130_fd_sc_hd__clkbuf_16 fanout1662 (.A(net1666),
    .X(net1662));
 sky130_fd_sc_hd__buf_12 fanout1663 (.A(net1664),
    .X(net1663));
 sky130_fd_sc_hd__buf_6 fanout1664 (.A(net1665),
    .X(net1664));
 sky130_fd_sc_hd__buf_12 fanout1665 (.A(net1666),
    .X(net1665));
 sky130_fd_sc_hd__buf_12 fanout1666 (.A(_04446_),
    .X(net1666));
 sky130_fd_sc_hd__buf_12 fanout1667 (.A(net1668),
    .X(net1667));
 sky130_fd_sc_hd__buf_12 fanout1668 (.A(_04445_),
    .X(net1668));
 sky130_fd_sc_hd__buf_4 fanout1669 (.A(net1671),
    .X(net1669));
 sky130_fd_sc_hd__buf_4 fanout1670 (.A(net1671),
    .X(net1670));
 sky130_fd_sc_hd__clkbuf_4 fanout1671 (.A(net1672),
    .X(net1671));
 sky130_fd_sc_hd__clkbuf_8 fanout1672 (.A(_04431_),
    .X(net1672));
 sky130_fd_sc_hd__buf_8 fanout1673 (.A(net1674),
    .X(net1673));
 sky130_fd_sc_hd__buf_6 fanout1674 (.A(net1675),
    .X(net1674));
 sky130_fd_sc_hd__buf_8 fanout1675 (.A(net1676),
    .X(net1675));
 sky130_fd_sc_hd__buf_8 fanout1676 (.A(_04430_),
    .X(net1676));
 sky130_fd_sc_hd__buf_6 fanout1677 (.A(net1678),
    .X(net1677));
 sky130_fd_sc_hd__buf_6 fanout1678 (.A(net1683),
    .X(net1678));
 sky130_fd_sc_hd__buf_6 fanout1679 (.A(net1681),
    .X(net1679));
 sky130_fd_sc_hd__buf_4 fanout1680 (.A(net1681),
    .X(net1680));
 sky130_fd_sc_hd__buf_4 fanout1681 (.A(net1683),
    .X(net1681));
 sky130_fd_sc_hd__buf_6 fanout1682 (.A(net1683),
    .X(net1682));
 sky130_fd_sc_hd__clkbuf_8 fanout1683 (.A(net1703),
    .X(net1683));
 sky130_fd_sc_hd__buf_6 fanout1684 (.A(net1688),
    .X(net1684));
 sky130_fd_sc_hd__buf_4 fanout1685 (.A(net1688),
    .X(net1685));
 sky130_fd_sc_hd__buf_6 fanout1686 (.A(net1688),
    .X(net1686));
 sky130_fd_sc_hd__buf_4 fanout1687 (.A(net1688),
    .X(net1687));
 sky130_fd_sc_hd__buf_12 fanout1688 (.A(net1703),
    .X(net1688));
 sky130_fd_sc_hd__buf_4 fanout1689 (.A(net1691),
    .X(net1689));
 sky130_fd_sc_hd__buf_6 fanout1690 (.A(net1694),
    .X(net1690));
 sky130_fd_sc_hd__buf_2 fanout1691 (.A(net1694),
    .X(net1691));
 sky130_fd_sc_hd__clkbuf_8 fanout1692 (.A(net1693),
    .X(net1692));
 sky130_fd_sc_hd__buf_6 fanout1693 (.A(net1694),
    .X(net1693));
 sky130_fd_sc_hd__clkbuf_16 fanout1694 (.A(net1703),
    .X(net1694));
 sky130_fd_sc_hd__buf_6 fanout1695 (.A(net1702),
    .X(net1695));
 sky130_fd_sc_hd__buf_4 fanout1696 (.A(net1702),
    .X(net1696));
 sky130_fd_sc_hd__clkbuf_8 fanout1697 (.A(net1698),
    .X(net1697));
 sky130_fd_sc_hd__buf_6 fanout1698 (.A(net1702),
    .X(net1698));
 sky130_fd_sc_hd__clkbuf_8 fanout1699 (.A(net1700),
    .X(net1699));
 sky130_fd_sc_hd__buf_6 fanout1700 (.A(net1702),
    .X(net1700));
 sky130_fd_sc_hd__clkbuf_8 fanout1701 (.A(net1702),
    .X(net1701));
 sky130_fd_sc_hd__buf_8 fanout1702 (.A(net1703),
    .X(net1702));
 sky130_fd_sc_hd__buf_12 fanout1703 (.A(_04422_),
    .X(net1703));
 sky130_fd_sc_hd__buf_6 fanout1704 (.A(net1705),
    .X(net1704));
 sky130_fd_sc_hd__buf_6 fanout1705 (.A(net1714),
    .X(net1705));
 sky130_fd_sc_hd__buf_6 fanout1706 (.A(net1714),
    .X(net1706));
 sky130_fd_sc_hd__buf_6 fanout1707 (.A(net1708),
    .X(net1707));
 sky130_fd_sc_hd__buf_6 fanout1708 (.A(net1714),
    .X(net1708));
 sky130_fd_sc_hd__buf_6 fanout1709 (.A(net1710),
    .X(net1709));
 sky130_fd_sc_hd__buf_6 fanout1710 (.A(net1713),
    .X(net1710));
 sky130_fd_sc_hd__buf_6 fanout1711 (.A(net1713),
    .X(net1711));
 sky130_fd_sc_hd__buf_4 fanout1712 (.A(net1713),
    .X(net1712));
 sky130_fd_sc_hd__buf_4 fanout1713 (.A(net1714),
    .X(net1713));
 sky130_fd_sc_hd__clkbuf_16 fanout1714 (.A(_04421_),
    .X(net1714));
 sky130_fd_sc_hd__buf_12 fanout1715 (.A(_04420_),
    .X(net1715));
 sky130_fd_sc_hd__buf_12 fanout1716 (.A(net1718),
    .X(net1716));
 sky130_fd_sc_hd__buf_8 fanout1717 (.A(net1718),
    .X(net1717));
 sky130_fd_sc_hd__buf_8 fanout1718 (.A(_04419_),
    .X(net1718));
 sky130_fd_sc_hd__buf_6 fanout1719 (.A(net1720),
    .X(net1719));
 sky130_fd_sc_hd__buf_8 fanout1720 (.A(net1721),
    .X(net1720));
 sky130_fd_sc_hd__clkbuf_16 fanout1721 (.A(net1725),
    .X(net1721));
 sky130_fd_sc_hd__buf_6 fanout1722 (.A(net1724),
    .X(net1722));
 sky130_fd_sc_hd__buf_6 fanout1723 (.A(net1724),
    .X(net1723));
 sky130_fd_sc_hd__buf_6 fanout1724 (.A(net1725),
    .X(net1724));
 sky130_fd_sc_hd__clkbuf_16 fanout1725 (.A(_04418_),
    .X(net1725));
 sky130_fd_sc_hd__buf_6 fanout1726 (.A(net1727),
    .X(net1726));
 sky130_fd_sc_hd__buf_6 fanout1727 (.A(net1730),
    .X(net1727));
 sky130_fd_sc_hd__buf_6 fanout1728 (.A(net1729),
    .X(net1728));
 sky130_fd_sc_hd__buf_6 fanout1729 (.A(net1730),
    .X(net1729));
 sky130_fd_sc_hd__clkbuf_16 fanout1730 (.A(_04418_),
    .X(net1730));
 sky130_fd_sc_hd__buf_6 fanout1731 (.A(net1734),
    .X(net1731));
 sky130_fd_sc_hd__buf_6 fanout1732 (.A(net1734),
    .X(net1732));
 sky130_fd_sc_hd__buf_6 fanout1733 (.A(net1734),
    .X(net1733));
 sky130_fd_sc_hd__buf_6 fanout1734 (.A(_04418_),
    .X(net1734));
 sky130_fd_sc_hd__buf_6 fanout1735 (.A(net1736),
    .X(net1735));
 sky130_fd_sc_hd__buf_6 fanout1736 (.A(net1738),
    .X(net1736));
 sky130_fd_sc_hd__buf_8 fanout1737 (.A(net1738),
    .X(net1737));
 sky130_fd_sc_hd__buf_8 fanout1738 (.A(_04417_),
    .X(net1738));
 sky130_fd_sc_hd__buf_6 fanout1739 (.A(net1741),
    .X(net1739));
 sky130_fd_sc_hd__buf_6 fanout1740 (.A(net1741),
    .X(net1740));
 sky130_fd_sc_hd__buf_6 fanout1741 (.A(net1742),
    .X(net1741));
 sky130_fd_sc_hd__buf_8 fanout1742 (.A(net1743),
    .X(net1742));
 sky130_fd_sc_hd__buf_12 fanout1743 (.A(_04417_),
    .X(net1743));
 sky130_fd_sc_hd__buf_8 fanout1744 (.A(net1745),
    .X(net1744));
 sky130_fd_sc_hd__buf_8 fanout1745 (.A(_04416_),
    .X(net1745));
 sky130_fd_sc_hd__buf_12 fanout1746 (.A(_04416_),
    .X(net1746));
 sky130_fd_sc_hd__clkbuf_8 fanout1747 (.A(_04416_),
    .X(net1747));
 sky130_fd_sc_hd__buf_8 fanout1748 (.A(net1749),
    .X(net1748));
 sky130_fd_sc_hd__buf_6 fanout1749 (.A(_04415_),
    .X(net1749));
 sky130_fd_sc_hd__buf_6 fanout1750 (.A(net1751),
    .X(net1750));
 sky130_fd_sc_hd__buf_8 fanout1751 (.A(net1752),
    .X(net1751));
 sky130_fd_sc_hd__buf_12 fanout1752 (.A(_04415_),
    .X(net1752));
 sky130_fd_sc_hd__buf_8 fanout1753 (.A(_04413_),
    .X(net1753));
 sky130_fd_sc_hd__buf_6 fanout1754 (.A(net1756),
    .X(net1754));
 sky130_fd_sc_hd__clkbuf_4 fanout1755 (.A(net1756),
    .X(net1755));
 sky130_fd_sc_hd__buf_6 fanout1756 (.A(_04413_),
    .X(net1756));
 sky130_fd_sc_hd__buf_8 fanout1757 (.A(net1758),
    .X(net1757));
 sky130_fd_sc_hd__buf_8 fanout1758 (.A(net1759),
    .X(net1758));
 sky130_fd_sc_hd__buf_6 fanout1759 (.A(_04409_),
    .X(net1759));
 sky130_fd_sc_hd__buf_6 fanout1760 (.A(_04402_),
    .X(net1760));
 sky130_fd_sc_hd__buf_2 fanout1761 (.A(_04402_),
    .X(net1761));
 sky130_fd_sc_hd__buf_6 fanout1762 (.A(net1763),
    .X(net1762));
 sky130_fd_sc_hd__clkbuf_8 fanout1763 (.A(net1764),
    .X(net1763));
 sky130_fd_sc_hd__buf_4 fanout1764 (.A(net1765),
    .X(net1764));
 sky130_fd_sc_hd__buf_6 fanout1765 (.A(_04402_),
    .X(net1765));
 sky130_fd_sc_hd__buf_6 fanout1766 (.A(net1767),
    .X(net1766));
 sky130_fd_sc_hd__buf_6 fanout1767 (.A(net1770),
    .X(net1767));
 sky130_fd_sc_hd__buf_4 fanout1768 (.A(net1770),
    .X(net1768));
 sky130_fd_sc_hd__buf_2 fanout1769 (.A(net1770),
    .X(net1769));
 sky130_fd_sc_hd__buf_4 fanout1770 (.A(net1776),
    .X(net1770));
 sky130_fd_sc_hd__buf_4 fanout1771 (.A(net1772),
    .X(net1771));
 sky130_fd_sc_hd__clkbuf_4 fanout1772 (.A(net1773),
    .X(net1772));
 sky130_fd_sc_hd__clkbuf_4 fanout1773 (.A(net1776),
    .X(net1773));
 sky130_fd_sc_hd__clkbuf_8 fanout1774 (.A(net1776),
    .X(net1774));
 sky130_fd_sc_hd__buf_4 fanout1775 (.A(net1776),
    .X(net1775));
 sky130_fd_sc_hd__buf_12 fanout1776 (.A(net482),
    .X(net1776));
 sky130_fd_sc_hd__clkbuf_4 fanout1777 (.A(net1778),
    .X(net1777));
 sky130_fd_sc_hd__buf_4 fanout1778 (.A(\jtag.state[1] ),
    .X(net1778));
 sky130_fd_sc_hd__clkbuf_8 fanout1779 (.A(\jtag.state[0] ),
    .X(net1779));
 sky130_fd_sc_hd__buf_2 fanout1780 (.A(\jtag.state[0] ),
    .X(net1780));
 sky130_fd_sc_hd__buf_6 fanout1781 (.A(\jtag.tckRisingEdge ),
    .X(net1781));
 sky130_fd_sc_hd__clkbuf_4 fanout1782 (.A(\jtag.tckRisingEdge ),
    .X(net1782));
 sky130_fd_sc_hd__clkbuf_16 fanout1783 (.A(net1785),
    .X(net1783));
 sky130_fd_sc_hd__buf_12 fanout1784 (.A(net1785),
    .X(net1784));
 sky130_fd_sc_hd__buf_12 fanout1785 (.A(net1787),
    .X(net1785));
 sky130_fd_sc_hd__buf_12 fanout1786 (.A(net1787),
    .X(net1786));
 sky130_fd_sc_hd__buf_12 fanout1787 (.A(net1796),
    .X(net1787));
 sky130_fd_sc_hd__buf_12 fanout1788 (.A(net1796),
    .X(net1788));
 sky130_fd_sc_hd__buf_6 fanout1789 (.A(net1790),
    .X(net1789));
 sky130_fd_sc_hd__buf_6 fanout1790 (.A(net1791),
    .X(net1790));
 sky130_fd_sc_hd__clkbuf_16 fanout1791 (.A(net1795),
    .X(net1791));
 sky130_fd_sc_hd__buf_6 fanout1792 (.A(net1795),
    .X(net1792));
 sky130_fd_sc_hd__buf_2 fanout1793 (.A(net1794),
    .X(net1793));
 sky130_fd_sc_hd__buf_4 fanout1794 (.A(net1795),
    .X(net1794));
 sky130_fd_sc_hd__buf_6 fanout1795 (.A(net1796),
    .X(net1795));
 sky130_fd_sc_hd__buf_8 fanout1796 (.A(\core.management_run ),
    .X(net1796));
 sky130_fd_sc_hd__buf_4 fanout1797 (.A(net1798),
    .X(net1797));
 sky130_fd_sc_hd__clkbuf_4 fanout1798 (.A(\core.management_interruptEnable ),
    .X(net1798));
 sky130_fd_sc_hd__clkbuf_8 fanout1799 (.A(net1804),
    .X(net1799));
 sky130_fd_sc_hd__clkbuf_8 fanout1800 (.A(net1804),
    .X(net1800));
 sky130_fd_sc_hd__buf_4 fanout1801 (.A(net1804),
    .X(net1801));
 sky130_fd_sc_hd__buf_12 fanout1802 (.A(net1804),
    .X(net1802));
 sky130_fd_sc_hd__buf_6 fanout1803 (.A(net1804),
    .X(net1803));
 sky130_fd_sc_hd__buf_4 fanout1804 (.A(\localMemoryInterface.lastRWBankSelect ),
    .X(net1804));
 sky130_fd_sc_hd__buf_6 fanout1806 (.A(net1808),
    .X(net1806));
 sky130_fd_sc_hd__buf_8 fanout1807 (.A(net1808),
    .X(net1807));
 sky130_fd_sc_hd__buf_4 fanout1808 (.A(net1809),
    .X(net1808));
 sky130_fd_sc_hd__buf_2 fanout1809 (.A(\core.pipe1_resultRegister[1] ),
    .X(net1809));
 sky130_fd_sc_hd__buf_6 fanout1810 (.A(\core.pipe1_resultRegister[0] ),
    .X(net1810));
 sky130_fd_sc_hd__buf_8 fanout1811 (.A(\core.pipe1_resultRegister[0] ),
    .X(net1811));
 sky130_fd_sc_hd__buf_4 fanout1812 (.A(net1813),
    .X(net1812));
 sky130_fd_sc_hd__clkbuf_4 fanout1813 (.A(net1814),
    .X(net1813));
 sky130_fd_sc_hd__buf_4 fanout1814 (.A(\core.useCachedLoad ),
    .X(net1814));
 sky130_fd_sc_hd__buf_8 fanout1815 (.A(\core.pipe0_currentInstruction[31] ),
    .X(net1815));
 sky130_fd_sc_hd__buf_4 fanout1816 (.A(\core.pipe0_currentInstruction[31] ),
    .X(net1816));
 sky130_fd_sc_hd__buf_8 fanout1817 (.A(net1818),
    .X(net1817));
 sky130_fd_sc_hd__buf_6 fanout1818 (.A(\core.pipe0_currentInstruction[30] ),
    .X(net1818));
 sky130_fd_sc_hd__buf_12 fanout1819 (.A(\core.pipe0_currentInstruction[28] ),
    .X(net1819));
 sky130_fd_sc_hd__clkbuf_16 fanout1820 (.A(\core.pipe0_currentInstruction[27] ),
    .X(net1820));
 sky130_fd_sc_hd__clkbuf_16 fanout1821 (.A(\core.pipe0_currentInstruction[26] ),
    .X(net1821));
 sky130_fd_sc_hd__buf_12 fanout1822 (.A(\core.pipe0_currentInstruction[25] ),
    .X(net1822));
 sky130_fd_sc_hd__buf_6 fanout1823 (.A(net1824),
    .X(net1823));
 sky130_fd_sc_hd__buf_6 fanout1824 (.A(net1825),
    .X(net1824));
 sky130_fd_sc_hd__buf_12 fanout1825 (.A(net1830),
    .X(net1825));
 sky130_fd_sc_hd__buf_6 fanout1826 (.A(net1827),
    .X(net1826));
 sky130_fd_sc_hd__clkbuf_16 fanout1827 (.A(net1828),
    .X(net1827));
 sky130_fd_sc_hd__buf_12 fanout1828 (.A(net1829),
    .X(net1828));
 sky130_fd_sc_hd__buf_12 fanout1829 (.A(net1830),
    .X(net1829));
 sky130_fd_sc_hd__buf_12 fanout1830 (.A(\core.pipe0_currentInstruction[24] ),
    .X(net1830));
 sky130_fd_sc_hd__buf_12 fanout1831 (.A(\core.pipe0_currentInstruction[23] ),
    .X(net1831));
 sky130_fd_sc_hd__buf_6 fanout1832 (.A(net1833),
    .X(net1832));
 sky130_fd_sc_hd__buf_6 fanout1833 (.A(\core.pipe0_currentInstruction[22] ),
    .X(net1833));
 sky130_fd_sc_hd__buf_8 fanout1834 (.A(net1836),
    .X(net1834));
 sky130_fd_sc_hd__buf_4 fanout1835 (.A(net1836),
    .X(net1835));
 sky130_fd_sc_hd__buf_12 fanout1836 (.A(net1837),
    .X(net1836));
 sky130_fd_sc_hd__buf_8 fanout1837 (.A(\core.pipe0_currentInstruction[22] ),
    .X(net1837));
 sky130_fd_sc_hd__buf_4 fanout1838 (.A(net1839),
    .X(net1838));
 sky130_fd_sc_hd__buf_6 fanout1839 (.A(net1840),
    .X(net1839));
 sky130_fd_sc_hd__buf_8 fanout1840 (.A(net1843),
    .X(net1840));
 sky130_fd_sc_hd__buf_6 fanout1841 (.A(net1842),
    .X(net1841));
 sky130_fd_sc_hd__buf_6 fanout1842 (.A(net1843),
    .X(net1842));
 sky130_fd_sc_hd__buf_8 fanout1843 (.A(\core.pipe0_currentInstruction[21] ),
    .X(net1843));
 sky130_fd_sc_hd__clkbuf_8 fanout1844 (.A(net1849),
    .X(net1844));
 sky130_fd_sc_hd__buf_8 fanout1845 (.A(net1849),
    .X(net1845));
 sky130_fd_sc_hd__buf_8 fanout1846 (.A(net1848),
    .X(net1846));
 sky130_fd_sc_hd__buf_4 fanout1847 (.A(net1849),
    .X(net1847));
 sky130_fd_sc_hd__buf_12 fanout1848 (.A(net1849),
    .X(net1848));
 sky130_fd_sc_hd__buf_12 fanout1849 (.A(\core.pipe0_currentInstruction[21] ),
    .X(net1849));
 sky130_fd_sc_hd__buf_8 fanout1850 (.A(net1851),
    .X(net1850));
 sky130_fd_sc_hd__buf_12 fanout1851 (.A(net1852),
    .X(net1851));
 sky130_fd_sc_hd__buf_12 fanout1852 (.A(\core.pipe0_currentInstruction[20] ),
    .X(net1852));
 sky130_fd_sc_hd__buf_6 fanout1853 (.A(net1854),
    .X(net1853));
 sky130_fd_sc_hd__buf_6 fanout1854 (.A(net1855),
    .X(net1854));
 sky130_fd_sc_hd__clkbuf_16 fanout1855 (.A(net1861),
    .X(net1855));
 sky130_fd_sc_hd__clkbuf_16 fanout1856 (.A(net1861),
    .X(net1856));
 sky130_fd_sc_hd__buf_6 fanout1857 (.A(net1860),
    .X(net1857));
 sky130_fd_sc_hd__buf_6 fanout1858 (.A(net1859),
    .X(net1858));
 sky130_fd_sc_hd__buf_6 fanout1859 (.A(net1860),
    .X(net1859));
 sky130_fd_sc_hd__clkbuf_16 fanout1860 (.A(net1861),
    .X(net1860));
 sky130_fd_sc_hd__buf_12 fanout1861 (.A(\core.pipe0_currentInstruction[19] ),
    .X(net1861));
 sky130_fd_sc_hd__buf_6 fanout1862 (.A(net1863),
    .X(net1862));
 sky130_fd_sc_hd__buf_12 fanout1863 (.A(net1867),
    .X(net1863));
 sky130_fd_sc_hd__buf_6 fanout1864 (.A(net1865),
    .X(net1864));
 sky130_fd_sc_hd__buf_8 fanout1865 (.A(net1866),
    .X(net1865));
 sky130_fd_sc_hd__buf_12 fanout1866 (.A(net1867),
    .X(net1866));
 sky130_fd_sc_hd__buf_12 fanout1867 (.A(\core.pipe0_currentInstruction[17] ),
    .X(net1867));
 sky130_fd_sc_hd__buf_6 fanout1868 (.A(net1869),
    .X(net1868));
 sky130_fd_sc_hd__clkbuf_8 fanout1869 (.A(\core.pipe0_currentInstruction[16] ),
    .X(net1869));
 sky130_fd_sc_hd__buf_6 fanout1870 (.A(net1871),
    .X(net1870));
 sky130_fd_sc_hd__buf_6 fanout1871 (.A(\core.pipe0_currentInstruction[16] ),
    .X(net1871));
 sky130_fd_sc_hd__buf_8 fanout1872 (.A(net1873),
    .X(net1872));
 sky130_fd_sc_hd__buf_6 fanout1873 (.A(\core.pipe0_currentInstruction[16] ),
    .X(net1873));
 sky130_fd_sc_hd__buf_6 fanout1874 (.A(net1877),
    .X(net1874));
 sky130_fd_sc_hd__buf_6 fanout1875 (.A(net1876),
    .X(net1875));
 sky130_fd_sc_hd__buf_6 fanout1876 (.A(net1877),
    .X(net1876));
 sky130_fd_sc_hd__buf_6 fanout1877 (.A(\core.pipe0_currentInstruction[16] ),
    .X(net1877));
 sky130_fd_sc_hd__buf_8 fanout1878 (.A(net1879),
    .X(net1878));
 sky130_fd_sc_hd__buf_6 fanout1879 (.A(\core.pipe0_currentInstruction[14] ),
    .X(net1879));
 sky130_fd_sc_hd__buf_12 fanout1880 (.A(\core.pipe0_currentInstruction[13] ),
    .X(net1880));
 sky130_fd_sc_hd__buf_8 fanout1881 (.A(net1882),
    .X(net1881));
 sky130_fd_sc_hd__buf_8 fanout1882 (.A(\core.pipe0_currentInstruction[12] ),
    .X(net1882));
 sky130_fd_sc_hd__buf_6 fanout1883 (.A(net1884),
    .X(net1883));
 sky130_fd_sc_hd__buf_4 fanout1884 (.A(\core.pipe1_operation.currentPipeStall ),
    .X(net1884));
 sky130_fd_sc_hd__buf_8 fanout1885 (.A(\core.csr.currentInstruction[13] ),
    .X(net1885));
 sky130_fd_sc_hd__clkbuf_8 fanout1886 (.A(net1889),
    .X(net1886));
 sky130_fd_sc_hd__buf_2 fanout1887 (.A(net1889),
    .X(net1887));
 sky130_fd_sc_hd__buf_4 fanout1888 (.A(net1889),
    .X(net1888));
 sky130_fd_sc_hd__clkbuf_4 fanout1889 (.A(net1919),
    .X(net1889));
 sky130_fd_sc_hd__buf_4 fanout1890 (.A(net1919),
    .X(net1890));
 sky130_fd_sc_hd__buf_4 fanout1891 (.A(net1892),
    .X(net1891));
 sky130_fd_sc_hd__clkbuf_4 fanout1892 (.A(net1919),
    .X(net1892));
 sky130_fd_sc_hd__buf_4 fanout1893 (.A(net1894),
    .X(net1893));
 sky130_fd_sc_hd__buf_6 fanout1894 (.A(net1905),
    .X(net1894));
 sky130_fd_sc_hd__buf_4 fanout1895 (.A(net1896),
    .X(net1895));
 sky130_fd_sc_hd__clkbuf_4 fanout1896 (.A(net1898),
    .X(net1896));
 sky130_fd_sc_hd__clkbuf_4 fanout1897 (.A(net1898),
    .X(net1897));
 sky130_fd_sc_hd__clkbuf_2 fanout1898 (.A(net1905),
    .X(net1898));
 sky130_fd_sc_hd__clkbuf_8 fanout1899 (.A(net1905),
    .X(net1899));
 sky130_fd_sc_hd__clkbuf_4 fanout1900 (.A(net1905),
    .X(net1900));
 sky130_fd_sc_hd__clkbuf_4 fanout1901 (.A(net1902),
    .X(net1901));
 sky130_fd_sc_hd__clkbuf_4 fanout1902 (.A(net1904),
    .X(net1902));
 sky130_fd_sc_hd__clkbuf_4 fanout1903 (.A(net1904),
    .X(net1903));
 sky130_fd_sc_hd__buf_2 fanout1904 (.A(net1905),
    .X(net1904));
 sky130_fd_sc_hd__clkbuf_8 fanout1905 (.A(net1919),
    .X(net1905));
 sky130_fd_sc_hd__buf_4 fanout1906 (.A(net1908),
    .X(net1906));
 sky130_fd_sc_hd__clkbuf_2 fanout1907 (.A(net1908),
    .X(net1907));
 sky130_fd_sc_hd__buf_6 fanout1908 (.A(net1919),
    .X(net1908));
 sky130_fd_sc_hd__buf_4 fanout1909 (.A(net1918),
    .X(net1909));
 sky130_fd_sc_hd__clkbuf_4 fanout1910 (.A(net1918),
    .X(net1910));
 sky130_fd_sc_hd__buf_4 fanout1911 (.A(net1912),
    .X(net1911));
 sky130_fd_sc_hd__buf_4 fanout1912 (.A(net1918),
    .X(net1912));
 sky130_fd_sc_hd__buf_4 fanout1913 (.A(net1914),
    .X(net1913));
 sky130_fd_sc_hd__buf_2 fanout1914 (.A(net1915),
    .X(net1914));
 sky130_fd_sc_hd__clkbuf_8 fanout1915 (.A(net1918),
    .X(net1915));
 sky130_fd_sc_hd__buf_4 fanout1916 (.A(net1918),
    .X(net1916));
 sky130_fd_sc_hd__clkbuf_4 fanout1917 (.A(net1918),
    .X(net1917));
 sky130_fd_sc_hd__buf_6 fanout1918 (.A(net1919),
    .X(net1918));
 sky130_fd_sc_hd__buf_12 fanout1919 (.A(_04429_),
    .X(net1919));
 sky130_fd_sc_hd__buf_4 fanout1920 (.A(net1921),
    .X(net1920));
 sky130_fd_sc_hd__clkbuf_2 fanout1921 (.A(net1922),
    .X(net1921));
 sky130_fd_sc_hd__clkbuf_4 fanout1922 (.A(net1929),
    .X(net1922));
 sky130_fd_sc_hd__buf_4 fanout1923 (.A(net1924),
    .X(net1923));
 sky130_fd_sc_hd__buf_4 fanout1924 (.A(net1925),
    .X(net1924));
 sky130_fd_sc_hd__clkbuf_8 fanout1925 (.A(net1929),
    .X(net1925));
 sky130_fd_sc_hd__buf_4 fanout1926 (.A(net1928),
    .X(net1926));
 sky130_fd_sc_hd__buf_4 fanout1927 (.A(net1928),
    .X(net1927));
 sky130_fd_sc_hd__buf_4 fanout1928 (.A(net1929),
    .X(net1928));
 sky130_fd_sc_hd__buf_4 fanout1929 (.A(_04429_),
    .X(net1929));
 sky130_fd_sc_hd__buf_4 fanout1930 (.A(net1931),
    .X(net1930));
 sky130_fd_sc_hd__clkbuf_8 fanout1931 (.A(net1938),
    .X(net1931));
 sky130_fd_sc_hd__buf_4 fanout1932 (.A(net1933),
    .X(net1932));
 sky130_fd_sc_hd__clkbuf_4 fanout1933 (.A(net1938),
    .X(net1933));
 sky130_fd_sc_hd__buf_4 fanout1934 (.A(net1935),
    .X(net1934));
 sky130_fd_sc_hd__clkbuf_4 fanout1935 (.A(net1938),
    .X(net1935));
 sky130_fd_sc_hd__clkbuf_4 fanout1936 (.A(net1937),
    .X(net1936));
 sky130_fd_sc_hd__buf_2 fanout1937 (.A(net1938),
    .X(net1937));
 sky130_fd_sc_hd__buf_4 fanout1938 (.A(_04429_),
    .X(net1938));
 sky130_fd_sc_hd__buf_4 fanout1939 (.A(net1941),
    .X(net1939));
 sky130_fd_sc_hd__buf_4 fanout1940 (.A(net1946),
    .X(net1940));
 sky130_fd_sc_hd__buf_2 fanout1941 (.A(net1946),
    .X(net1941));
 sky130_fd_sc_hd__buf_4 fanout1942 (.A(net1943),
    .X(net1942));
 sky130_fd_sc_hd__buf_4 fanout1943 (.A(net1946),
    .X(net1943));
 sky130_fd_sc_hd__buf_4 fanout1944 (.A(net1945),
    .X(net1944));
 sky130_fd_sc_hd__buf_2 fanout1945 (.A(net1946),
    .X(net1945));
 sky130_fd_sc_hd__clkbuf_4 fanout1946 (.A(net1960),
    .X(net1946));
 sky130_fd_sc_hd__buf_4 fanout1947 (.A(net1948),
    .X(net1947));
 sky130_fd_sc_hd__clkbuf_2 fanout1948 (.A(net1960),
    .X(net1948));
 sky130_fd_sc_hd__buf_4 fanout1949 (.A(net1952),
    .X(net1949));
 sky130_fd_sc_hd__buf_4 fanout1950 (.A(net1951),
    .X(net1950));
 sky130_fd_sc_hd__clkbuf_4 fanout1951 (.A(net1952),
    .X(net1951));
 sky130_fd_sc_hd__buf_2 fanout1952 (.A(net1960),
    .X(net1952));
 sky130_fd_sc_hd__buf_4 fanout1953 (.A(net1954),
    .X(net1953));
 sky130_fd_sc_hd__clkbuf_4 fanout1954 (.A(net1956),
    .X(net1954));
 sky130_fd_sc_hd__clkbuf_4 fanout1955 (.A(net1956),
    .X(net1955));
 sky130_fd_sc_hd__buf_2 fanout1956 (.A(net1960),
    .X(net1956));
 sky130_fd_sc_hd__buf_4 fanout1957 (.A(net1958),
    .X(net1957));
 sky130_fd_sc_hd__buf_4 fanout1958 (.A(net1959),
    .X(net1958));
 sky130_fd_sc_hd__buf_4 fanout1959 (.A(net1960),
    .X(net1959));
 sky130_fd_sc_hd__buf_4 fanout1960 (.A(_04429_),
    .X(net1960));
 sky130_fd_sc_hd__buf_6 fanout1961 (.A(net1969),
    .X(net1961));
 sky130_fd_sc_hd__buf_4 fanout1962 (.A(net1964),
    .X(net1962));
 sky130_fd_sc_hd__buf_2 fanout1963 (.A(net1964),
    .X(net1963));
 sky130_fd_sc_hd__buf_4 fanout1964 (.A(net1968),
    .X(net1964));
 sky130_fd_sc_hd__buf_4 fanout1965 (.A(net1967),
    .X(net1965));
 sky130_fd_sc_hd__buf_4 fanout1966 (.A(net1967),
    .X(net1966));
 sky130_fd_sc_hd__buf_6 fanout1967 (.A(net1968),
    .X(net1967));
 sky130_fd_sc_hd__buf_4 fanout1968 (.A(net1969),
    .X(net1968));
 sky130_fd_sc_hd__buf_8 fanout1969 (.A(net1979),
    .X(net1969));
 sky130_fd_sc_hd__clkbuf_16 fanout1970 (.A(net1979),
    .X(net1970));
 sky130_fd_sc_hd__buf_4 fanout1971 (.A(net1974),
    .X(net1971));
 sky130_fd_sc_hd__buf_4 fanout1972 (.A(net1974),
    .X(net1972));
 sky130_fd_sc_hd__buf_2 fanout1973 (.A(net1974),
    .X(net1973));
 sky130_fd_sc_hd__buf_4 fanout1974 (.A(net1979),
    .X(net1974));
 sky130_fd_sc_hd__buf_6 fanout1975 (.A(net1978),
    .X(net1975));
 sky130_fd_sc_hd__buf_4 fanout1976 (.A(net1978),
    .X(net1976));
 sky130_fd_sc_hd__clkbuf_4 fanout1977 (.A(net1978),
    .X(net1977));
 sky130_fd_sc_hd__clkbuf_8 fanout1978 (.A(net1979),
    .X(net1978));
 sky130_fd_sc_hd__clkbuf_16 fanout1979 (.A(net284),
    .X(net1979));
 sky130_fd_sc_hd__buf_6 fanout1980 (.A(net1983),
    .X(net1980));
 sky130_fd_sc_hd__buf_6 fanout1981 (.A(net1983),
    .X(net1981));
 sky130_fd_sc_hd__clkbuf_4 fanout1982 (.A(net1983),
    .X(net1982));
 sky130_fd_sc_hd__clkbuf_8 fanout1983 (.A(net1989),
    .X(net1983));
 sky130_fd_sc_hd__buf_4 fanout1984 (.A(net1988),
    .X(net1984));
 sky130_fd_sc_hd__buf_4 fanout1985 (.A(net1986),
    .X(net1985));
 sky130_fd_sc_hd__buf_4 fanout1986 (.A(net1988),
    .X(net1986));
 sky130_fd_sc_hd__buf_2 fanout1987 (.A(net1988),
    .X(net1987));
 sky130_fd_sc_hd__buf_4 fanout1988 (.A(net1989),
    .X(net1988));
 sky130_fd_sc_hd__buf_8 fanout1989 (.A(net2002),
    .X(net1989));
 sky130_fd_sc_hd__buf_4 fanout1990 (.A(net1994),
    .X(net1990));
 sky130_fd_sc_hd__buf_4 fanout1991 (.A(net1994),
    .X(net1991));
 sky130_fd_sc_hd__buf_4 fanout1992 (.A(net1993),
    .X(net1992));
 sky130_fd_sc_hd__clkbuf_4 fanout1993 (.A(net1994),
    .X(net1993));
 sky130_fd_sc_hd__clkbuf_4 fanout1994 (.A(net2002),
    .X(net1994));
 sky130_fd_sc_hd__buf_4 fanout1995 (.A(net1996),
    .X(net1995));
 sky130_fd_sc_hd__clkbuf_8 fanout1996 (.A(net2002),
    .X(net1996));
 sky130_fd_sc_hd__buf_4 fanout1997 (.A(net1998),
    .X(net1997));
 sky130_fd_sc_hd__buf_4 fanout1998 (.A(net2002),
    .X(net1998));
 sky130_fd_sc_hd__buf_4 fanout1999 (.A(net2001),
    .X(net1999));
 sky130_fd_sc_hd__buf_2 fanout2000 (.A(net2001),
    .X(net2000));
 sky130_fd_sc_hd__buf_6 fanout2001 (.A(net2002),
    .X(net2001));
 sky130_fd_sc_hd__buf_8 fanout2002 (.A(net284),
    .X(net2002));
 sky130_fd_sc_hd__buf_4 fanout2003 (.A(net2005),
    .X(net2003));
 sky130_fd_sc_hd__buf_4 fanout2004 (.A(net2005),
    .X(net2004));
 sky130_fd_sc_hd__clkbuf_4 fanout2005 (.A(net2006),
    .X(net2005));
 sky130_fd_sc_hd__buf_4 fanout2006 (.A(net205),
    .X(net2006));
 sky130_fd_sc_hd__buf_12 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__buf_6 fanout489 (.A(_03614_),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_16 fanout490 (.A(net491),
    .X(net490));
 sky130_fd_sc_hd__buf_12 fanout491 (.A(_03614_),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_16 fanout492 (.A(_03612_),
    .X(net492));
 sky130_fd_sc_hd__buf_6 fanout493 (.A(_03612_),
    .X(net493));
 sky130_fd_sc_hd__buf_12 fanout494 (.A(_03612_),
    .X(net494));
 sky130_fd_sc_hd__buf_6 fanout495 (.A(_03612_),
    .X(net495));
 sky130_fd_sc_hd__buf_12 fanout496 (.A(_03610_),
    .X(net496));
 sky130_fd_sc_hd__buf_4 fanout497 (.A(_03610_),
    .X(net497));
 sky130_fd_sc_hd__buf_12 fanout498 (.A(_03610_),
    .X(net498));
 sky130_fd_sc_hd__buf_6 fanout499 (.A(_03610_),
    .X(net499));
 sky130_fd_sc_hd__buf_12 fanout500 (.A(_03608_),
    .X(net500));
 sky130_fd_sc_hd__buf_4 fanout501 (.A(_03608_),
    .X(net501));
 sky130_fd_sc_hd__buf_12 fanout502 (.A(_03608_),
    .X(net502));
 sky130_fd_sc_hd__buf_6 fanout503 (.A(_03608_),
    .X(net503));
 sky130_fd_sc_hd__buf_12 fanout504 (.A(_03606_),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_8 fanout505 (.A(_03606_),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_16 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_16 fanout507 (.A(_03606_),
    .X(net507));
 sky130_fd_sc_hd__buf_12 fanout508 (.A(_03604_),
    .X(net508));
 sky130_fd_sc_hd__buf_4 fanout509 (.A(_03604_),
    .X(net509));
 sky130_fd_sc_hd__buf_12 fanout510 (.A(_03604_),
    .X(net510));
 sky130_fd_sc_hd__buf_6 fanout511 (.A(_03604_),
    .X(net511));
 sky130_fd_sc_hd__buf_12 fanout512 (.A(_03602_),
    .X(net512));
 sky130_fd_sc_hd__buf_4 fanout513 (.A(_03602_),
    .X(net513));
 sky130_fd_sc_hd__buf_12 fanout514 (.A(_03602_),
    .X(net514));
 sky130_fd_sc_hd__buf_6 fanout515 (.A(_03602_),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_16 fanout516 (.A(_03599_),
    .X(net516));
 sky130_fd_sc_hd__buf_4 fanout517 (.A(_03599_),
    .X(net517));
 sky130_fd_sc_hd__buf_12 fanout518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__buf_12 fanout519 (.A(_03599_),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_16 fanout520 (.A(_03597_),
    .X(net520));
 sky130_fd_sc_hd__buf_6 fanout521 (.A(_03597_),
    .X(net521));
 sky130_fd_sc_hd__buf_12 fanout522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__buf_12 fanout523 (.A(_03597_),
    .X(net523));
 sky130_fd_sc_hd__clkbuf_16 fanout524 (.A(_03595_),
    .X(net524));
 sky130_fd_sc_hd__buf_6 fanout525 (.A(_03595_),
    .X(net525));
 sky130_fd_sc_hd__buf_12 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_12 fanout527 (.A(_03595_),
    .X(net527));
 sky130_fd_sc_hd__buf_12 fanout528 (.A(_03593_),
    .X(net528));
 sky130_fd_sc_hd__buf_4 fanout529 (.A(_03593_),
    .X(net529));
 sky130_fd_sc_hd__buf_12 fanout530 (.A(_03593_),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_8 fanout531 (.A(_03593_),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_16 fanout532 (.A(_03591_),
    .X(net532));
 sky130_fd_sc_hd__buf_4 fanout533 (.A(_03591_),
    .X(net533));
 sky130_fd_sc_hd__buf_12 fanout534 (.A(net535),
    .X(net534));
 sky130_fd_sc_hd__buf_12 fanout535 (.A(_03591_),
    .X(net535));
 sky130_fd_sc_hd__buf_8 fanout536 (.A(net539),
    .X(net536));
 sky130_fd_sc_hd__buf_12 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__buf_12 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_12 fanout539 (.A(_03387_),
    .X(net539));
 sky130_fd_sc_hd__buf_12 fanout540 (.A(net543),
    .X(net540));
 sky130_fd_sc_hd__buf_12 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__buf_12 fanout542 (.A(net543),
    .X(net542));
 sky130_fd_sc_hd__buf_12 fanout543 (.A(_03385_),
    .X(net543));
 sky130_fd_sc_hd__buf_12 fanout544 (.A(net547),
    .X(net544));
 sky130_fd_sc_hd__buf_12 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__buf_12 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__buf_12 fanout547 (.A(_03383_),
    .X(net547));
 sky130_fd_sc_hd__buf_12 fanout548 (.A(_03381_),
    .X(net548));
 sky130_fd_sc_hd__buf_6 fanout549 (.A(_03381_),
    .X(net549));
 sky130_fd_sc_hd__buf_12 fanout550 (.A(_03381_),
    .X(net550));
 sky130_fd_sc_hd__buf_6 fanout551 (.A(_03381_),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_16 fanout552 (.A(net553),
    .X(net552));
 sky130_fd_sc_hd__buf_6 fanout553 (.A(_03379_),
    .X(net553));
 sky130_fd_sc_hd__buf_12 fanout554 (.A(_03379_),
    .X(net554));
 sky130_fd_sc_hd__buf_6 fanout555 (.A(_03379_),
    .X(net555));
 sky130_fd_sc_hd__buf_12 fanout556 (.A(_03096_),
    .X(net556));
 sky130_fd_sc_hd__buf_4 fanout557 (.A(_03096_),
    .X(net557));
 sky130_fd_sc_hd__buf_12 fanout558 (.A(_03096_),
    .X(net558));
 sky130_fd_sc_hd__buf_6 fanout559 (.A(_03096_),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_16 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__buf_6 fanout561 (.A(_03094_),
    .X(net561));
 sky130_fd_sc_hd__buf_12 fanout562 (.A(_03094_),
    .X(net562));
 sky130_fd_sc_hd__buf_6 fanout563 (.A(_03094_),
    .X(net563));
 sky130_fd_sc_hd__buf_12 fanout564 (.A(_03092_),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_8 fanout565 (.A(_03092_),
    .X(net565));
 sky130_fd_sc_hd__buf_12 fanout566 (.A(net567),
    .X(net566));
 sky130_fd_sc_hd__buf_12 fanout567 (.A(_03092_),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_16 fanout568 (.A(_03044_),
    .X(net568));
 sky130_fd_sc_hd__buf_6 fanout569 (.A(_03044_),
    .X(net569));
 sky130_fd_sc_hd__buf_12 fanout570 (.A(_03044_),
    .X(net570));
 sky130_fd_sc_hd__buf_8 fanout571 (.A(_03044_),
    .X(net571));
 sky130_fd_sc_hd__buf_12 fanout572 (.A(_03042_),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_8 fanout573 (.A(_03042_),
    .X(net573));
 sky130_fd_sc_hd__buf_12 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__buf_12 fanout575 (.A(_03042_),
    .X(net575));
 sky130_fd_sc_hd__buf_8 fanout576 (.A(net579),
    .X(net576));
 sky130_fd_sc_hd__buf_12 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__buf_12 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__buf_12 fanout579 (.A(_02934_),
    .X(net579));
 sky130_fd_sc_hd__buf_12 fanout580 (.A(_02927_),
    .X(net580));
 sky130_fd_sc_hd__buf_4 fanout581 (.A(_02927_),
    .X(net581));
 sky130_fd_sc_hd__buf_12 fanout582 (.A(_02927_),
    .X(net582));
 sky130_fd_sc_hd__buf_6 fanout583 (.A(_02927_),
    .X(net583));
 sky130_fd_sc_hd__buf_4 fanout584 (.A(net585),
    .X(net584));
 sky130_fd_sc_hd__buf_4 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__buf_4 fanout586 (.A(_02860_),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_8 fanout587 (.A(_09111_),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_4 fanout588 (.A(_09111_),
    .X(net588));
 sky130_fd_sc_hd__buf_4 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__buf_4 fanout590 (.A(_09111_),
    .X(net590));
 sky130_fd_sc_hd__buf_12 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__buf_8 fanout592 (.A(_09109_),
    .X(net592));
 sky130_fd_sc_hd__buf_12 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__buf_12 fanout594 (.A(_09109_),
    .X(net594));
 sky130_fd_sc_hd__buf_12 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__buf_12 fanout596 (.A(_09107_),
    .X(net596));
 sky130_fd_sc_hd__buf_12 fanout597 (.A(net598),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_16 fanout598 (.A(_09107_),
    .X(net598));
 sky130_fd_sc_hd__buf_12 fanout599 (.A(_09104_),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_8 fanout600 (.A(_09104_),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_16 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_12 fanout602 (.A(_09104_),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_16 fanout603 (.A(_09102_),
    .X(net603));
 sky130_fd_sc_hd__buf_6 fanout604 (.A(_09102_),
    .X(net604));
 sky130_fd_sc_hd__buf_12 fanout605 (.A(_09102_),
    .X(net605));
 sky130_fd_sc_hd__buf_6 fanout606 (.A(_09102_),
    .X(net606));
 sky130_fd_sc_hd__buf_12 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__buf_6 fanout608 (.A(_09100_),
    .X(net608));
 sky130_fd_sc_hd__buf_12 fanout609 (.A(net610),
    .X(net609));
 sky130_fd_sc_hd__buf_12 fanout610 (.A(_09100_),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_16 fanout611 (.A(_09096_),
    .X(net611));
 sky130_fd_sc_hd__buf_6 fanout612 (.A(_09096_),
    .X(net612));
 sky130_fd_sc_hd__buf_12 fanout613 (.A(_09096_),
    .X(net613));
 sky130_fd_sc_hd__buf_8 fanout614 (.A(_09096_),
    .X(net614));
 sky130_fd_sc_hd__buf_12 fanout615 (.A(_09088_),
    .X(net615));
 sky130_fd_sc_hd__buf_6 fanout616 (.A(_09088_),
    .X(net616));
 sky130_fd_sc_hd__buf_12 fanout617 (.A(_09088_),
    .X(net617));
 sky130_fd_sc_hd__buf_6 fanout618 (.A(_09088_),
    .X(net618));
 sky130_fd_sc_hd__buf_6 fanout619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_8 fanout620 (.A(net622),
    .X(net620));
 sky130_fd_sc_hd__buf_6 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__buf_6 fanout622 (.A(_08768_),
    .X(net622));
 sky130_fd_sc_hd__buf_6 fanout623 (.A(_08653_),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_8 fanout624 (.A(_08653_),
    .X(net624));
 sky130_fd_sc_hd__buf_4 fanout625 (.A(net627),
    .X(net625));
 sky130_fd_sc_hd__buf_2 fanout626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_8 fanout627 (.A(_08652_),
    .X(net627));
 sky130_fd_sc_hd__buf_6 fanout628 (.A(_08652_),
    .X(net628));
 sky130_fd_sc_hd__buf_4 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_4 fanout630 (.A(net631),
    .X(net630));
 sky130_fd_sc_hd__buf_4 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__buf_6 fanout632 (.A(_08646_),
    .X(net632));
 sky130_fd_sc_hd__buf_12 fanout633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_16 fanout634 (.A(_03098_),
    .X(net634));
 sky130_fd_sc_hd__buf_4 fanout635 (.A(net636),
    .X(net635));
 sky130_fd_sc_hd__buf_4 fanout636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__buf_12 fanout637 (.A(_03098_),
    .X(net637));
 sky130_fd_sc_hd__buf_4 fanout638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_8 fanout639 (.A(_03098_),
    .X(net639));
 sky130_fd_sc_hd__buf_8 fanout640 (.A(net645),
    .X(net640));
 sky130_fd_sc_hd__buf_4 fanout641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__buf_4 fanout642 (.A(net645),
    .X(net642));
 sky130_fd_sc_hd__buf_4 fanout643 (.A(net645),
    .X(net643));
 sky130_fd_sc_hd__buf_2 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_8 fanout645 (.A(_02893_),
    .X(net645));
 sky130_fd_sc_hd__buf_6 fanout646 (.A(_02859_),
    .X(net646));
 sky130_fd_sc_hd__buf_4 fanout647 (.A(net650),
    .X(net647));
 sky130_fd_sc_hd__buf_4 fanout648 (.A(net650),
    .X(net648));
 sky130_fd_sc_hd__buf_2 fanout649 (.A(net650),
    .X(net649));
 sky130_fd_sc_hd__buf_2 fanout650 (.A(_02859_),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 fanout651 (.A(net654),
    .X(net651));
 sky130_fd_sc_hd__buf_4 fanout652 (.A(net654),
    .X(net652));
 sky130_fd_sc_hd__buf_4 fanout653 (.A(net654),
    .X(net653));
 sky130_fd_sc_hd__buf_4 fanout654 (.A(_09150_),
    .X(net654));
 sky130_fd_sc_hd__buf_4 fanout655 (.A(net656),
    .X(net655));
 sky130_fd_sc_hd__buf_4 fanout656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__buf_8 fanout657 (.A(_09150_),
    .X(net657));
 sky130_fd_sc_hd__buf_4 fanout658 (.A(_09110_),
    .X(net658));
 sky130_fd_sc_hd__buf_2 fanout659 (.A(_09110_),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_4 fanout660 (.A(net661),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_4 fanout661 (.A(_09110_),
    .X(net661));
 sky130_fd_sc_hd__buf_4 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__buf_4 fanout663 (.A(_08767_),
    .X(net663));
 sky130_fd_sc_hd__buf_6 fanout664 (.A(_08767_),
    .X(net664));
 sky130_fd_sc_hd__buf_2 fanout665 (.A(_08767_),
    .X(net665));
 sky130_fd_sc_hd__buf_4 fanout666 (.A(net668),
    .X(net666));
 sky130_fd_sc_hd__buf_2 fanout667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__buf_6 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__buf_8 fanout669 (.A(_08729_),
    .X(net669));
 sky130_fd_sc_hd__buf_6 fanout670 (.A(net674),
    .X(net670));
 sky130_fd_sc_hd__buf_4 fanout671 (.A(net672),
    .X(net671));
 sky130_fd_sc_hd__buf_4 fanout672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__buf_4 fanout673 (.A(net674),
    .X(net673));
 sky130_fd_sc_hd__buf_6 fanout674 (.A(_08651_),
    .X(net674));
 sky130_fd_sc_hd__clkbuf_4 fanout675 (.A(net677),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_2 fanout676 (.A(net677),
    .X(net676));
 sky130_fd_sc_hd__buf_6 fanout677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__buf_6 fanout678 (.A(_08645_),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_4 fanout679 (.A(net681),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_2 fanout680 (.A(net681),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_4 fanout681 (.A(net685),
    .X(net681));
 sky130_fd_sc_hd__buf_4 fanout682 (.A(net684),
    .X(net682));
 sky130_fd_sc_hd__buf_4 fanout683 (.A(net684),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_4 fanout684 (.A(net685),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_4 fanout685 (.A(_08645_),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_8 fanout686 (.A(net688),
    .X(net686));
 sky130_fd_sc_hd__buf_4 fanout687 (.A(net688),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_4 fanout688 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__buf_4 fanout689 (.A(_08645_),
    .X(net689));
 sky130_fd_sc_hd__buf_8 fanout690 (.A(net691),
    .X(net690));
 sky130_fd_sc_hd__buf_6 fanout691 (.A(net693),
    .X(net691));
 sky130_fd_sc_hd__buf_4 fanout692 (.A(net693),
    .X(net692));
 sky130_fd_sc_hd__buf_6 fanout693 (.A(_08619_),
    .X(net693));
 sky130_fd_sc_hd__buf_4 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__buf_4 fanout695 (.A(net696),
    .X(net695));
 sky130_fd_sc_hd__buf_6 fanout696 (.A(_08644_),
    .X(net696));
 sky130_fd_sc_hd__buf_6 fanout697 (.A(_08644_),
    .X(net697));
 sky130_fd_sc_hd__buf_4 fanout698 (.A(net700),
    .X(net698));
 sky130_fd_sc_hd__buf_2 fanout699 (.A(net700),
    .X(net699));
 sky130_fd_sc_hd__buf_4 fanout700 (.A(_08638_),
    .X(net700));
 sky130_fd_sc_hd__buf_6 fanout701 (.A(_08638_),
    .X(net701));
 sky130_fd_sc_hd__buf_8 fanout702 (.A(_08378_),
    .X(net702));
 sky130_fd_sc_hd__buf_4 fanout703 (.A(net704),
    .X(net703));
 sky130_fd_sc_hd__buf_4 fanout704 (.A(net705),
    .X(net704));
 sky130_fd_sc_hd__buf_6 fanout705 (.A(net706),
    .X(net705));
 sky130_fd_sc_hd__buf_4 fanout706 (.A(_03049_),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_4 fanout707 (.A(net708),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_2 fanout708 (.A(net710),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_4 fanout709 (.A(net710),
    .X(net709));
 sky130_fd_sc_hd__buf_2 fanout710 (.A(net711),
    .X(net710));
 sky130_fd_sc_hd__buf_4 fanout711 (.A(net713),
    .X(net711));
 sky130_fd_sc_hd__buf_12 fanout712 (.A(net713),
    .X(net712));
 sky130_fd_sc_hd__buf_12 fanout713 (.A(_08369_),
    .X(net713));
 sky130_fd_sc_hd__buf_4 fanout714 (.A(net715),
    .X(net714));
 sky130_fd_sc_hd__buf_4 fanout715 (.A(net716),
    .X(net715));
 sky130_fd_sc_hd__buf_6 fanout716 (.A(net717),
    .X(net716));
 sky130_fd_sc_hd__buf_4 fanout717 (.A(_03050_),
    .X(net717));
 sky130_fd_sc_hd__buf_6 fanout718 (.A(net722),
    .X(net718));
 sky130_fd_sc_hd__buf_4 fanout719 (.A(net720),
    .X(net719));
 sky130_fd_sc_hd__buf_6 fanout720 (.A(net722),
    .X(net720));
 sky130_fd_sc_hd__buf_2 fanout721 (.A(net722),
    .X(net721));
 sky130_fd_sc_hd__buf_8 fanout722 (.A(_08380_),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_16 fanout723 (.A(_08380_),
    .X(net723));
 sky130_fd_sc_hd__buf_8 fanout724 (.A(_08346_),
    .X(net724));
 sky130_fd_sc_hd__buf_6 fanout725 (.A(_08152_),
    .X(net725));
 sky130_fd_sc_hd__buf_4 fanout726 (.A(net727),
    .X(net726));
 sky130_fd_sc_hd__buf_4 fanout727 (.A(_00577_),
    .X(net727));
 sky130_fd_sc_hd__buf_6 fanout728 (.A(_00577_),
    .X(net728));
 sky130_fd_sc_hd__buf_8 fanout729 (.A(_00577_),
    .X(net729));
 sky130_fd_sc_hd__buf_8 fanout730 (.A(_04357_),
    .X(net730));
 sky130_fd_sc_hd__buf_4 fanout731 (.A(_04357_),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_8 fanout732 (.A(net733),
    .X(net732));
 sky130_fd_sc_hd__buf_6 fanout733 (.A(net735),
    .X(net733));
 sky130_fd_sc_hd__buf_6 fanout734 (.A(net735),
    .X(net734));
 sky130_fd_sc_hd__buf_6 fanout735 (.A(_04355_),
    .X(net735));
 sky130_fd_sc_hd__buf_6 fanout736 (.A(_04354_),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_4 fanout737 (.A(_04354_),
    .X(net737));
 sky130_fd_sc_hd__buf_4 fanout738 (.A(net739),
    .X(net738));
 sky130_fd_sc_hd__buf_4 fanout739 (.A(net741),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_8 fanout740 (.A(net741),
    .X(net740));
 sky130_fd_sc_hd__buf_4 fanout741 (.A(_08766_),
    .X(net741));
 sky130_fd_sc_hd__buf_6 fanout742 (.A(_04373_),
    .X(net742));
 sky130_fd_sc_hd__buf_6 fanout743 (.A(net746),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_4 fanout744 (.A(net746),
    .X(net744));
 sky130_fd_sc_hd__buf_6 fanout745 (.A(net746),
    .X(net745));
 sky130_fd_sc_hd__buf_6 fanout746 (.A(_04171_),
    .X(net746));
 sky130_fd_sc_hd__buf_4 fanout747 (.A(net749),
    .X(net747));
 sky130_fd_sc_hd__buf_4 fanout748 (.A(net749),
    .X(net748));
 sky130_fd_sc_hd__buf_6 fanout749 (.A(_03971_),
    .X(net749));
 sky130_fd_sc_hd__buf_4 fanout750 (.A(_03960_),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_4 fanout751 (.A(_03960_),
    .X(net751));
 sky130_fd_sc_hd__buf_6 fanout752 (.A(_03960_),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_4 fanout753 (.A(_03960_),
    .X(net753));
 sky130_fd_sc_hd__buf_4 fanout754 (.A(net755),
    .X(net754));
 sky130_fd_sc_hd__buf_6 fanout755 (.A(net757),
    .X(net755));
 sky130_fd_sc_hd__buf_4 fanout756 (.A(net757),
    .X(net756));
 sky130_fd_sc_hd__buf_4 fanout757 (.A(_04173_),
    .X(net757));
 sky130_fd_sc_hd__buf_4 fanout758 (.A(net760),
    .X(net758));
 sky130_fd_sc_hd__buf_6 fanout759 (.A(net760),
    .X(net759));
 sky130_fd_sc_hd__buf_6 fanout760 (.A(_04173_),
    .X(net760));
 sky130_fd_sc_hd__buf_6 fanout761 (.A(net762),
    .X(net761));
 sky130_fd_sc_hd__buf_4 fanout762 (.A(_04035_),
    .X(net762));
 sky130_fd_sc_hd__buf_6 fanout763 (.A(_04035_),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_4 fanout764 (.A(_04035_),
    .X(net764));
 sky130_fd_sc_hd__buf_8 fanout765 (.A(_08094_),
    .X(net765));
 sky130_fd_sc_hd__buf_6 fanout766 (.A(net768),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_16 fanout767 (.A(net768),
    .X(net767));
 sky130_fd_sc_hd__buf_6 fanout768 (.A(_04444_),
    .X(net768));
 sky130_fd_sc_hd__buf_4 fanout769 (.A(net770),
    .X(net769));
 sky130_fd_sc_hd__buf_6 fanout770 (.A(net776),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_8 fanout771 (.A(net773),
    .X(net771));
 sky130_fd_sc_hd__buf_2 fanout772 (.A(net773),
    .X(net772));
 sky130_fd_sc_hd__buf_4 fanout773 (.A(net776),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_8 fanout774 (.A(net776),
    .X(net774));
 sky130_fd_sc_hd__buf_6 fanout775 (.A(net776),
    .X(net775));
 sky130_fd_sc_hd__buf_6 fanout776 (.A(\core.csr.inTrap ),
    .X(net776));
 sky130_fd_sc_hd__buf_4 fanout777 (.A(net779),
    .X(net777));
 sky130_fd_sc_hd__buf_4 fanout778 (.A(net779),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_4 fanout779 (.A(net784),
    .X(net779));
 sky130_fd_sc_hd__buf_4 fanout780 (.A(net782),
    .X(net780));
 sky130_fd_sc_hd__buf_4 fanout781 (.A(net782),
    .X(net781));
 sky130_fd_sc_hd__buf_4 fanout782 (.A(net784),
    .X(net782));
 sky130_fd_sc_hd__buf_8 fanout783 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__buf_4 fanout784 (.A(\core.csr.inTrap ),
    .X(net784));
 sky130_fd_sc_hd__buf_8 fanout785 (.A(net786),
    .X(net785));
 sky130_fd_sc_hd__buf_4 fanout786 (.A(_07506_),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_8 fanout787 (.A(_07438_),
    .X(net787));
 sky130_fd_sc_hd__buf_6 fanout788 (.A(_07438_),
    .X(net788));
 sky130_fd_sc_hd__buf_6 fanout789 (.A(_07532_),
    .X(net789));
 sky130_fd_sc_hd__buf_4 fanout790 (.A(net791),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_4 fanout791 (.A(_07531_),
    .X(net791));
 sky130_fd_sc_hd__buf_6 fanout792 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__buf_8 fanout793 (.A(_07401_),
    .X(net793));
 sky130_fd_sc_hd__buf_8 fanout794 (.A(net796),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_8 fanout795 (.A(net796),
    .X(net795));
 sky130_fd_sc_hd__buf_8 fanout796 (.A(_07401_),
    .X(net796));
 sky130_fd_sc_hd__buf_8 fanout797 (.A(_07400_),
    .X(net797));
 sky130_fd_sc_hd__buf_4 fanout798 (.A(_07400_),
    .X(net798));
 sky130_fd_sc_hd__buf_12 fanout799 (.A(net801),
    .X(net799));
 sky130_fd_sc_hd__buf_6 fanout800 (.A(net801),
    .X(net800));
 sky130_fd_sc_hd__buf_6 fanout801 (.A(_07389_),
    .X(net801));
 sky130_fd_sc_hd__buf_4 fanout802 (.A(net803),
    .X(net802));
 sky130_fd_sc_hd__buf_6 fanout803 (.A(_03547_),
    .X(net803));
 sky130_fd_sc_hd__buf_6 fanout804 (.A(net805),
    .X(net804));
 sky130_fd_sc_hd__buf_8 fanout805 (.A(_03547_),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_8 fanout806 (.A(net807),
    .X(net806));
 sky130_fd_sc_hd__buf_4 fanout807 (.A(_08095_),
    .X(net807));
 sky130_fd_sc_hd__buf_4 fanout808 (.A(net809),
    .X(net808));
 sky130_fd_sc_hd__buf_2 fanout809 (.A(net810),
    .X(net809));
 sky130_fd_sc_hd__buf_2 fanout810 (.A(net811),
    .X(net810));
 sky130_fd_sc_hd__buf_6 fanout811 (.A(_07503_),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_8 fanout812 (.A(net813),
    .X(net812));
 sky130_fd_sc_hd__buf_8 fanout813 (.A(net814),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_16 fanout814 (.A(_07476_),
    .X(net814));
 sky130_fd_sc_hd__buf_8 fanout815 (.A(net817),
    .X(net815));
 sky130_fd_sc_hd__buf_4 fanout816 (.A(net817),
    .X(net816));
 sky130_fd_sc_hd__buf_8 fanout817 (.A(_07474_),
    .X(net817));
 sky130_fd_sc_hd__buf_4 fanout818 (.A(_02441_),
    .X(net818));
 sky130_fd_sc_hd__buf_2 fanout819 (.A(_02441_),
    .X(net819));
 sky130_fd_sc_hd__buf_6 fanout820 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__clkbuf_8 fanout821 (.A(net823),
    .X(net821));
 sky130_fd_sc_hd__buf_8 fanout822 (.A(net823),
    .X(net822));
 sky130_fd_sc_hd__buf_6 fanout823 (.A(_09357_),
    .X(net823));
 sky130_fd_sc_hd__buf_4 fanout824 (.A(_09353_),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_16 fanout825 (.A(_09224_),
    .X(net825));
 sky130_fd_sc_hd__buf_4 fanout826 (.A(_09224_),
    .X(net826));
 sky130_fd_sc_hd__buf_6 fanout827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_4 fanout828 (.A(net829),
    .X(net828));
 sky130_fd_sc_hd__buf_2 fanout829 (.A(net830),
    .X(net829));
 sky130_fd_sc_hd__buf_4 fanout830 (.A(net831),
    .X(net830));
 sky130_fd_sc_hd__buf_4 fanout831 (.A(_06698_),
    .X(net831));
 sky130_fd_sc_hd__buf_8 fanout832 (.A(_04353_),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_8 fanout833 (.A(_04353_),
    .X(net833));
 sky130_fd_sc_hd__buf_6 fanout834 (.A(net835),
    .X(net834));
 sky130_fd_sc_hd__buf_6 fanout835 (.A(_04128_),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_16 fanout836 (.A(_04128_),
    .X(net836));
 sky130_fd_sc_hd__buf_4 fanout837 (.A(_04128_),
    .X(net837));
 sky130_fd_sc_hd__buf_4 fanout838 (.A(net841),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_4 fanout839 (.A(net841),
    .X(net839));
 sky130_fd_sc_hd__buf_6 fanout840 (.A(net841),
    .X(net840));
 sky130_fd_sc_hd__buf_6 fanout841 (.A(_03959_),
    .X(net841));
 sky130_fd_sc_hd__buf_4 fanout842 (.A(net843),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_4 fanout843 (.A(net844),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_4 fanout844 (.A(net846),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_8 fanout845 (.A(net846),
    .X(net845));
 sky130_fd_sc_hd__buf_4 fanout846 (.A(_03890_),
    .X(net846));
 sky130_fd_sc_hd__buf_6 fanout847 (.A(net849),
    .X(net847));
 sky130_fd_sc_hd__buf_6 fanout848 (.A(net849),
    .X(net848));
 sky130_fd_sc_hd__buf_6 fanout849 (.A(_03890_),
    .X(net849));
 sky130_fd_sc_hd__buf_8 fanout850 (.A(_03755_),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_4 fanout851 (.A(_03755_),
    .X(net851));
 sky130_fd_sc_hd__buf_6 fanout852 (.A(net853),
    .X(net852));
 sky130_fd_sc_hd__buf_6 fanout853 (.A(_03755_),
    .X(net853));
 sky130_fd_sc_hd__buf_6 fanout854 (.A(net857),
    .X(net854));
 sky130_fd_sc_hd__buf_6 fanout855 (.A(net856),
    .X(net855));
 sky130_fd_sc_hd__buf_6 fanout856 (.A(net857),
    .X(net856));
 sky130_fd_sc_hd__buf_8 fanout857 (.A(_09355_),
    .X(net857));
 sky130_fd_sc_hd__buf_6 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_8 fanout859 (.A(net861),
    .X(net859));
 sky130_fd_sc_hd__buf_8 fanout860 (.A(net861),
    .X(net860));
 sky130_fd_sc_hd__buf_6 fanout861 (.A(_09304_),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_8 fanout862 (.A(net863),
    .X(net862));
 sky130_fd_sc_hd__buf_6 fanout863 (.A(net865),
    .X(net863));
 sky130_fd_sc_hd__buf_6 fanout864 (.A(net865),
    .X(net864));
 sky130_fd_sc_hd__buf_8 fanout865 (.A(_09303_),
    .X(net865));
 sky130_fd_sc_hd__buf_8 fanout866 (.A(net867),
    .X(net866));
 sky130_fd_sc_hd__buf_8 fanout867 (.A(net869),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_16 fanout868 (.A(net869),
    .X(net868));
 sky130_fd_sc_hd__buf_8 fanout869 (.A(_09297_),
    .X(net869));
 sky130_fd_sc_hd__buf_6 fanout870 (.A(net871),
    .X(net870));
 sky130_fd_sc_hd__buf_6 fanout871 (.A(net873),
    .X(net871));
 sky130_fd_sc_hd__buf_8 fanout872 (.A(net873),
    .X(net872));
 sky130_fd_sc_hd__buf_8 fanout873 (.A(_09294_),
    .X(net873));
 sky130_fd_sc_hd__buf_4 fanout874 (.A(net875),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_4 fanout875 (.A(_09288_),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_8 fanout876 (.A(net877),
    .X(net876));
 sky130_fd_sc_hd__buf_4 fanout877 (.A(_09288_),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_4 fanout878 (.A(net879),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_4 fanout879 (.A(_09280_),
    .X(net879));
 sky130_fd_sc_hd__buf_6 fanout880 (.A(net881),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_8 fanout881 (.A(_09280_),
    .X(net881));
 sky130_fd_sc_hd__buf_4 fanout882 (.A(net883),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_4 fanout883 (.A(net884),
    .X(net883));
 sky130_fd_sc_hd__buf_6 fanout884 (.A(_09279_),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_8 fanout885 (.A(_06101_),
    .X(net885));
 sky130_fd_sc_hd__buf_4 fanout886 (.A(_05931_),
    .X(net886));
 sky130_fd_sc_hd__buf_4 fanout887 (.A(_05931_),
    .X(net887));
 sky130_fd_sc_hd__buf_6 fanout888 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__buf_4 fanout889 (.A(_04033_),
    .X(net889));
 sky130_fd_sc_hd__buf_6 fanout890 (.A(_04033_),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_4 fanout891 (.A(_04033_),
    .X(net891));
 sky130_fd_sc_hd__buf_8 fanout892 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__buf_6 fanout893 (.A(_03924_),
    .X(net893));
 sky130_fd_sc_hd__buf_6 fanout894 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__buf_4 fanout895 (.A(_03924_),
    .X(net895));
 sky130_fd_sc_hd__buf_6 fanout896 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__buf_6 fanout897 (.A(_03109_),
    .X(net897));
 sky130_fd_sc_hd__buf_6 fanout898 (.A(_03109_),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_8 fanout899 (.A(net900),
    .X(net899));
 sky130_fd_sc_hd__buf_6 fanout900 (.A(net902),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_16 fanout901 (.A(net902),
    .X(net901));
 sky130_fd_sc_hd__buf_6 fanout902 (.A(_09360_),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_8 fanout903 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__buf_6 fanout904 (.A(net906),
    .X(net904));
 sky130_fd_sc_hd__clkbuf_16 fanout905 (.A(net906),
    .X(net905));
 sky130_fd_sc_hd__buf_6 fanout906 (.A(_09358_),
    .X(net906));
 sky130_fd_sc_hd__buf_6 fanout907 (.A(net908),
    .X(net907));
 sky130_fd_sc_hd__buf_4 fanout908 (.A(_09336_),
    .X(net908));
 sky130_fd_sc_hd__buf_6 fanout909 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_4 fanout910 (.A(_09336_),
    .X(net910));
 sky130_fd_sc_hd__buf_6 fanout911 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__clkbuf_8 fanout912 (.A(net913),
    .X(net912));
 sky130_fd_sc_hd__buf_6 fanout913 (.A(_09335_),
    .X(net913));
 sky130_fd_sc_hd__buf_4 fanout914 (.A(net915),
    .X(net914));
 sky130_fd_sc_hd__buf_8 fanout915 (.A(net916),
    .X(net915));
 sky130_fd_sc_hd__buf_6 fanout916 (.A(net917),
    .X(net916));
 sky130_fd_sc_hd__buf_12 fanout917 (.A(_09286_),
    .X(net917));
 sky130_fd_sc_hd__buf_4 fanout918 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__buf_8 fanout919 (.A(net920),
    .X(net919));
 sky130_fd_sc_hd__buf_6 fanout920 (.A(net921),
    .X(net920));
 sky130_fd_sc_hd__buf_12 fanout921 (.A(_09285_),
    .X(net921));
 sky130_fd_sc_hd__buf_6 fanout922 (.A(_09278_),
    .X(net922));
 sky130_fd_sc_hd__buf_4 fanout923 (.A(net924),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_4 fanout924 (.A(_09275_),
    .X(net924));
 sky130_fd_sc_hd__buf_6 fanout925 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__buf_4 fanout926 (.A(_09275_),
    .X(net926));
 sky130_fd_sc_hd__buf_4 fanout927 (.A(net928),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_4 fanout928 (.A(_09273_),
    .X(net928));
 sky130_fd_sc_hd__buf_6 fanout929 (.A(net930),
    .X(net929));
 sky130_fd_sc_hd__buf_4 fanout930 (.A(_09273_),
    .X(net930));
 sky130_fd_sc_hd__buf_6 fanout931 (.A(_06196_),
    .X(net931));
 sky130_fd_sc_hd__buf_8 fanout932 (.A(net934),
    .X(net932));
 sky130_fd_sc_hd__buf_6 fanout933 (.A(net934),
    .X(net933));
 sky130_fd_sc_hd__buf_4 fanout934 (.A(_06195_),
    .X(net934));
 sky130_fd_sc_hd__buf_6 fanout935 (.A(net938),
    .X(net935));
 sky130_fd_sc_hd__clkbuf_4 fanout936 (.A(net938),
    .X(net936));
 sky130_fd_sc_hd__buf_4 fanout937 (.A(net938),
    .X(net937));
 sky130_fd_sc_hd__buf_4 fanout938 (.A(_06100_),
    .X(net938));
 sky130_fd_sc_hd__buf_4 fanout939 (.A(net941),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_4 fanout940 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__clkbuf_8 fanout941 (.A(net943),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_8 fanout942 (.A(net943),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_4 fanout943 (.A(_06015_),
    .X(net943));
 sky130_fd_sc_hd__buf_4 fanout944 (.A(net945),
    .X(net944));
 sky130_fd_sc_hd__buf_6 fanout945 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__buf_6 fanout946 (.A(_05930_),
    .X(net946));
 sky130_fd_sc_hd__buf_6 fanout947 (.A(_05847_),
    .X(net947));
 sky130_fd_sc_hd__buf_6 fanout948 (.A(_05847_),
    .X(net948));
 sky130_fd_sc_hd__buf_8 fanout949 (.A(_05846_),
    .X(net949));
 sky130_fd_sc_hd__buf_12 fanout950 (.A(_05846_),
    .X(net950));
 sky130_fd_sc_hd__buf_6 fanout951 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__buf_4 fanout952 (.A(_08773_),
    .X(net952));
 sky130_fd_sc_hd__buf_6 fanout953 (.A(_08773_),
    .X(net953));
 sky130_fd_sc_hd__buf_4 fanout954 (.A(net956),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_2 fanout955 (.A(net956),
    .X(net955));
 sky130_fd_sc_hd__buf_8 fanout956 (.A(_08772_),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_4 fanout957 (.A(net958),
    .X(net957));
 sky130_fd_sc_hd__buf_2 fanout958 (.A(net961),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_4 fanout959 (.A(net961),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_2 fanout960 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__buf_6 fanout961 (.A(_06244_),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 fanout962 (.A(net964),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_4 fanout963 (.A(net964),
    .X(net963));
 sky130_fd_sc_hd__buf_4 fanout964 (.A(net965),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_8 fanout965 (.A(_05475_),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_4 fanout966 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__buf_2 fanout967 (.A(net968),
    .X(net967));
 sky130_fd_sc_hd__buf_2 fanout968 (.A(_05387_),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_4 fanout969 (.A(_05387_),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_4 fanout970 (.A(net972),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_2 fanout971 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__buf_4 fanout972 (.A(net973),
    .X(net972));
 sky130_fd_sc_hd__buf_6 fanout973 (.A(_05299_),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_4 fanout974 (.A(net977),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_2 fanout975 (.A(net977),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_4 fanout976 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__buf_2 fanout977 (.A(net978),
    .X(net977));
 sky130_fd_sc_hd__buf_6 fanout978 (.A(_05207_),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_4 fanout979 (.A(net980),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_4 fanout980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__buf_4 fanout981 (.A(net982),
    .X(net981));
 sky130_fd_sc_hd__buf_6 fanout982 (.A(_05120_),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout983 (.A(net984),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_4 fanout984 (.A(_05041_),
    .X(net984));
 sky130_fd_sc_hd__buf_6 fanout985 (.A(_05041_),
    .X(net985));
 sky130_fd_sc_hd__buf_2 fanout986 (.A(_05041_),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_4 fanout987 (.A(net989),
    .X(net987));
 sky130_fd_sc_hd__buf_2 fanout988 (.A(net989),
    .X(net988));
 sky130_fd_sc_hd__buf_4 fanout989 (.A(net990),
    .X(net989));
 sky130_fd_sc_hd__buf_4 fanout990 (.A(_04958_),
    .X(net990));
 sky130_fd_sc_hd__buf_4 fanout991 (.A(net992),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_4 fanout992 (.A(_03110_),
    .X(net992));
 sky130_fd_sc_hd__buf_4 fanout993 (.A(net994),
    .X(net993));
 sky130_fd_sc_hd__buf_4 fanout994 (.A(_03110_),
    .X(net994));
 sky130_fd_sc_hd__buf_4 fanout995 (.A(net996),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_4 fanout996 (.A(_03100_),
    .X(net996));
 sky130_fd_sc_hd__buf_4 fanout997 (.A(net998),
    .X(net997));
 sky130_fd_sc_hd__buf_4 fanout998 (.A(_03100_),
    .X(net998));
 sky130_fd_sc_hd__buf_6 fanout999 (.A(net1001),
    .X(net999));
 sky130_fd_sc_hd__buf_6 input1 (.A(coreIndex[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input10 (.A(core_wb_data_i[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(dout0[61]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(dout0[62]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(dout0[63]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(dout0[6]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(dout0[7]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(dout0[8]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 input106 (.A(dout0[9]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(dout1[0]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(dout1[10]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(dout1[11]),
    .X(net109));
 sky130_fd_sc_hd__buf_4 input11 (.A(core_wb_data_i[10]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(dout1[12]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(dout1[13]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(dout1[14]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(dout1[15]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(dout1[16]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(dout1[17]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(dout1[18]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(dout1[19]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(dout1[1]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(dout1[20]),
    .X(net119));
 sky130_fd_sc_hd__buf_4 input12 (.A(core_wb_data_i[11]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(dout1[21]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(dout1[22]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(dout1[23]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(dout1[24]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(dout1[25]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(dout1[26]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(dout1[27]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(dout1[28]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(dout1[29]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(dout1[2]),
    .X(net129));
 sky130_fd_sc_hd__buf_4 input13 (.A(core_wb_data_i[12]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(dout1[30]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(dout1[31]),
    .X(net131));
 sky130_fd_sc_hd__buf_2 input132 (.A(dout1[32]),
    .X(net132));
 sky130_fd_sc_hd__buf_2 input133 (.A(dout1[33]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 input134 (.A(dout1[34]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 input135 (.A(dout1[35]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(dout1[36]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(dout1[37]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_2 input138 (.A(dout1[38]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 input139 (.A(dout1[39]),
    .X(net139));
 sky130_fd_sc_hd__buf_4 input14 (.A(core_wb_data_i[13]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input140 (.A(dout1[3]),
    .X(net140));
 sky130_fd_sc_hd__buf_2 input141 (.A(dout1[40]),
    .X(net141));
 sky130_fd_sc_hd__buf_2 input142 (.A(dout1[41]),
    .X(net142));
 sky130_fd_sc_hd__buf_2 input143 (.A(dout1[42]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 input144 (.A(dout1[43]),
    .X(net144));
 sky130_fd_sc_hd__buf_2 input145 (.A(dout1[44]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 input146 (.A(dout1[45]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(dout1[46]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 input148 (.A(dout1[47]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 input149 (.A(dout1[48]),
    .X(net149));
 sky130_fd_sc_hd__buf_4 input15 (.A(core_wb_data_i[14]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input150 (.A(dout1[49]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_2 input151 (.A(dout1[4]),
    .X(net151));
 sky130_fd_sc_hd__buf_2 input152 (.A(dout1[50]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_2 input153 (.A(dout1[51]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 input154 (.A(dout1[52]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 input155 (.A(dout1[53]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 input156 (.A(dout1[54]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 input157 (.A(dout1[55]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 input158 (.A(dout1[56]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(dout1[57]),
    .X(net159));
 sky130_fd_sc_hd__buf_4 input16 (.A(core_wb_data_i[15]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input160 (.A(dout1[58]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 input161 (.A(dout1[59]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 input162 (.A(dout1[5]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(dout1[60]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 input164 (.A(dout1[61]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 input165 (.A(dout1[62]),
    .X(net165));
 sky130_fd_sc_hd__buf_2 input166 (.A(dout1[63]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 input167 (.A(dout1[6]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 input168 (.A(dout1[7]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 input169 (.A(dout1[8]),
    .X(net169));
 sky130_fd_sc_hd__buf_4 input17 (.A(core_wb_data_i[16]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input170 (.A(dout1[9]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 input171 (.A(irq[0]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(irq[10]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 input173 (.A(irq[11]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 input174 (.A(irq[12]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 input175 (.A(irq[13]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 input176 (.A(irq[14]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 input177 (.A(irq[15]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 input178 (.A(irq[1]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 input179 (.A(irq[2]),
    .X(net179));
 sky130_fd_sc_hd__buf_4 input18 (.A(core_wb_data_i[17]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(irq[3]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 input181 (.A(irq[4]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 input182 (.A(irq[5]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 input183 (.A(irq[6]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 input184 (.A(irq[7]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 input185 (.A(irq[8]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(irq[9]),
    .X(net186));
 sky130_fd_sc_hd__buf_4 input187 (.A(jtag_tck),
    .X(net187));
 sky130_fd_sc_hd__buf_12 input188 (.A(jtag_tdi),
    .X(net188));
 sky130_fd_sc_hd__buf_6 input189 (.A(jtag_tms),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(core_wb_data_i[18]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(localMemory_wb_adr_i[0]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 input191 (.A(localMemory_wb_adr_i[10]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 input192 (.A(localMemory_wb_adr_i[11]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 input193 (.A(localMemory_wb_adr_i[12]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 input194 (.A(localMemory_wb_adr_i[13]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 input195 (.A(localMemory_wb_adr_i[14]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 input196 (.A(localMemory_wb_adr_i[15]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 input197 (.A(localMemory_wb_adr_i[16]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(localMemory_wb_adr_i[17]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 input199 (.A(localMemory_wb_adr_i[18]),
    .X(net199));
 sky130_fd_sc_hd__buf_6 input2 (.A(coreIndex[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input20 (.A(core_wb_data_i[19]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input200 (.A(localMemory_wb_adr_i[19]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 input201 (.A(localMemory_wb_adr_i[1]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 input202 (.A(localMemory_wb_adr_i[20]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 input203 (.A(localMemory_wb_adr_i[21]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 input204 (.A(localMemory_wb_adr_i[22]),
    .X(net204));
 sky130_fd_sc_hd__buf_6 input205 (.A(localMemory_wb_adr_i[23]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 input206 (.A(localMemory_wb_adr_i[2]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 input207 (.A(localMemory_wb_adr_i[3]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 input208 (.A(localMemory_wb_adr_i[4]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 input209 (.A(localMemory_wb_adr_i[5]),
    .X(net209));
 sky130_fd_sc_hd__buf_4 input21 (.A(core_wb_data_i[1]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input210 (.A(localMemory_wb_adr_i[6]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 input211 (.A(localMemory_wb_adr_i[7]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 input212 (.A(localMemory_wb_adr_i[8]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(localMemory_wb_adr_i[9]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 input214 (.A(localMemory_wb_cyc_i),
    .X(net214));
 sky130_fd_sc_hd__buf_12 input215 (.A(localMemory_wb_data_i[0]),
    .X(net215));
 sky130_fd_sc_hd__buf_12 input216 (.A(localMemory_wb_data_i[10]),
    .X(net216));
 sky130_fd_sc_hd__buf_12 input217 (.A(localMemory_wb_data_i[11]),
    .X(net217));
 sky130_fd_sc_hd__buf_12 input218 (.A(localMemory_wb_data_i[12]),
    .X(net218));
 sky130_fd_sc_hd__buf_12 input219 (.A(localMemory_wb_data_i[13]),
    .X(net219));
 sky130_fd_sc_hd__buf_4 input22 (.A(core_wb_data_i[20]),
    .X(net22));
 sky130_fd_sc_hd__buf_12 input220 (.A(localMemory_wb_data_i[14]),
    .X(net220));
 sky130_fd_sc_hd__buf_12 input221 (.A(localMemory_wb_data_i[15]),
    .X(net221));
 sky130_fd_sc_hd__buf_12 input222 (.A(localMemory_wb_data_i[16]),
    .X(net222));
 sky130_fd_sc_hd__buf_12 input223 (.A(localMemory_wb_data_i[17]),
    .X(net223));
 sky130_fd_sc_hd__buf_12 input224 (.A(localMemory_wb_data_i[18]),
    .X(net224));
 sky130_fd_sc_hd__buf_12 input225 (.A(localMemory_wb_data_i[19]),
    .X(net225));
 sky130_fd_sc_hd__buf_12 input226 (.A(localMemory_wb_data_i[1]),
    .X(net226));
 sky130_fd_sc_hd__buf_12 input227 (.A(localMemory_wb_data_i[20]),
    .X(net227));
 sky130_fd_sc_hd__buf_12 input228 (.A(localMemory_wb_data_i[21]),
    .X(net228));
 sky130_fd_sc_hd__buf_12 input229 (.A(localMemory_wb_data_i[22]),
    .X(net229));
 sky130_fd_sc_hd__buf_4 input23 (.A(core_wb_data_i[21]),
    .X(net23));
 sky130_fd_sc_hd__buf_12 input230 (.A(localMemory_wb_data_i[23]),
    .X(net230));
 sky130_fd_sc_hd__buf_12 input231 (.A(localMemory_wb_data_i[24]),
    .X(net231));
 sky130_fd_sc_hd__buf_12 input232 (.A(localMemory_wb_data_i[25]),
    .X(net232));
 sky130_fd_sc_hd__buf_12 input233 (.A(localMemory_wb_data_i[26]),
    .X(net233));
 sky130_fd_sc_hd__buf_12 input234 (.A(localMemory_wb_data_i[27]),
    .X(net234));
 sky130_fd_sc_hd__buf_12 input235 (.A(localMemory_wb_data_i[28]),
    .X(net235));
 sky130_fd_sc_hd__buf_12 input236 (.A(localMemory_wb_data_i[29]),
    .X(net236));
 sky130_fd_sc_hd__buf_12 input237 (.A(localMemory_wb_data_i[2]),
    .X(net237));
 sky130_fd_sc_hd__buf_12 input238 (.A(localMemory_wb_data_i[30]),
    .X(net238));
 sky130_fd_sc_hd__buf_12 input239 (.A(localMemory_wb_data_i[31]),
    .X(net239));
 sky130_fd_sc_hd__buf_4 input24 (.A(core_wb_data_i[22]),
    .X(net24));
 sky130_fd_sc_hd__buf_12 input240 (.A(localMemory_wb_data_i[3]),
    .X(net240));
 sky130_fd_sc_hd__buf_12 input241 (.A(localMemory_wb_data_i[4]),
    .X(net241));
 sky130_fd_sc_hd__buf_12 input242 (.A(localMemory_wb_data_i[5]),
    .X(net242));
 sky130_fd_sc_hd__buf_12 input243 (.A(localMemory_wb_data_i[6]),
    .X(net243));
 sky130_fd_sc_hd__buf_12 input244 (.A(localMemory_wb_data_i[7]),
    .X(net244));
 sky130_fd_sc_hd__buf_12 input245 (.A(localMemory_wb_data_i[8]),
    .X(net245));
 sky130_fd_sc_hd__buf_12 input246 (.A(localMemory_wb_data_i[9]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 input247 (.A(localMemory_wb_sel_i[0]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 input248 (.A(localMemory_wb_sel_i[1]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 input249 (.A(localMemory_wb_sel_i[2]),
    .X(net249));
 sky130_fd_sc_hd__buf_4 input25 (.A(core_wb_data_i[23]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input250 (.A(localMemory_wb_sel_i[3]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 input251 (.A(localMemory_wb_stb_i),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 input252 (.A(localMemory_wb_we_i),
    .X(net252));
 sky130_fd_sc_hd__buf_4 input253 (.A(manufacturerID[0]),
    .X(net253));
 sky130_fd_sc_hd__buf_2 input254 (.A(manufacturerID[10]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_4 input255 (.A(manufacturerID[1]),
    .X(net255));
 sky130_fd_sc_hd__buf_2 input256 (.A(manufacturerID[2]),
    .X(net256));
 sky130_fd_sc_hd__buf_2 input257 (.A(manufacturerID[3]),
    .X(net257));
 sky130_fd_sc_hd__buf_2 input258 (.A(manufacturerID[4]),
    .X(net258));
 sky130_fd_sc_hd__buf_2 input259 (.A(manufacturerID[5]),
    .X(net259));
 sky130_fd_sc_hd__buf_4 input26 (.A(core_wb_data_i[24]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input260 (.A(manufacturerID[6]),
    .X(net260));
 sky130_fd_sc_hd__buf_2 input261 (.A(manufacturerID[7]),
    .X(net261));
 sky130_fd_sc_hd__buf_2 input262 (.A(manufacturerID[8]),
    .X(net262));
 sky130_fd_sc_hd__buf_2 input263 (.A(manufacturerID[9]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_4 input264 (.A(partID[0]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 input265 (.A(partID[10]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_2 input266 (.A(partID[11]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 input267 (.A(partID[12]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 input268 (.A(partID[13]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 input269 (.A(partID[14]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(core_wb_data_i[25]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input270 (.A(partID[15]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 input271 (.A(partID[1]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 input272 (.A(partID[2]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_2 input273 (.A(partID[3]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_2 input274 (.A(partID[4]),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 input275 (.A(partID[5]),
    .X(net275));
 sky130_fd_sc_hd__buf_2 input276 (.A(partID[6]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 input277 (.A(partID[7]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_2 input278 (.A(partID[8]),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 input279 (.A(partID[9]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(core_wb_data_i[26]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input280 (.A(versionID[0]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 input281 (.A(versionID[1]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 input282 (.A(versionID[2]),
    .X(net282));
 sky130_fd_sc_hd__buf_2 input283 (.A(versionID[3]),
    .X(net283));
 sky130_fd_sc_hd__buf_12 input284 (.A(wb_rst_i),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(core_wb_data_i[27]),
    .X(net29));
 sky130_fd_sc_hd__buf_6 input3 (.A(coreIndex[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(core_wb_data_i[28]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(core_wb_data_i[29]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_8 input32 (.A(core_wb_data_i[2]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 input33 (.A(core_wb_data_i[30]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(core_wb_data_i[31]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(core_wb_data_i[3]),
    .X(net35));
 sky130_fd_sc_hd__buf_6 input36 (.A(core_wb_data_i[4]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(core_wb_data_i[5]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(core_wb_data_i[6]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(core_wb_data_i[7]),
    .X(net39));
 sky130_fd_sc_hd__buf_6 input4 (.A(coreIndex[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(core_wb_data_i[8]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(core_wb_data_i[9]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(core_wb_error_i),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(dout0[0]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(dout0[10]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(dout0[11]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(dout0[12]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(dout0[13]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(dout0[14]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(dout0[15]),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input5 (.A(coreIndex[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(dout0[16]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(dout0[17]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(dout0[18]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(dout0[19]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(dout0[1]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(dout0[20]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(dout0[21]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(dout0[22]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(dout0[23]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(dout0[24]),
    .X(net59));
 sky130_fd_sc_hd__buf_4 input6 (.A(coreIndex[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(dout0[25]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(dout0[26]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(dout0[27]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(dout0[28]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(dout0[29]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(dout0[2]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(dout0[30]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(dout0[31]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(dout0[32]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(dout0[33]),
    .X(net69));
 sky130_fd_sc_hd__buf_4 input7 (.A(coreIndex[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(dout0[34]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(dout0[35]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(dout0[36]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(dout0[37]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(dout0[38]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(dout0[39]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(dout0[3]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(dout0[40]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(dout0[41]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(dout0[42]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(coreIndex[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(dout0[43]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(dout0[44]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(dout0[45]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(dout0[46]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(dout0[47]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(dout0[48]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(dout0[49]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(dout0[4]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(dout0[50]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(dout0[51]),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input9 (.A(core_wb_ack_i),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(dout0[52]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input91 (.A(dout0[53]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(dout0[54]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 input93 (.A(dout0[55]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(dout0[56]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(dout0[57]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(dout0[58]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(dout0[59]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(dout0[5]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(dout0[60]),
    .X(net99));
 sky130_fd_sc_hd__buf_6 max_cap1275 (.A(_04467_),
    .X(net1275));
 sky130_fd_sc_hd__buf_12 max_cap1805 (.A(\localMemoryInterface.lastRBankSelect ),
    .X(net1805));
 sky130_fd_sc_hd__buf_4 output285 (.A(net285),
    .X(addr0[0]));
 sky130_fd_sc_hd__buf_4 output286 (.A(net286),
    .X(addr0[1]));
 sky130_fd_sc_hd__buf_4 output287 (.A(net287),
    .X(addr0[2]));
 sky130_fd_sc_hd__buf_4 output288 (.A(net288),
    .X(addr0[3]));
 sky130_fd_sc_hd__buf_4 output289 (.A(net289),
    .X(addr0[4]));
 sky130_fd_sc_hd__buf_4 output290 (.A(net290),
    .X(addr0[5]));
 sky130_fd_sc_hd__buf_4 output291 (.A(net291),
    .X(addr0[6]));
 sky130_fd_sc_hd__buf_4 output292 (.A(net292),
    .X(addr0[7]));
 sky130_fd_sc_hd__buf_4 output293 (.A(net293),
    .X(addr0[8]));
 sky130_fd_sc_hd__buf_4 output294 (.A(net294),
    .X(addr1[0]));
 sky130_fd_sc_hd__buf_4 output295 (.A(net295),
    .X(addr1[1]));
 sky130_fd_sc_hd__buf_4 output296 (.A(net296),
    .X(addr1[2]));
 sky130_fd_sc_hd__buf_4 output297 (.A(net297),
    .X(addr1[3]));
 sky130_fd_sc_hd__buf_4 output298 (.A(net298),
    .X(addr1[4]));
 sky130_fd_sc_hd__buf_4 output299 (.A(net299),
    .X(addr1[5]));
 sky130_fd_sc_hd__buf_4 output300 (.A(net300),
    .X(addr1[6]));
 sky130_fd_sc_hd__buf_4 output301 (.A(net301),
    .X(addr1[7]));
 sky130_fd_sc_hd__buf_4 output302 (.A(net302),
    .X(addr1[8]));
 sky130_fd_sc_hd__clkbuf_2 output303 (.A(net303),
    .X(clk0));
 sky130_fd_sc_hd__clkbuf_2 output304 (.A(net304),
    .X(clk1));
 sky130_fd_sc_hd__buf_4 output305 (.A(net305),
    .X(core_wb_adr_o[0]));
 sky130_fd_sc_hd__buf_4 output306 (.A(net306),
    .X(core_wb_adr_o[10]));
 sky130_fd_sc_hd__buf_4 output307 (.A(net307),
    .X(core_wb_adr_o[11]));
 sky130_fd_sc_hd__buf_4 output308 (.A(net308),
    .X(core_wb_adr_o[12]));
 sky130_fd_sc_hd__buf_4 output309 (.A(net309),
    .X(core_wb_adr_o[13]));
 sky130_fd_sc_hd__buf_4 output310 (.A(net310),
    .X(core_wb_adr_o[14]));
 sky130_fd_sc_hd__buf_4 output311 (.A(net311),
    .X(core_wb_adr_o[15]));
 sky130_fd_sc_hd__buf_4 output312 (.A(net312),
    .X(core_wb_adr_o[16]));
 sky130_fd_sc_hd__buf_4 output313 (.A(net313),
    .X(core_wb_adr_o[17]));
 sky130_fd_sc_hd__buf_4 output314 (.A(net314),
    .X(core_wb_adr_o[18]));
 sky130_fd_sc_hd__buf_4 output315 (.A(net315),
    .X(core_wb_adr_o[19]));
 sky130_fd_sc_hd__buf_4 output316 (.A(net316),
    .X(core_wb_adr_o[1]));
 sky130_fd_sc_hd__buf_4 output317 (.A(net317),
    .X(core_wb_adr_o[20]));
 sky130_fd_sc_hd__buf_4 output318 (.A(net318),
    .X(core_wb_adr_o[21]));
 sky130_fd_sc_hd__buf_4 output319 (.A(net319),
    .X(core_wb_adr_o[22]));
 sky130_fd_sc_hd__buf_4 output320 (.A(net320),
    .X(core_wb_adr_o[23]));
 sky130_fd_sc_hd__buf_4 output321 (.A(net321),
    .X(core_wb_adr_o[24]));
 sky130_fd_sc_hd__buf_4 output322 (.A(net322),
    .X(core_wb_adr_o[25]));
 sky130_fd_sc_hd__buf_4 output323 (.A(net323),
    .X(core_wb_adr_o[26]));
 sky130_fd_sc_hd__buf_4 output324 (.A(net324),
    .X(core_wb_adr_o[27]));
 sky130_fd_sc_hd__buf_4 output325 (.A(net325),
    .X(core_wb_adr_o[2]));
 sky130_fd_sc_hd__buf_4 output326 (.A(net326),
    .X(core_wb_adr_o[3]));
 sky130_fd_sc_hd__buf_4 output327 (.A(net327),
    .X(core_wb_adr_o[4]));
 sky130_fd_sc_hd__buf_4 output328 (.A(net328),
    .X(core_wb_adr_o[5]));
 sky130_fd_sc_hd__buf_4 output329 (.A(net329),
    .X(core_wb_adr_o[6]));
 sky130_fd_sc_hd__buf_4 output330 (.A(net330),
    .X(core_wb_adr_o[7]));
 sky130_fd_sc_hd__buf_4 output331 (.A(net331),
    .X(core_wb_adr_o[8]));
 sky130_fd_sc_hd__buf_4 output332 (.A(net332),
    .X(core_wb_adr_o[9]));
 sky130_fd_sc_hd__buf_4 output333 (.A(net333),
    .X(core_wb_cyc_o));
 sky130_fd_sc_hd__buf_4 output334 (.A(net334),
    .X(core_wb_data_o[0]));
 sky130_fd_sc_hd__buf_4 output335 (.A(net335),
    .X(core_wb_data_o[10]));
 sky130_fd_sc_hd__buf_4 output336 (.A(net336),
    .X(core_wb_data_o[11]));
 sky130_fd_sc_hd__buf_4 output337 (.A(net337),
    .X(core_wb_data_o[12]));
 sky130_fd_sc_hd__buf_4 output338 (.A(net338),
    .X(core_wb_data_o[13]));
 sky130_fd_sc_hd__buf_4 output339 (.A(net339),
    .X(core_wb_data_o[14]));
 sky130_fd_sc_hd__buf_4 output340 (.A(net340),
    .X(core_wb_data_o[15]));
 sky130_fd_sc_hd__buf_4 output341 (.A(net341),
    .X(core_wb_data_o[16]));
 sky130_fd_sc_hd__buf_4 output342 (.A(net342),
    .X(core_wb_data_o[17]));
 sky130_fd_sc_hd__buf_4 output343 (.A(net343),
    .X(core_wb_data_o[18]));
 sky130_fd_sc_hd__buf_4 output344 (.A(net344),
    .X(core_wb_data_o[19]));
 sky130_fd_sc_hd__buf_4 output345 (.A(net345),
    .X(core_wb_data_o[1]));
 sky130_fd_sc_hd__buf_4 output346 (.A(net346),
    .X(core_wb_data_o[20]));
 sky130_fd_sc_hd__buf_4 output347 (.A(net347),
    .X(core_wb_data_o[21]));
 sky130_fd_sc_hd__buf_4 output348 (.A(net348),
    .X(core_wb_data_o[22]));
 sky130_fd_sc_hd__buf_4 output349 (.A(net349),
    .X(core_wb_data_o[23]));
 sky130_fd_sc_hd__buf_4 output350 (.A(net350),
    .X(core_wb_data_o[24]));
 sky130_fd_sc_hd__buf_4 output351 (.A(net351),
    .X(core_wb_data_o[25]));
 sky130_fd_sc_hd__buf_4 output352 (.A(net352),
    .X(core_wb_data_o[26]));
 sky130_fd_sc_hd__buf_4 output353 (.A(net353),
    .X(core_wb_data_o[27]));
 sky130_fd_sc_hd__buf_4 output354 (.A(net354),
    .X(core_wb_data_o[28]));
 sky130_fd_sc_hd__buf_4 output355 (.A(net355),
    .X(core_wb_data_o[29]));
 sky130_fd_sc_hd__buf_4 output356 (.A(net356),
    .X(core_wb_data_o[2]));
 sky130_fd_sc_hd__buf_4 output357 (.A(net357),
    .X(core_wb_data_o[30]));
 sky130_fd_sc_hd__buf_4 output358 (.A(net358),
    .X(core_wb_data_o[31]));
 sky130_fd_sc_hd__buf_4 output359 (.A(net359),
    .X(core_wb_data_o[3]));
 sky130_fd_sc_hd__buf_4 output360 (.A(net360),
    .X(core_wb_data_o[4]));
 sky130_fd_sc_hd__buf_4 output361 (.A(net361),
    .X(core_wb_data_o[5]));
 sky130_fd_sc_hd__buf_4 output362 (.A(net362),
    .X(core_wb_data_o[6]));
 sky130_fd_sc_hd__buf_4 output363 (.A(net363),
    .X(core_wb_data_o[7]));
 sky130_fd_sc_hd__buf_4 output364 (.A(net364),
    .X(core_wb_data_o[8]));
 sky130_fd_sc_hd__buf_4 output365 (.A(net365),
    .X(core_wb_data_o[9]));
 sky130_fd_sc_hd__buf_4 output366 (.A(net366),
    .X(core_wb_sel_o[0]));
 sky130_fd_sc_hd__buf_4 output367 (.A(net367),
    .X(core_wb_sel_o[1]));
 sky130_fd_sc_hd__buf_4 output368 (.A(net368),
    .X(core_wb_sel_o[2]));
 sky130_fd_sc_hd__buf_4 output369 (.A(net369),
    .X(core_wb_sel_o[3]));
 sky130_fd_sc_hd__buf_4 output370 (.A(net370),
    .X(core_wb_stb_o));
 sky130_fd_sc_hd__buf_4 output371 (.A(net371),
    .X(core_wb_we_o));
 sky130_fd_sc_hd__buf_4 output372 (.A(net372),
    .X(csb0[0]));
 sky130_fd_sc_hd__buf_4 output373 (.A(net373),
    .X(csb0[1]));
 sky130_fd_sc_hd__buf_4 output374 (.A(net374),
    .X(csb1[0]));
 sky130_fd_sc_hd__buf_4 output375 (.A(net375),
    .X(csb1[1]));
 sky130_fd_sc_hd__buf_6 output376 (.A(net376),
    .X(din0[0]));
 sky130_fd_sc_hd__buf_4 output377 (.A(net377),
    .X(din0[10]));
 sky130_fd_sc_hd__buf_4 output378 (.A(net378),
    .X(din0[11]));
 sky130_fd_sc_hd__buf_4 output379 (.A(net379),
    .X(din0[12]));
 sky130_fd_sc_hd__buf_4 output380 (.A(net380),
    .X(din0[13]));
 sky130_fd_sc_hd__buf_4 output381 (.A(net381),
    .X(din0[14]));
 sky130_fd_sc_hd__buf_4 output382 (.A(net382),
    .X(din0[15]));
 sky130_fd_sc_hd__buf_4 output383 (.A(net383),
    .X(din0[16]));
 sky130_fd_sc_hd__buf_4 output384 (.A(net384),
    .X(din0[17]));
 sky130_fd_sc_hd__buf_4 output385 (.A(net385),
    .X(din0[18]));
 sky130_fd_sc_hd__buf_4 output386 (.A(net386),
    .X(din0[19]));
 sky130_fd_sc_hd__buf_6 output387 (.A(net387),
    .X(din0[1]));
 sky130_fd_sc_hd__buf_4 output388 (.A(net388),
    .X(din0[20]));
 sky130_fd_sc_hd__buf_4 output389 (.A(net389),
    .X(din0[21]));
 sky130_fd_sc_hd__buf_4 output390 (.A(net390),
    .X(din0[22]));
 sky130_fd_sc_hd__buf_4 output391 (.A(net391),
    .X(din0[23]));
 sky130_fd_sc_hd__buf_4 output392 (.A(net392),
    .X(din0[24]));
 sky130_fd_sc_hd__buf_4 output393 (.A(net393),
    .X(din0[25]));
 sky130_fd_sc_hd__buf_4 output394 (.A(net394),
    .X(din0[26]));
 sky130_fd_sc_hd__buf_4 output395 (.A(net395),
    .X(din0[27]));
 sky130_fd_sc_hd__buf_4 output396 (.A(net396),
    .X(din0[28]));
 sky130_fd_sc_hd__buf_4 output397 (.A(net397),
    .X(din0[29]));
 sky130_fd_sc_hd__buf_6 output398 (.A(net398),
    .X(din0[2]));
 sky130_fd_sc_hd__buf_4 output399 (.A(net399),
    .X(din0[30]));
 sky130_fd_sc_hd__buf_4 output400 (.A(net400),
    .X(din0[31]));
 sky130_fd_sc_hd__buf_6 output401 (.A(net401),
    .X(din0[3]));
 sky130_fd_sc_hd__buf_4 output402 (.A(net402),
    .X(din0[4]));
 sky130_fd_sc_hd__buf_4 output403 (.A(net403),
    .X(din0[5]));
 sky130_fd_sc_hd__buf_4 output404 (.A(net404),
    .X(din0[6]));
 sky130_fd_sc_hd__buf_4 output405 (.A(net405),
    .X(din0[7]));
 sky130_fd_sc_hd__buf_4 output406 (.A(net406),
    .X(din0[8]));
 sky130_fd_sc_hd__buf_4 output407 (.A(net407),
    .X(din0[9]));
 sky130_fd_sc_hd__buf_4 output408 (.A(net408),
    .X(jtag_tdo));
 sky130_fd_sc_hd__buf_4 output409 (.A(net409),
    .X(localMemory_wb_ack_o));
 sky130_fd_sc_hd__buf_4 output410 (.A(net410),
    .X(localMemory_wb_data_o[0]));
 sky130_fd_sc_hd__buf_4 output411 (.A(net411),
    .X(localMemory_wb_data_o[10]));
 sky130_fd_sc_hd__buf_4 output412 (.A(net412),
    .X(localMemory_wb_data_o[11]));
 sky130_fd_sc_hd__buf_4 output413 (.A(net413),
    .X(localMemory_wb_data_o[12]));
 sky130_fd_sc_hd__buf_4 output414 (.A(net414),
    .X(localMemory_wb_data_o[13]));
 sky130_fd_sc_hd__buf_4 output415 (.A(net415),
    .X(localMemory_wb_data_o[14]));
 sky130_fd_sc_hd__buf_4 output416 (.A(net416),
    .X(localMemory_wb_data_o[15]));
 sky130_fd_sc_hd__buf_4 output417 (.A(net417),
    .X(localMemory_wb_data_o[16]));
 sky130_fd_sc_hd__buf_4 output418 (.A(net418),
    .X(localMemory_wb_data_o[17]));
 sky130_fd_sc_hd__buf_4 output419 (.A(net419),
    .X(localMemory_wb_data_o[18]));
 sky130_fd_sc_hd__buf_4 output420 (.A(net420),
    .X(localMemory_wb_data_o[19]));
 sky130_fd_sc_hd__buf_4 output421 (.A(net421),
    .X(localMemory_wb_data_o[1]));
 sky130_fd_sc_hd__buf_4 output422 (.A(net422),
    .X(localMemory_wb_data_o[20]));
 sky130_fd_sc_hd__buf_4 output423 (.A(net423),
    .X(localMemory_wb_data_o[21]));
 sky130_fd_sc_hd__buf_4 output424 (.A(net424),
    .X(localMemory_wb_data_o[22]));
 sky130_fd_sc_hd__buf_4 output425 (.A(net425),
    .X(localMemory_wb_data_o[23]));
 sky130_fd_sc_hd__buf_4 output426 (.A(net426),
    .X(localMemory_wb_data_o[24]));
 sky130_fd_sc_hd__buf_4 output427 (.A(net427),
    .X(localMemory_wb_data_o[25]));
 sky130_fd_sc_hd__buf_4 output428 (.A(net428),
    .X(localMemory_wb_data_o[26]));
 sky130_fd_sc_hd__buf_4 output429 (.A(net429),
    .X(localMemory_wb_data_o[27]));
 sky130_fd_sc_hd__buf_4 output430 (.A(net430),
    .X(localMemory_wb_data_o[28]));
 sky130_fd_sc_hd__buf_4 output431 (.A(net431),
    .X(localMemory_wb_data_o[29]));
 sky130_fd_sc_hd__buf_4 output432 (.A(net432),
    .X(localMemory_wb_data_o[2]));
 sky130_fd_sc_hd__buf_4 output433 (.A(net433),
    .X(localMemory_wb_data_o[30]));
 sky130_fd_sc_hd__buf_4 output434 (.A(net434),
    .X(localMemory_wb_data_o[31]));
 sky130_fd_sc_hd__buf_4 output435 (.A(net435),
    .X(localMemory_wb_data_o[3]));
 sky130_fd_sc_hd__buf_4 output436 (.A(net436),
    .X(localMemory_wb_data_o[4]));
 sky130_fd_sc_hd__buf_4 output437 (.A(net437),
    .X(localMemory_wb_data_o[5]));
 sky130_fd_sc_hd__buf_4 output438 (.A(net438),
    .X(localMemory_wb_data_o[6]));
 sky130_fd_sc_hd__buf_4 output439 (.A(net439),
    .X(localMemory_wb_data_o[7]));
 sky130_fd_sc_hd__buf_4 output440 (.A(net440),
    .X(localMemory_wb_data_o[8]));
 sky130_fd_sc_hd__buf_4 output441 (.A(net441),
    .X(localMemory_wb_data_o[9]));
 sky130_fd_sc_hd__buf_4 output442 (.A(net442),
    .X(localMemory_wb_stall_o));
 sky130_fd_sc_hd__buf_4 output443 (.A(net1078),
    .X(probe_env[0]));
 sky130_fd_sc_hd__buf_4 output444 (.A(net444),
    .X(probe_env[1]));
 sky130_fd_sc_hd__buf_4 output445 (.A(net445),
    .X(probe_jtagInstruction[0]));
 sky130_fd_sc_hd__buf_4 output446 (.A(net446),
    .X(probe_jtagInstruction[1]));
 sky130_fd_sc_hd__buf_4 output447 (.A(net447),
    .X(probe_jtagInstruction[2]));
 sky130_fd_sc_hd__buf_4 output448 (.A(net448),
    .X(probe_jtagInstruction[3]));
 sky130_fd_sc_hd__buf_4 output449 (.A(net449),
    .X(probe_jtagInstruction[4]));
 sky130_fd_sc_hd__buf_4 output450 (.A(net450),
    .X(probe_programCounter[0]));
 sky130_fd_sc_hd__buf_4 output451 (.A(net451),
    .X(probe_programCounter[10]));
 sky130_fd_sc_hd__buf_4 output452 (.A(net452),
    .X(probe_programCounter[11]));
 sky130_fd_sc_hd__buf_4 output453 (.A(net453),
    .X(probe_programCounter[12]));
 sky130_fd_sc_hd__buf_4 output454 (.A(net454),
    .X(probe_programCounter[13]));
 sky130_fd_sc_hd__buf_4 output455 (.A(net455),
    .X(probe_programCounter[14]));
 sky130_fd_sc_hd__buf_4 output456 (.A(net456),
    .X(probe_programCounter[15]));
 sky130_fd_sc_hd__buf_4 output457 (.A(net457),
    .X(probe_programCounter[16]));
 sky130_fd_sc_hd__buf_4 output458 (.A(net458),
    .X(probe_programCounter[17]));
 sky130_fd_sc_hd__buf_4 output459 (.A(net459),
    .X(probe_programCounter[18]));
 sky130_fd_sc_hd__buf_4 output460 (.A(net460),
    .X(probe_programCounter[19]));
 sky130_fd_sc_hd__buf_4 output461 (.A(net461),
    .X(probe_programCounter[1]));
 sky130_fd_sc_hd__buf_4 output462 (.A(net462),
    .X(probe_programCounter[20]));
 sky130_fd_sc_hd__buf_4 output463 (.A(net463),
    .X(probe_programCounter[21]));
 sky130_fd_sc_hd__buf_4 output464 (.A(net464),
    .X(probe_programCounter[22]));
 sky130_fd_sc_hd__buf_4 output465 (.A(net465),
    .X(probe_programCounter[23]));
 sky130_fd_sc_hd__buf_4 output466 (.A(net466),
    .X(probe_programCounter[24]));
 sky130_fd_sc_hd__buf_4 output467 (.A(net467),
    .X(probe_programCounter[25]));
 sky130_fd_sc_hd__buf_4 output468 (.A(net468),
    .X(probe_programCounter[26]));
 sky130_fd_sc_hd__buf_4 output469 (.A(net469),
    .X(probe_programCounter[27]));
 sky130_fd_sc_hd__buf_4 output470 (.A(net470),
    .X(probe_programCounter[28]));
 sky130_fd_sc_hd__buf_4 output471 (.A(net471),
    .X(probe_programCounter[29]));
 sky130_fd_sc_hd__buf_4 output472 (.A(net472),
    .X(probe_programCounter[2]));
 sky130_fd_sc_hd__buf_4 output473 (.A(net473),
    .X(probe_programCounter[30]));
 sky130_fd_sc_hd__buf_4 output474 (.A(net474),
    .X(probe_programCounter[31]));
 sky130_fd_sc_hd__buf_4 output475 (.A(net475),
    .X(probe_programCounter[3]));
 sky130_fd_sc_hd__buf_4 output476 (.A(net476),
    .X(probe_programCounter[4]));
 sky130_fd_sc_hd__buf_4 output477 (.A(net477),
    .X(probe_programCounter[5]));
 sky130_fd_sc_hd__buf_4 output478 (.A(net478),
    .X(probe_programCounter[6]));
 sky130_fd_sc_hd__buf_4 output479 (.A(net479),
    .X(probe_programCounter[7]));
 sky130_fd_sc_hd__buf_4 output480 (.A(net480),
    .X(probe_programCounter[8]));
 sky130_fd_sc_hd__buf_4 output481 (.A(net481),
    .X(probe_programCounter[9]));
 sky130_fd_sc_hd__buf_4 output482 (.A(net1776),
    .X(probe_state));
 sky130_fd_sc_hd__buf_4 output483 (.A(net483),
    .X(web0));
 sky130_fd_sc_hd__buf_6 output484 (.A(net484),
    .X(wmask0[0]));
 sky130_fd_sc_hd__buf_6 output485 (.A(net485),
    .X(wmask0[1]));
 sky130_fd_sc_hd__buf_6 output486 (.A(net486),
    .X(wmask0[2]));
 sky130_fd_sc_hd__buf_6 output487 (.A(net487),
    .X(wmask0[3]));
 sky130_fd_sc_hd__buf_2 rebuffer5 (.A(_06321_),
    .X(net2012));
 sky130_fd_sc_hd__clkbuf_4 split1 (.A(net702),
    .X(net2008));
 sky130_fd_sc_hd__clkbuf_4 split2 (.A(net712),
    .X(net2009));
 sky130_fd_sc_hd__buf_4 split3 (.A(net724),
    .X(net2010));
 sky130_fd_sc_hd__buf_2 split4 (.A(net973),
    .X(net2011));
 sky130_fd_sc_hd__clkbuf_4 split6 (.A(net794),
    .X(net2013));
 sky130_fd_sc_hd__clkbuf_4 split7 (.A(net1236),
    .X(net2014));
 sky130_fd_sc_hd__clkbuf_4 split8 (.A(net799),
    .X(net2015));
 sky130_fd_sc_hd__clkbuf_2 split9 (.A(net693),
    .X(net2016));
 sky130_fd_sc_hd__buf_12 wire1254 (.A(_08374_),
    .X(net1254));
 assign localMemory_wb_error_o = net2007;
endmodule

