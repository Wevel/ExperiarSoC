VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ExperiarCore
  CLASS BLOCK ;
  FOREIGN ExperiarCore ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 900.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END addr0[8]
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.080 4.000 580.680 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END addr1[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END clk0
  PIN clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END clk1
  PIN coreIndex[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 896.000 5.890 900.000 ;
    END
  END coreIndex[0]
  PIN coreIndex[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 896.000 17.390 900.000 ;
    END
  END coreIndex[1]
  PIN coreIndex[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 896.000 28.890 900.000 ;
    END
  END coreIndex[2]
  PIN coreIndex[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 896.000 40.390 900.000 ;
    END
  END coreIndex[3]
  PIN coreIndex[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 896.000 51.890 900.000 ;
    END
  END coreIndex[4]
  PIN coreIndex[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 896.000 63.390 900.000 ;
    END
  END coreIndex[5]
  PIN coreIndex[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 896.000 74.890 900.000 ;
    END
  END coreIndex[6]
  PIN coreIndex[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 896.000 86.390 900.000 ;
    END
  END coreIndex[7]
  PIN core_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 10.920 450.000 11.520 ;
    END
  END core_wb_ack_i
  PIN core_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 37.440 450.000 38.040 ;
    END
  END core_wb_adr_o[0]
  PIN core_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 189.080 450.000 189.680 ;
    END
  END core_wb_adr_o[10]
  PIN core_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 202.000 450.000 202.600 ;
    END
  END core_wb_adr_o[11]
  PIN core_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 215.600 450.000 216.200 ;
    END
  END core_wb_adr_o[12]
  PIN core_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 229.200 450.000 229.800 ;
    END
  END core_wb_adr_o[13]
  PIN core_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 242.120 450.000 242.720 ;
    END
  END core_wb_adr_o[14]
  PIN core_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 255.720 450.000 256.320 ;
    END
  END core_wb_adr_o[15]
  PIN core_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 269.320 450.000 269.920 ;
    END
  END core_wb_adr_o[16]
  PIN core_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 282.240 450.000 282.840 ;
    END
  END core_wb_adr_o[17]
  PIN core_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 295.840 450.000 296.440 ;
    END
  END core_wb_adr_o[18]
  PIN core_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 309.440 450.000 310.040 ;
    END
  END core_wb_adr_o[19]
  PIN core_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 55.120 450.000 55.720 ;
    END
  END core_wb_adr_o[1]
  PIN core_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 322.360 450.000 322.960 ;
    END
  END core_wb_adr_o[20]
  PIN core_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 335.960 450.000 336.560 ;
    END
  END core_wb_adr_o[21]
  PIN core_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 349.560 450.000 350.160 ;
    END
  END core_wb_adr_o[22]
  PIN core_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 362.480 450.000 363.080 ;
    END
  END core_wb_adr_o[23]
  PIN core_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 376.080 450.000 376.680 ;
    END
  END core_wb_adr_o[24]
  PIN core_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 389.680 450.000 390.280 ;
    END
  END core_wb_adr_o[25]
  PIN core_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 402.600 450.000 403.200 ;
    END
  END core_wb_adr_o[26]
  PIN core_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 416.200 450.000 416.800 ;
    END
  END core_wb_adr_o[27]
  PIN core_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 72.800 450.000 73.400 ;
    END
  END core_wb_adr_o[2]
  PIN core_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 91.160 450.000 91.760 ;
    END
  END core_wb_adr_o[3]
  PIN core_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 108.840 450.000 109.440 ;
    END
  END core_wb_adr_o[4]
  PIN core_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 121.760 450.000 122.360 ;
    END
  END core_wb_adr_o[5]
  PIN core_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 135.360 450.000 135.960 ;
    END
  END core_wb_adr_o[6]
  PIN core_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 148.960 450.000 149.560 ;
    END
  END core_wb_adr_o[7]
  PIN core_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 161.880 450.000 162.480 ;
    END
  END core_wb_adr_o[8]
  PIN core_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 175.480 450.000 176.080 ;
    END
  END core_wb_adr_o[9]
  PIN core_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 15.000 450.000 15.600 ;
    END
  END core_wb_cyc_o
  PIN core_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 41.520 450.000 42.120 ;
    END
  END core_wb_data_i[0]
  PIN core_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 193.160 450.000 193.760 ;
    END
  END core_wb_data_i[10]
  PIN core_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 206.760 450.000 207.360 ;
    END
  END core_wb_data_i[11]
  PIN core_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 220.360 450.000 220.960 ;
    END
  END core_wb_data_i[12]
  PIN core_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 233.280 450.000 233.880 ;
    END
  END core_wb_data_i[13]
  PIN core_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 246.880 450.000 247.480 ;
    END
  END core_wb_data_i[14]
  PIN core_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 260.480 450.000 261.080 ;
    END
  END core_wb_data_i[15]
  PIN core_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 273.400 450.000 274.000 ;
    END
  END core_wb_data_i[16]
  PIN core_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 287.000 450.000 287.600 ;
    END
  END core_wb_data_i[17]
  PIN core_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 300.600 450.000 301.200 ;
    END
  END core_wb_data_i[18]
  PIN core_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 313.520 450.000 314.120 ;
    END
  END core_wb_data_i[19]
  PIN core_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 59.880 450.000 60.480 ;
    END
  END core_wb_data_i[1]
  PIN core_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 327.120 450.000 327.720 ;
    END
  END core_wb_data_i[20]
  PIN core_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 340.720 450.000 341.320 ;
    END
  END core_wb_data_i[21]
  PIN core_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 353.640 450.000 354.240 ;
    END
  END core_wb_data_i[22]
  PIN core_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 367.240 450.000 367.840 ;
    END
  END core_wb_data_i[23]
  PIN core_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 380.840 450.000 381.440 ;
    END
  END core_wb_data_i[24]
  PIN core_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 393.760 450.000 394.360 ;
    END
  END core_wb_data_i[25]
  PIN core_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 407.360 450.000 407.960 ;
    END
  END core_wb_data_i[26]
  PIN core_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 420.960 450.000 421.560 ;
    END
  END core_wb_data_i[27]
  PIN core_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 429.800 450.000 430.400 ;
    END
  END core_wb_data_i[28]
  PIN core_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 438.640 450.000 439.240 ;
    END
  END core_wb_data_i[29]
  PIN core_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 77.560 450.000 78.160 ;
    END
  END core_wb_data_i[2]
  PIN core_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 447.480 450.000 448.080 ;
    END
  END core_wb_data_i[30]
  PIN core_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 456.320 450.000 456.920 ;
    END
  END core_wb_data_i[31]
  PIN core_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 95.240 450.000 95.840 ;
    END
  END core_wb_data_i[3]
  PIN core_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 112.920 450.000 113.520 ;
    END
  END core_wb_data_i[4]
  PIN core_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 126.520 450.000 127.120 ;
    END
  END core_wb_data_i[5]
  PIN core_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 140.120 450.000 140.720 ;
    END
  END core_wb_data_i[6]
  PIN core_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 153.040 450.000 153.640 ;
    END
  END core_wb_data_i[7]
  PIN core_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 166.640 450.000 167.240 ;
    END
  END core_wb_data_i[8]
  PIN core_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 180.240 450.000 180.840 ;
    END
  END core_wb_data_i[9]
  PIN core_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 46.280 450.000 46.880 ;
    END
  END core_wb_data_o[0]
  PIN core_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 197.920 450.000 198.520 ;
    END
  END core_wb_data_o[10]
  PIN core_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 211.520 450.000 212.120 ;
    END
  END core_wb_data_o[11]
  PIN core_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 224.440 450.000 225.040 ;
    END
  END core_wb_data_o[12]
  PIN core_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 238.040 450.000 238.640 ;
    END
  END core_wb_data_o[13]
  PIN core_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 251.640 450.000 252.240 ;
    END
  END core_wb_data_o[14]
  PIN core_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 264.560 450.000 265.160 ;
    END
  END core_wb_data_o[15]
  PIN core_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 278.160 450.000 278.760 ;
    END
  END core_wb_data_o[16]
  PIN core_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 291.760 450.000 292.360 ;
    END
  END core_wb_data_o[17]
  PIN core_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 304.680 450.000 305.280 ;
    END
  END core_wb_data_o[18]
  PIN core_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 318.280 450.000 318.880 ;
    END
  END core_wb_data_o[19]
  PIN core_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 63.960 450.000 64.560 ;
    END
  END core_wb_data_o[1]
  PIN core_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 331.880 450.000 332.480 ;
    END
  END core_wb_data_o[20]
  PIN core_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 344.800 450.000 345.400 ;
    END
  END core_wb_data_o[21]
  PIN core_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 358.400 450.000 359.000 ;
    END
  END core_wb_data_o[22]
  PIN core_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 372.000 450.000 372.600 ;
    END
  END core_wb_data_o[23]
  PIN core_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 384.920 450.000 385.520 ;
    END
  END core_wb_data_o[24]
  PIN core_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 398.520 450.000 399.120 ;
    END
  END core_wb_data_o[25]
  PIN core_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 412.120 450.000 412.720 ;
    END
  END core_wb_data_o[26]
  PIN core_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 425.040 450.000 425.640 ;
    END
  END core_wb_data_o[27]
  PIN core_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 433.880 450.000 434.480 ;
    END
  END core_wb_data_o[28]
  PIN core_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 442.720 450.000 443.320 ;
    END
  END core_wb_data_o[29]
  PIN core_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 81.640 450.000 82.240 ;
    END
  END core_wb_data_o[2]
  PIN core_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 452.240 450.000 452.840 ;
    END
  END core_wb_data_o[30]
  PIN core_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 461.080 450.000 461.680 ;
    END
  END core_wb_data_o[31]
  PIN core_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 100.000 450.000 100.600 ;
    END
  END core_wb_data_o[3]
  PIN core_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 117.680 450.000 118.280 ;
    END
  END core_wb_data_o[4]
  PIN core_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 131.280 450.000 131.880 ;
    END
  END core_wb_data_o[5]
  PIN core_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 144.200 450.000 144.800 ;
    END
  END core_wb_data_o[6]
  PIN core_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 157.800 450.000 158.400 ;
    END
  END core_wb_data_o[7]
  PIN core_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 171.400 450.000 172.000 ;
    END
  END core_wb_data_o[8]
  PIN core_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 184.320 450.000 184.920 ;
    END
  END core_wb_data_o[9]
  PIN core_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 19.760 450.000 20.360 ;
    END
  END core_wb_error_i
  PIN core_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 51.040 450.000 51.640 ;
    END
  END core_wb_sel_o[0]
  PIN core_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 68.720 450.000 69.320 ;
    END
  END core_wb_sel_o[1]
  PIN core_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 86.400 450.000 87.000 ;
    END
  END core_wb_sel_o[2]
  PIN core_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 104.080 450.000 104.680 ;
    END
  END core_wb_sel_o[3]
  PIN core_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 23.840 450.000 24.440 ;
    END
  END core_wb_stall_i
  PIN core_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 28.600 450.000 29.200 ;
    END
  END core_wb_stb_o
  PIN core_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 32.680 450.000 33.280 ;
    END
  END core_wb_we_o
  PIN csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END csb0[0]
  PIN csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END csb0[1]
  PIN csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END csb1[0]
  PIN csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END csb1[1]
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END din0[9]
  PIN dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END dout0[32]
  PIN dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END dout0[33]
  PIN dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END dout0[34]
  PIN dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END dout0[35]
  PIN dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 4.000 417.480 ;
    END
  END dout0[36]
  PIN dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END dout0[37]
  PIN dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END dout0[38]
  PIN dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END dout0[39]
  PIN dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END dout0[3]
  PIN dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END dout0[40]
  PIN dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END dout0[41]
  PIN dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END dout0[42]
  PIN dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END dout0[43]
  PIN dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END dout0[44]
  PIN dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END dout0[45]
  PIN dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END dout0[46]
  PIN dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END dout0[47]
  PIN dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END dout0[48]
  PIN dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END dout0[49]
  PIN dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END dout0[4]
  PIN dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END dout0[50]
  PIN dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END dout0[51]
  PIN dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 4.000 492.280 ;
    END
  END dout0[52]
  PIN dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END dout0[53]
  PIN dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END dout0[54]
  PIN dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 4.000 505.880 ;
    END
  END dout0[55]
  PIN dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END dout0[56]
  PIN dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END dout0[57]
  PIN dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END dout0[58]
  PIN dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END dout0[59]
  PIN dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END dout0[5]
  PIN dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END dout0[60]
  PIN dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END dout0[61]
  PIN dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END dout0[62]
  PIN dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END dout0[63]
  PIN dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.880 4.000 655.480 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.520 4.000 688.120 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.280 4.000 692.880 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END dout1[31]
  PIN dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.800 4.000 753.400 ;
    END
  END dout1[32]
  PIN dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END dout1[33]
  PIN dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 762.320 4.000 762.920 ;
    END
  END dout1[34]
  PIN dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 767.080 4.000 767.680 ;
    END
  END dout1[35]
  PIN dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.160 4.000 771.760 ;
    END
  END dout1[36]
  PIN dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.920 4.000 776.520 ;
    END
  END dout1[37]
  PIN dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END dout1[38]
  PIN dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END dout1[39]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END dout1[3]
  PIN dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.200 4.000 790.800 ;
    END
  END dout1[40]
  PIN dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.960 4.000 795.560 ;
    END
  END dout1[41]
  PIN dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.720 4.000 800.320 ;
    END
  END dout1[42]
  PIN dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.800 4.000 804.400 ;
    END
  END dout1[43]
  PIN dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 808.560 4.000 809.160 ;
    END
  END dout1[44]
  PIN dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END dout1[45]
  PIN dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END dout1[46]
  PIN dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END dout1[47]
  PIN dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 827.600 4.000 828.200 ;
    END
  END dout1[48]
  PIN dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END dout1[49]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END dout1[4]
  PIN dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END dout1[50]
  PIN dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.200 4.000 841.800 ;
    END
  END dout1[51]
  PIN dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.960 4.000 846.560 ;
    END
  END dout1[52]
  PIN dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.720 4.000 851.320 ;
    END
  END dout1[53]
  PIN dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END dout1[54]
  PIN dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END dout1[55]
  PIN dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END dout1[56]
  PIN dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 869.080 4.000 869.680 ;
    END
  END dout1[57]
  PIN dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END dout1[58]
  PIN dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END dout1[59]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END dout1[5]
  PIN dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 883.360 4.000 883.960 ;
    END
  END dout1[60]
  PIN dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END dout1[61]
  PIN dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.880 4.000 893.480 ;
    END
  END dout1[62]
  PIN dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END dout1[63]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 645.360 4.000 645.960 ;
    END
  END dout1[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END jtag_tms
  PIN localMemory_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 465.160 450.000 465.760 ;
    END
  END localMemory_wb_ack_o
  PIN localMemory_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 491.680 450.000 492.280 ;
    END
  END localMemory_wb_adr_i[0]
  PIN localMemory_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 643.320 450.000 643.920 ;
    END
  END localMemory_wb_adr_i[10]
  PIN localMemory_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 656.920 450.000 657.520 ;
    END
  END localMemory_wb_adr_i[11]
  PIN localMemory_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 670.520 450.000 671.120 ;
    END
  END localMemory_wb_adr_i[12]
  PIN localMemory_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 683.440 450.000 684.040 ;
    END
  END localMemory_wb_adr_i[13]
  PIN localMemory_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 697.040 450.000 697.640 ;
    END
  END localMemory_wb_adr_i[14]
  PIN localMemory_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 710.640 450.000 711.240 ;
    END
  END localMemory_wb_adr_i[15]
  PIN localMemory_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 723.560 450.000 724.160 ;
    END
  END localMemory_wb_adr_i[16]
  PIN localMemory_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 737.160 450.000 737.760 ;
    END
  END localMemory_wb_adr_i[17]
  PIN localMemory_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 750.760 450.000 751.360 ;
    END
  END localMemory_wb_adr_i[18]
  PIN localMemory_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 763.680 450.000 764.280 ;
    END
  END localMemory_wb_adr_i[19]
  PIN localMemory_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 510.040 450.000 510.640 ;
    END
  END localMemory_wb_adr_i[1]
  PIN localMemory_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 777.280 450.000 777.880 ;
    END
  END localMemory_wb_adr_i[20]
  PIN localMemory_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 790.880 450.000 791.480 ;
    END
  END localMemory_wb_adr_i[21]
  PIN localMemory_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 803.800 450.000 804.400 ;
    END
  END localMemory_wb_adr_i[22]
  PIN localMemory_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 817.400 450.000 818.000 ;
    END
  END localMemory_wb_adr_i[23]
  PIN localMemory_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 527.720 450.000 528.320 ;
    END
  END localMemory_wb_adr_i[2]
  PIN localMemory_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 545.400 450.000 546.000 ;
    END
  END localMemory_wb_adr_i[3]
  PIN localMemory_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 563.080 450.000 563.680 ;
    END
  END localMemory_wb_adr_i[4]
  PIN localMemory_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 576.680 450.000 577.280 ;
    END
  END localMemory_wb_adr_i[5]
  PIN localMemory_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 590.280 450.000 590.880 ;
    END
  END localMemory_wb_adr_i[6]
  PIN localMemory_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 603.200 450.000 603.800 ;
    END
  END localMemory_wb_adr_i[7]
  PIN localMemory_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 616.800 450.000 617.400 ;
    END
  END localMemory_wb_adr_i[8]
  PIN localMemory_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 630.400 450.000 631.000 ;
    END
  END localMemory_wb_adr_i[9]
  PIN localMemory_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 469.920 450.000 470.520 ;
    END
  END localMemory_wb_cyc_i
  PIN localMemory_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 496.440 450.000 497.040 ;
    END
  END localMemory_wb_data_i[0]
  PIN localMemory_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 648.080 450.000 648.680 ;
    END
  END localMemory_wb_data_i[10]
  PIN localMemory_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 661.680 450.000 662.280 ;
    END
  END localMemory_wb_data_i[11]
  PIN localMemory_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 674.600 450.000 675.200 ;
    END
  END localMemory_wb_data_i[12]
  PIN localMemory_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 688.200 450.000 688.800 ;
    END
  END localMemory_wb_data_i[13]
  PIN localMemory_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 701.800 450.000 702.400 ;
    END
  END localMemory_wb_data_i[14]
  PIN localMemory_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 714.720 450.000 715.320 ;
    END
  END localMemory_wb_data_i[15]
  PIN localMemory_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 728.320 450.000 728.920 ;
    END
  END localMemory_wb_data_i[16]
  PIN localMemory_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 741.920 450.000 742.520 ;
    END
  END localMemory_wb_data_i[17]
  PIN localMemory_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 754.840 450.000 755.440 ;
    END
  END localMemory_wb_data_i[18]
  PIN localMemory_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 768.440 450.000 769.040 ;
    END
  END localMemory_wb_data_i[19]
  PIN localMemory_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 514.120 450.000 514.720 ;
    END
  END localMemory_wb_data_i[1]
  PIN localMemory_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 782.040 450.000 782.640 ;
    END
  END localMemory_wb_data_i[20]
  PIN localMemory_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 794.960 450.000 795.560 ;
    END
  END localMemory_wb_data_i[21]
  PIN localMemory_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 808.560 450.000 809.160 ;
    END
  END localMemory_wb_data_i[22]
  PIN localMemory_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 822.160 450.000 822.760 ;
    END
  END localMemory_wb_data_i[23]
  PIN localMemory_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 831.000 450.000 831.600 ;
    END
  END localMemory_wb_data_i[24]
  PIN localMemory_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 839.840 450.000 840.440 ;
    END
  END localMemory_wb_data_i[25]
  PIN localMemory_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 848.680 450.000 849.280 ;
    END
  END localMemory_wb_data_i[26]
  PIN localMemory_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 857.520 450.000 858.120 ;
    END
  END localMemory_wb_data_i[27]
  PIN localMemory_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 866.360 450.000 866.960 ;
    END
  END localMemory_wb_data_i[28]
  PIN localMemory_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 875.200 450.000 875.800 ;
    END
  END localMemory_wb_data_i[29]
  PIN localMemory_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 531.800 450.000 532.400 ;
    END
  END localMemory_wb_data_i[2]
  PIN localMemory_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 884.040 450.000 884.640 ;
    END
  END localMemory_wb_data_i[30]
  PIN localMemory_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 892.880 450.000 893.480 ;
    END
  END localMemory_wb_data_i[31]
  PIN localMemory_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 550.160 450.000 550.760 ;
    END
  END localMemory_wb_data_i[3]
  PIN localMemory_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 567.840 450.000 568.440 ;
    END
  END localMemory_wb_data_i[4]
  PIN localMemory_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 581.440 450.000 582.040 ;
    END
  END localMemory_wb_data_i[5]
  PIN localMemory_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 594.360 450.000 594.960 ;
    END
  END localMemory_wb_data_i[6]
  PIN localMemory_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 607.960 450.000 608.560 ;
    END
  END localMemory_wb_data_i[7]
  PIN localMemory_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 621.560 450.000 622.160 ;
    END
  END localMemory_wb_data_i[8]
  PIN localMemory_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 634.480 450.000 635.080 ;
    END
  END localMemory_wb_data_i[9]
  PIN localMemory_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 501.200 450.000 501.800 ;
    END
  END localMemory_wb_data_o[0]
  PIN localMemory_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 652.160 450.000 652.760 ;
    END
  END localMemory_wb_data_o[10]
  PIN localMemory_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 665.760 450.000 666.360 ;
    END
  END localMemory_wb_data_o[11]
  PIN localMemory_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 679.360 450.000 679.960 ;
    END
  END localMemory_wb_data_o[12]
  PIN localMemory_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 692.280 450.000 692.880 ;
    END
  END localMemory_wb_data_o[13]
  PIN localMemory_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 705.880 450.000 706.480 ;
    END
  END localMemory_wb_data_o[14]
  PIN localMemory_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 719.480 450.000 720.080 ;
    END
  END localMemory_wb_data_o[15]
  PIN localMemory_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 732.400 450.000 733.000 ;
    END
  END localMemory_wb_data_o[16]
  PIN localMemory_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 746.000 450.000 746.600 ;
    END
  END localMemory_wb_data_o[17]
  PIN localMemory_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 759.600 450.000 760.200 ;
    END
  END localMemory_wb_data_o[18]
  PIN localMemory_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 772.520 450.000 773.120 ;
    END
  END localMemory_wb_data_o[19]
  PIN localMemory_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 518.880 450.000 519.480 ;
    END
  END localMemory_wb_data_o[1]
  PIN localMemory_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 786.120 450.000 786.720 ;
    END
  END localMemory_wb_data_o[20]
  PIN localMemory_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 799.720 450.000 800.320 ;
    END
  END localMemory_wb_data_o[21]
  PIN localMemory_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 812.640 450.000 813.240 ;
    END
  END localMemory_wb_data_o[22]
  PIN localMemory_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 826.240 450.000 826.840 ;
    END
  END localMemory_wb_data_o[23]
  PIN localMemory_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 835.080 450.000 835.680 ;
    END
  END localMemory_wb_data_o[24]
  PIN localMemory_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 843.920 450.000 844.520 ;
    END
  END localMemory_wb_data_o[25]
  PIN localMemory_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 852.760 450.000 853.360 ;
    END
  END localMemory_wb_data_o[26]
  PIN localMemory_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 862.280 450.000 862.880 ;
    END
  END localMemory_wb_data_o[27]
  PIN localMemory_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 871.120 450.000 871.720 ;
    END
  END localMemory_wb_data_o[28]
  PIN localMemory_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 879.960 450.000 880.560 ;
    END
  END localMemory_wb_data_o[29]
  PIN localMemory_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 536.560 450.000 537.160 ;
    END
  END localMemory_wb_data_o[2]
  PIN localMemory_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 888.800 450.000 889.400 ;
    END
  END localMemory_wb_data_o[30]
  PIN localMemory_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 897.640 450.000 898.240 ;
    END
  END localMemory_wb_data_o[31]
  PIN localMemory_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 554.240 450.000 554.840 ;
    END
  END localMemory_wb_data_o[3]
  PIN localMemory_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 571.920 450.000 572.520 ;
    END
  END localMemory_wb_data_o[4]
  PIN localMemory_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 585.520 450.000 586.120 ;
    END
  END localMemory_wb_data_o[5]
  PIN localMemory_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 599.120 450.000 599.720 ;
    END
  END localMemory_wb_data_o[6]
  PIN localMemory_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 612.040 450.000 612.640 ;
    END
  END localMemory_wb_data_o[7]
  PIN localMemory_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 625.640 450.000 626.240 ;
    END
  END localMemory_wb_data_o[8]
  PIN localMemory_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 639.240 450.000 639.840 ;
    END
  END localMemory_wb_data_o[9]
  PIN localMemory_wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 474.000 450.000 474.600 ;
    END
  END localMemory_wb_error_o
  PIN localMemory_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 505.280 450.000 505.880 ;
    END
  END localMemory_wb_sel_i[0]
  PIN localMemory_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 522.960 450.000 523.560 ;
    END
  END localMemory_wb_sel_i[1]
  PIN localMemory_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 541.320 450.000 541.920 ;
    END
  END localMemory_wb_sel_i[2]
  PIN localMemory_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 559.000 450.000 559.600 ;
    END
  END localMemory_wb_sel_i[3]
  PIN localMemory_wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 478.760 450.000 479.360 ;
    END
  END localMemory_wb_stall_o
  PIN localMemory_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 482.840 450.000 483.440 ;
    END
  END localMemory_wb_stb_i
  PIN localMemory_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 487.600 450.000 488.200 ;
    END
  END localMemory_wb_we_i
  PIN manufacturerID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 896.000 97.890 900.000 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 896.000 213.350 900.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 896.000 109.390 900.000 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 896.000 120.890 900.000 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 896.000 132.390 900.000 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 896.000 143.890 900.000 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 896.000 155.850 900.000 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 896.000 167.350 900.000 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 896.000 178.850 900.000 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 896.000 190.350 900.000 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 896.000 201.850 900.000 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 896.000 224.850 900.000 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 896.000 340.310 900.000 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 896.000 351.810 900.000 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 896.000 363.310 900.000 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 896.000 374.810 900.000 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 896.000 386.310 900.000 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 896.000 397.810 900.000 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 896.000 236.350 900.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 896.000 247.850 900.000 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 896.000 259.350 900.000 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 896.000 270.850 900.000 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 896.000 282.350 900.000 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 896.000 293.850 900.000 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 896.000 305.810 900.000 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 896.000 317.310 900.000 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 896.000 328.810 900.000 ;
    END
  END partID[9]
  PIN probe_errorCode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END probe_errorCode[0]
  PIN probe_errorCode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END probe_errorCode[1]
  PIN probe_errorCode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END probe_errorCode[2]
  PIN probe_errorCode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END probe_errorCode[3]
  PIN probe_isBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END probe_isBranch
  PIN probe_isCompressed
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END probe_isCompressed
  PIN probe_isLoad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END probe_isLoad
  PIN probe_isStore
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END probe_isStore
  PIN probe_jtagInstruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END probe_jtagInstruction[0]
  PIN probe_jtagInstruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END probe_jtagInstruction[1]
  PIN probe_jtagInstruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END probe_jtagInstruction[2]
  PIN probe_jtagInstruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END probe_jtagInstruction[3]
  PIN probe_jtagInstruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END probe_jtagInstruction[4]
  PIN probe_opcode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END probe_opcode[0]
  PIN probe_opcode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END probe_opcode[1]
  PIN probe_opcode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END probe_opcode[2]
  PIN probe_opcode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END probe_opcode[3]
  PIN probe_opcode[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END probe_opcode[4]
  PIN probe_opcode[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END probe_opcode[5]
  PIN probe_opcode[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END probe_opcode[6]
  PIN probe_programCounter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END probe_programCounter[0]
  PIN probe_programCounter[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END probe_programCounter[10]
  PIN probe_programCounter[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END probe_programCounter[11]
  PIN probe_programCounter[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END probe_programCounter[12]
  PIN probe_programCounter[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END probe_programCounter[13]
  PIN probe_programCounter[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END probe_programCounter[14]
  PIN probe_programCounter[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END probe_programCounter[15]
  PIN probe_programCounter[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END probe_programCounter[16]
  PIN probe_programCounter[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END probe_programCounter[17]
  PIN probe_programCounter[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END probe_programCounter[18]
  PIN probe_programCounter[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END probe_programCounter[19]
  PIN probe_programCounter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END probe_programCounter[1]
  PIN probe_programCounter[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END probe_programCounter[20]
  PIN probe_programCounter[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END probe_programCounter[21]
  PIN probe_programCounter[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END probe_programCounter[22]
  PIN probe_programCounter[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END probe_programCounter[23]
  PIN probe_programCounter[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END probe_programCounter[24]
  PIN probe_programCounter[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END probe_programCounter[25]
  PIN probe_programCounter[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END probe_programCounter[26]
  PIN probe_programCounter[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END probe_programCounter[27]
  PIN probe_programCounter[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END probe_programCounter[28]
  PIN probe_programCounter[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END probe_programCounter[29]
  PIN probe_programCounter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END probe_programCounter[2]
  PIN probe_programCounter[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END probe_programCounter[30]
  PIN probe_programCounter[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END probe_programCounter[31]
  PIN probe_programCounter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END probe_programCounter[3]
  PIN probe_programCounter[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END probe_programCounter[4]
  PIN probe_programCounter[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END probe_programCounter[5]
  PIN probe_programCounter[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END probe_programCounter[6]
  PIN probe_programCounter[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END probe_programCounter[7]
  PIN probe_programCounter[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END probe_programCounter[8]
  PIN probe_programCounter[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END probe_programCounter[9]
  PIN probe_state[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END probe_state[0]
  PIN probe_state[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END probe_state[1]
  PIN probe_takeBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END probe_takeBranch
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 886.960 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 896.000 409.310 900.000 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 896.000 420.810 900.000 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 896.000 432.310 900.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 896.000 443.810 900.000 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 886.960 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 2.080 450.000 2.680 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 6.160 450.000 6.760 ;
    END
  END wb_rst_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 444.360 886.805 ;
      LAYER met1 ;
        RECT 0.070 6.500 449.810 890.420 ;
      LAYER met2 ;
        RECT 0.100 895.720 5.330 898.125 ;
        RECT 6.170 895.720 16.830 898.125 ;
        RECT 17.670 895.720 28.330 898.125 ;
        RECT 29.170 895.720 39.830 898.125 ;
        RECT 40.670 895.720 51.330 898.125 ;
        RECT 52.170 895.720 62.830 898.125 ;
        RECT 63.670 895.720 74.330 898.125 ;
        RECT 75.170 895.720 85.830 898.125 ;
        RECT 86.670 895.720 97.330 898.125 ;
        RECT 98.170 895.720 108.830 898.125 ;
        RECT 109.670 895.720 120.330 898.125 ;
        RECT 121.170 895.720 131.830 898.125 ;
        RECT 132.670 895.720 143.330 898.125 ;
        RECT 144.170 895.720 155.290 898.125 ;
        RECT 156.130 895.720 166.790 898.125 ;
        RECT 167.630 895.720 178.290 898.125 ;
        RECT 179.130 895.720 189.790 898.125 ;
        RECT 190.630 895.720 201.290 898.125 ;
        RECT 202.130 895.720 212.790 898.125 ;
        RECT 213.630 895.720 224.290 898.125 ;
        RECT 225.130 895.720 235.790 898.125 ;
        RECT 236.630 895.720 247.290 898.125 ;
        RECT 248.130 895.720 258.790 898.125 ;
        RECT 259.630 895.720 270.290 898.125 ;
        RECT 271.130 895.720 281.790 898.125 ;
        RECT 282.630 895.720 293.290 898.125 ;
        RECT 294.130 895.720 305.250 898.125 ;
        RECT 306.090 895.720 316.750 898.125 ;
        RECT 317.590 895.720 328.250 898.125 ;
        RECT 329.090 895.720 339.750 898.125 ;
        RECT 340.590 895.720 351.250 898.125 ;
        RECT 352.090 895.720 362.750 898.125 ;
        RECT 363.590 895.720 374.250 898.125 ;
        RECT 375.090 895.720 385.750 898.125 ;
        RECT 386.590 895.720 397.250 898.125 ;
        RECT 398.090 895.720 408.750 898.125 ;
        RECT 409.590 895.720 420.250 898.125 ;
        RECT 421.090 895.720 431.750 898.125 ;
        RECT 432.590 895.720 443.250 898.125 ;
        RECT 444.090 895.720 449.790 898.125 ;
        RECT 0.100 4.280 449.790 895.720 ;
        RECT 0.100 2.195 3.490 4.280 ;
        RECT 4.330 2.195 11.310 4.280 ;
        RECT 12.150 2.195 19.590 4.280 ;
        RECT 20.430 2.195 27.870 4.280 ;
        RECT 28.710 2.195 36.150 4.280 ;
        RECT 36.990 2.195 43.970 4.280 ;
        RECT 44.810 2.195 52.250 4.280 ;
        RECT 53.090 2.195 60.530 4.280 ;
        RECT 61.370 2.195 68.810 4.280 ;
        RECT 69.650 2.195 77.090 4.280 ;
        RECT 77.930 2.195 84.910 4.280 ;
        RECT 85.750 2.195 93.190 4.280 ;
        RECT 94.030 2.195 101.470 4.280 ;
        RECT 102.310 2.195 109.750 4.280 ;
        RECT 110.590 2.195 117.570 4.280 ;
        RECT 118.410 2.195 125.850 4.280 ;
        RECT 126.690 2.195 134.130 4.280 ;
        RECT 134.970 2.195 142.410 4.280 ;
        RECT 143.250 2.195 150.690 4.280 ;
        RECT 151.530 2.195 158.510 4.280 ;
        RECT 159.350 2.195 166.790 4.280 ;
        RECT 167.630 2.195 175.070 4.280 ;
        RECT 175.910 2.195 183.350 4.280 ;
        RECT 184.190 2.195 191.170 4.280 ;
        RECT 192.010 2.195 199.450 4.280 ;
        RECT 200.290 2.195 207.730 4.280 ;
        RECT 208.570 2.195 216.010 4.280 ;
        RECT 216.850 2.195 224.290 4.280 ;
        RECT 225.130 2.195 232.110 4.280 ;
        RECT 232.950 2.195 240.390 4.280 ;
        RECT 241.230 2.195 248.670 4.280 ;
        RECT 249.510 2.195 256.950 4.280 ;
        RECT 257.790 2.195 265.230 4.280 ;
        RECT 266.070 2.195 273.050 4.280 ;
        RECT 273.890 2.195 281.330 4.280 ;
        RECT 282.170 2.195 289.610 4.280 ;
        RECT 290.450 2.195 297.890 4.280 ;
        RECT 298.730 2.195 305.710 4.280 ;
        RECT 306.550 2.195 313.990 4.280 ;
        RECT 314.830 2.195 322.270 4.280 ;
        RECT 323.110 2.195 330.550 4.280 ;
        RECT 331.390 2.195 338.830 4.280 ;
        RECT 339.670 2.195 346.650 4.280 ;
        RECT 347.490 2.195 354.930 4.280 ;
        RECT 355.770 2.195 363.210 4.280 ;
        RECT 364.050 2.195 371.490 4.280 ;
        RECT 372.330 2.195 379.310 4.280 ;
        RECT 380.150 2.195 387.590 4.280 ;
        RECT 388.430 2.195 395.870 4.280 ;
        RECT 396.710 2.195 404.150 4.280 ;
        RECT 404.990 2.195 412.430 4.280 ;
        RECT 413.270 2.195 420.250 4.280 ;
        RECT 421.090 2.195 428.530 4.280 ;
        RECT 429.370 2.195 436.810 4.280 ;
        RECT 437.650 2.195 445.090 4.280 ;
        RECT 445.930 2.195 449.790 4.280 ;
      LAYER met3 ;
        RECT 4.400 897.240 445.600 898.105 ;
        RECT 0.270 893.880 449.815 897.240 ;
        RECT 4.400 892.480 445.600 893.880 ;
        RECT 0.270 889.800 449.815 892.480 ;
        RECT 0.270 889.120 445.600 889.800 ;
        RECT 4.400 888.400 445.600 889.120 ;
        RECT 4.400 887.720 449.815 888.400 ;
        RECT 0.270 885.040 449.815 887.720 ;
        RECT 0.270 884.360 445.600 885.040 ;
        RECT 4.400 883.640 445.600 884.360 ;
        RECT 4.400 882.960 449.815 883.640 ;
        RECT 0.270 880.960 449.815 882.960 ;
        RECT 0.270 879.600 445.600 880.960 ;
        RECT 4.400 879.560 445.600 879.600 ;
        RECT 4.400 878.200 449.815 879.560 ;
        RECT 0.270 876.200 449.815 878.200 ;
        RECT 0.270 874.840 445.600 876.200 ;
        RECT 4.400 874.800 445.600 874.840 ;
        RECT 4.400 873.440 449.815 874.800 ;
        RECT 0.270 872.120 449.815 873.440 ;
        RECT 0.270 870.720 445.600 872.120 ;
        RECT 0.270 870.080 449.815 870.720 ;
        RECT 4.400 868.680 449.815 870.080 ;
        RECT 0.270 867.360 449.815 868.680 ;
        RECT 0.270 866.000 445.600 867.360 ;
        RECT 4.400 865.960 445.600 866.000 ;
        RECT 4.400 864.600 449.815 865.960 ;
        RECT 0.270 863.280 449.815 864.600 ;
        RECT 0.270 861.880 445.600 863.280 ;
        RECT 0.270 861.240 449.815 861.880 ;
        RECT 4.400 859.840 449.815 861.240 ;
        RECT 0.270 858.520 449.815 859.840 ;
        RECT 0.270 857.120 445.600 858.520 ;
        RECT 0.270 856.480 449.815 857.120 ;
        RECT 4.400 855.080 449.815 856.480 ;
        RECT 0.270 853.760 449.815 855.080 ;
        RECT 0.270 852.360 445.600 853.760 ;
        RECT 0.270 851.720 449.815 852.360 ;
        RECT 4.400 850.320 449.815 851.720 ;
        RECT 0.270 849.680 449.815 850.320 ;
        RECT 0.270 848.280 445.600 849.680 ;
        RECT 0.270 846.960 449.815 848.280 ;
        RECT 4.400 845.560 449.815 846.960 ;
        RECT 0.270 844.920 449.815 845.560 ;
        RECT 0.270 843.520 445.600 844.920 ;
        RECT 0.270 842.200 449.815 843.520 ;
        RECT 4.400 840.840 449.815 842.200 ;
        RECT 4.400 840.800 445.600 840.840 ;
        RECT 0.270 839.440 445.600 840.800 ;
        RECT 0.270 837.440 449.815 839.440 ;
        RECT 4.400 836.080 449.815 837.440 ;
        RECT 4.400 836.040 445.600 836.080 ;
        RECT 0.270 834.680 445.600 836.040 ;
        RECT 0.270 833.360 449.815 834.680 ;
        RECT 4.400 832.000 449.815 833.360 ;
        RECT 4.400 831.960 445.600 832.000 ;
        RECT 0.270 830.600 445.600 831.960 ;
        RECT 0.270 828.600 449.815 830.600 ;
        RECT 4.400 827.240 449.815 828.600 ;
        RECT 4.400 827.200 445.600 827.240 ;
        RECT 0.270 825.840 445.600 827.200 ;
        RECT 0.270 823.840 449.815 825.840 ;
        RECT 4.400 823.160 449.815 823.840 ;
        RECT 4.400 822.440 445.600 823.160 ;
        RECT 0.270 821.760 445.600 822.440 ;
        RECT 0.270 819.080 449.815 821.760 ;
        RECT 4.400 818.400 449.815 819.080 ;
        RECT 4.400 817.680 445.600 818.400 ;
        RECT 0.270 817.000 445.600 817.680 ;
        RECT 0.270 814.320 449.815 817.000 ;
        RECT 4.400 813.640 449.815 814.320 ;
        RECT 4.400 812.920 445.600 813.640 ;
        RECT 0.270 812.240 445.600 812.920 ;
        RECT 0.270 809.560 449.815 812.240 ;
        RECT 4.400 808.160 445.600 809.560 ;
        RECT 0.270 804.800 449.815 808.160 ;
        RECT 4.400 803.400 445.600 804.800 ;
        RECT 0.270 800.720 449.815 803.400 ;
        RECT 4.400 799.320 445.600 800.720 ;
        RECT 0.270 795.960 449.815 799.320 ;
        RECT 4.400 794.560 445.600 795.960 ;
        RECT 0.270 791.880 449.815 794.560 ;
        RECT 0.270 791.200 445.600 791.880 ;
        RECT 4.400 790.480 445.600 791.200 ;
        RECT 4.400 789.800 449.815 790.480 ;
        RECT 0.270 787.120 449.815 789.800 ;
        RECT 0.270 786.440 445.600 787.120 ;
        RECT 4.400 785.720 445.600 786.440 ;
        RECT 4.400 785.040 449.815 785.720 ;
        RECT 0.270 783.040 449.815 785.040 ;
        RECT 0.270 781.680 445.600 783.040 ;
        RECT 4.400 781.640 445.600 781.680 ;
        RECT 4.400 780.280 449.815 781.640 ;
        RECT 0.270 778.280 449.815 780.280 ;
        RECT 0.270 776.920 445.600 778.280 ;
        RECT 4.400 776.880 445.600 776.920 ;
        RECT 4.400 775.520 449.815 776.880 ;
        RECT 0.270 773.520 449.815 775.520 ;
        RECT 0.270 772.160 445.600 773.520 ;
        RECT 4.400 772.120 445.600 772.160 ;
        RECT 4.400 770.760 449.815 772.120 ;
        RECT 0.270 769.440 449.815 770.760 ;
        RECT 0.270 768.080 445.600 769.440 ;
        RECT 4.400 768.040 445.600 768.080 ;
        RECT 4.400 766.680 449.815 768.040 ;
        RECT 0.270 764.680 449.815 766.680 ;
        RECT 0.270 763.320 445.600 764.680 ;
        RECT 4.400 763.280 445.600 763.320 ;
        RECT 4.400 761.920 449.815 763.280 ;
        RECT 0.270 760.600 449.815 761.920 ;
        RECT 0.270 759.200 445.600 760.600 ;
        RECT 0.270 758.560 449.815 759.200 ;
        RECT 4.400 757.160 449.815 758.560 ;
        RECT 0.270 755.840 449.815 757.160 ;
        RECT 0.270 754.440 445.600 755.840 ;
        RECT 0.270 753.800 449.815 754.440 ;
        RECT 4.400 752.400 449.815 753.800 ;
        RECT 0.270 751.760 449.815 752.400 ;
        RECT 0.270 750.360 445.600 751.760 ;
        RECT 0.270 749.040 449.815 750.360 ;
        RECT 4.400 747.640 449.815 749.040 ;
        RECT 0.270 747.000 449.815 747.640 ;
        RECT 0.270 745.600 445.600 747.000 ;
        RECT 0.270 744.280 449.815 745.600 ;
        RECT 4.400 742.920 449.815 744.280 ;
        RECT 4.400 742.880 445.600 742.920 ;
        RECT 0.270 741.520 445.600 742.880 ;
        RECT 0.270 739.520 449.815 741.520 ;
        RECT 4.400 738.160 449.815 739.520 ;
        RECT 4.400 738.120 445.600 738.160 ;
        RECT 0.270 736.760 445.600 738.120 ;
        RECT 0.270 735.440 449.815 736.760 ;
        RECT 4.400 734.040 449.815 735.440 ;
        RECT 0.270 733.400 449.815 734.040 ;
        RECT 0.270 732.000 445.600 733.400 ;
        RECT 0.270 730.680 449.815 732.000 ;
        RECT 4.400 729.320 449.815 730.680 ;
        RECT 4.400 729.280 445.600 729.320 ;
        RECT 0.270 727.920 445.600 729.280 ;
        RECT 0.270 725.920 449.815 727.920 ;
        RECT 4.400 724.560 449.815 725.920 ;
        RECT 4.400 724.520 445.600 724.560 ;
        RECT 0.270 723.160 445.600 724.520 ;
        RECT 0.270 721.160 449.815 723.160 ;
        RECT 4.400 720.480 449.815 721.160 ;
        RECT 4.400 719.760 445.600 720.480 ;
        RECT 0.270 719.080 445.600 719.760 ;
        RECT 0.270 716.400 449.815 719.080 ;
        RECT 4.400 715.720 449.815 716.400 ;
        RECT 4.400 715.000 445.600 715.720 ;
        RECT 0.270 714.320 445.600 715.000 ;
        RECT 0.270 711.640 449.815 714.320 ;
        RECT 4.400 710.240 445.600 711.640 ;
        RECT 0.270 706.880 449.815 710.240 ;
        RECT 4.400 705.480 445.600 706.880 ;
        RECT 0.270 702.800 449.815 705.480 ;
        RECT 4.400 701.400 445.600 702.800 ;
        RECT 0.270 698.040 449.815 701.400 ;
        RECT 4.400 696.640 445.600 698.040 ;
        RECT 0.270 693.280 449.815 696.640 ;
        RECT 4.400 691.880 445.600 693.280 ;
        RECT 0.270 689.200 449.815 691.880 ;
        RECT 0.270 688.520 445.600 689.200 ;
        RECT 4.400 687.800 445.600 688.520 ;
        RECT 4.400 687.120 449.815 687.800 ;
        RECT 0.270 684.440 449.815 687.120 ;
        RECT 0.270 683.760 445.600 684.440 ;
        RECT 4.400 683.040 445.600 683.760 ;
        RECT 4.400 682.360 449.815 683.040 ;
        RECT 0.270 680.360 449.815 682.360 ;
        RECT 0.270 679.000 445.600 680.360 ;
        RECT 4.400 678.960 445.600 679.000 ;
        RECT 4.400 677.600 449.815 678.960 ;
        RECT 0.270 675.600 449.815 677.600 ;
        RECT 0.270 674.240 445.600 675.600 ;
        RECT 4.400 674.200 445.600 674.240 ;
        RECT 4.400 672.840 449.815 674.200 ;
        RECT 0.270 671.520 449.815 672.840 ;
        RECT 0.270 670.120 445.600 671.520 ;
        RECT 0.270 669.480 449.815 670.120 ;
        RECT 4.400 668.080 449.815 669.480 ;
        RECT 0.270 666.760 449.815 668.080 ;
        RECT 0.270 665.400 445.600 666.760 ;
        RECT 4.400 665.360 445.600 665.400 ;
        RECT 4.400 664.000 449.815 665.360 ;
        RECT 0.270 662.680 449.815 664.000 ;
        RECT 0.270 661.280 445.600 662.680 ;
        RECT 0.270 660.640 449.815 661.280 ;
        RECT 4.400 659.240 449.815 660.640 ;
        RECT 0.270 657.920 449.815 659.240 ;
        RECT 0.270 656.520 445.600 657.920 ;
        RECT 0.270 655.880 449.815 656.520 ;
        RECT 4.400 654.480 449.815 655.880 ;
        RECT 0.270 653.160 449.815 654.480 ;
        RECT 0.270 651.760 445.600 653.160 ;
        RECT 0.270 651.120 449.815 651.760 ;
        RECT 4.400 649.720 449.815 651.120 ;
        RECT 0.270 649.080 449.815 649.720 ;
        RECT 0.270 647.680 445.600 649.080 ;
        RECT 0.270 646.360 449.815 647.680 ;
        RECT 4.400 644.960 449.815 646.360 ;
        RECT 0.270 644.320 449.815 644.960 ;
        RECT 0.270 642.920 445.600 644.320 ;
        RECT 0.270 641.600 449.815 642.920 ;
        RECT 4.400 640.240 449.815 641.600 ;
        RECT 4.400 640.200 445.600 640.240 ;
        RECT 0.270 638.840 445.600 640.200 ;
        RECT 0.270 636.840 449.815 638.840 ;
        RECT 4.400 635.480 449.815 636.840 ;
        RECT 4.400 635.440 445.600 635.480 ;
        RECT 0.270 634.080 445.600 635.440 ;
        RECT 0.270 632.760 449.815 634.080 ;
        RECT 4.400 631.400 449.815 632.760 ;
        RECT 4.400 631.360 445.600 631.400 ;
        RECT 0.270 630.000 445.600 631.360 ;
        RECT 0.270 628.000 449.815 630.000 ;
        RECT 4.400 626.640 449.815 628.000 ;
        RECT 4.400 626.600 445.600 626.640 ;
        RECT 0.270 625.240 445.600 626.600 ;
        RECT 0.270 623.240 449.815 625.240 ;
        RECT 4.400 622.560 449.815 623.240 ;
        RECT 4.400 621.840 445.600 622.560 ;
        RECT 0.270 621.160 445.600 621.840 ;
        RECT 0.270 618.480 449.815 621.160 ;
        RECT 4.400 617.800 449.815 618.480 ;
        RECT 4.400 617.080 445.600 617.800 ;
        RECT 0.270 616.400 445.600 617.080 ;
        RECT 0.270 613.720 449.815 616.400 ;
        RECT 4.400 613.040 449.815 613.720 ;
        RECT 4.400 612.320 445.600 613.040 ;
        RECT 0.270 611.640 445.600 612.320 ;
        RECT 0.270 608.960 449.815 611.640 ;
        RECT 4.400 607.560 445.600 608.960 ;
        RECT 0.270 604.200 449.815 607.560 ;
        RECT 4.400 602.800 445.600 604.200 ;
        RECT 0.270 600.120 449.815 602.800 ;
        RECT 4.400 598.720 445.600 600.120 ;
        RECT 0.270 595.360 449.815 598.720 ;
        RECT 4.400 593.960 445.600 595.360 ;
        RECT 0.270 591.280 449.815 593.960 ;
        RECT 0.270 590.600 445.600 591.280 ;
        RECT 4.400 589.880 445.600 590.600 ;
        RECT 4.400 589.200 449.815 589.880 ;
        RECT 0.270 586.520 449.815 589.200 ;
        RECT 0.270 585.840 445.600 586.520 ;
        RECT 4.400 585.120 445.600 585.840 ;
        RECT 4.400 584.440 449.815 585.120 ;
        RECT 0.270 582.440 449.815 584.440 ;
        RECT 0.270 581.080 445.600 582.440 ;
        RECT 4.400 581.040 445.600 581.080 ;
        RECT 4.400 579.680 449.815 581.040 ;
        RECT 0.270 577.680 449.815 579.680 ;
        RECT 0.270 576.320 445.600 577.680 ;
        RECT 4.400 576.280 445.600 576.320 ;
        RECT 4.400 574.920 449.815 576.280 ;
        RECT 0.270 572.920 449.815 574.920 ;
        RECT 0.270 571.560 445.600 572.920 ;
        RECT 4.400 571.520 445.600 571.560 ;
        RECT 4.400 570.160 449.815 571.520 ;
        RECT 0.270 568.840 449.815 570.160 ;
        RECT 0.270 567.480 445.600 568.840 ;
        RECT 4.400 567.440 445.600 567.480 ;
        RECT 4.400 566.080 449.815 567.440 ;
        RECT 0.270 564.080 449.815 566.080 ;
        RECT 0.270 562.720 445.600 564.080 ;
        RECT 4.400 562.680 445.600 562.720 ;
        RECT 4.400 561.320 449.815 562.680 ;
        RECT 0.270 560.000 449.815 561.320 ;
        RECT 0.270 558.600 445.600 560.000 ;
        RECT 0.270 557.960 449.815 558.600 ;
        RECT 4.400 556.560 449.815 557.960 ;
        RECT 0.270 555.240 449.815 556.560 ;
        RECT 0.270 553.840 445.600 555.240 ;
        RECT 0.270 553.200 449.815 553.840 ;
        RECT 4.400 551.800 449.815 553.200 ;
        RECT 0.270 551.160 449.815 551.800 ;
        RECT 0.270 549.760 445.600 551.160 ;
        RECT 0.270 548.440 449.815 549.760 ;
        RECT 4.400 547.040 449.815 548.440 ;
        RECT 0.270 546.400 449.815 547.040 ;
        RECT 0.270 545.000 445.600 546.400 ;
        RECT 0.270 543.680 449.815 545.000 ;
        RECT 4.400 542.320 449.815 543.680 ;
        RECT 4.400 542.280 445.600 542.320 ;
        RECT 0.270 540.920 445.600 542.280 ;
        RECT 0.270 538.920 449.815 540.920 ;
        RECT 4.400 537.560 449.815 538.920 ;
        RECT 4.400 537.520 445.600 537.560 ;
        RECT 0.270 536.160 445.600 537.520 ;
        RECT 0.270 534.840 449.815 536.160 ;
        RECT 4.400 533.440 449.815 534.840 ;
        RECT 0.270 532.800 449.815 533.440 ;
        RECT 0.270 531.400 445.600 532.800 ;
        RECT 0.270 530.080 449.815 531.400 ;
        RECT 4.400 528.720 449.815 530.080 ;
        RECT 4.400 528.680 445.600 528.720 ;
        RECT 0.270 527.320 445.600 528.680 ;
        RECT 0.270 525.320 449.815 527.320 ;
        RECT 4.400 523.960 449.815 525.320 ;
        RECT 4.400 523.920 445.600 523.960 ;
        RECT 0.270 522.560 445.600 523.920 ;
        RECT 0.270 520.560 449.815 522.560 ;
        RECT 4.400 519.880 449.815 520.560 ;
        RECT 4.400 519.160 445.600 519.880 ;
        RECT 0.270 518.480 445.600 519.160 ;
        RECT 0.270 515.800 449.815 518.480 ;
        RECT 4.400 515.120 449.815 515.800 ;
        RECT 4.400 514.400 445.600 515.120 ;
        RECT 0.270 513.720 445.600 514.400 ;
        RECT 0.270 511.040 449.815 513.720 ;
        RECT 4.400 509.640 445.600 511.040 ;
        RECT 0.270 506.280 449.815 509.640 ;
        RECT 4.400 504.880 445.600 506.280 ;
        RECT 0.270 502.200 449.815 504.880 ;
        RECT 4.400 500.800 445.600 502.200 ;
        RECT 0.270 497.440 449.815 500.800 ;
        RECT 4.400 496.040 445.600 497.440 ;
        RECT 0.270 492.680 449.815 496.040 ;
        RECT 4.400 491.280 445.600 492.680 ;
        RECT 0.270 488.600 449.815 491.280 ;
        RECT 0.270 487.920 445.600 488.600 ;
        RECT 4.400 487.200 445.600 487.920 ;
        RECT 4.400 486.520 449.815 487.200 ;
        RECT 0.270 483.840 449.815 486.520 ;
        RECT 0.270 483.160 445.600 483.840 ;
        RECT 4.400 482.440 445.600 483.160 ;
        RECT 4.400 481.760 449.815 482.440 ;
        RECT 0.270 479.760 449.815 481.760 ;
        RECT 0.270 478.400 445.600 479.760 ;
        RECT 4.400 478.360 445.600 478.400 ;
        RECT 4.400 477.000 449.815 478.360 ;
        RECT 0.270 475.000 449.815 477.000 ;
        RECT 0.270 473.640 445.600 475.000 ;
        RECT 4.400 473.600 445.600 473.640 ;
        RECT 4.400 472.240 449.815 473.600 ;
        RECT 0.270 470.920 449.815 472.240 ;
        RECT 0.270 469.560 445.600 470.920 ;
        RECT 4.400 469.520 445.600 469.560 ;
        RECT 4.400 468.160 449.815 469.520 ;
        RECT 0.270 466.160 449.815 468.160 ;
        RECT 0.270 464.800 445.600 466.160 ;
        RECT 4.400 464.760 445.600 464.800 ;
        RECT 4.400 463.400 449.815 464.760 ;
        RECT 0.270 462.080 449.815 463.400 ;
        RECT 0.270 460.680 445.600 462.080 ;
        RECT 0.270 460.040 449.815 460.680 ;
        RECT 4.400 458.640 449.815 460.040 ;
        RECT 0.270 457.320 449.815 458.640 ;
        RECT 0.270 455.920 445.600 457.320 ;
        RECT 0.270 455.280 449.815 455.920 ;
        RECT 4.400 453.880 449.815 455.280 ;
        RECT 0.270 453.240 449.815 453.880 ;
        RECT 0.270 451.840 445.600 453.240 ;
        RECT 0.270 450.520 449.815 451.840 ;
        RECT 4.400 449.120 449.815 450.520 ;
        RECT 0.270 448.480 449.815 449.120 ;
        RECT 0.270 447.080 445.600 448.480 ;
        RECT 0.270 445.760 449.815 447.080 ;
        RECT 4.400 444.360 449.815 445.760 ;
        RECT 0.270 443.720 449.815 444.360 ;
        RECT 0.270 442.320 445.600 443.720 ;
        RECT 0.270 441.000 449.815 442.320 ;
        RECT 4.400 439.640 449.815 441.000 ;
        RECT 4.400 439.600 445.600 439.640 ;
        RECT 0.270 438.240 445.600 439.600 ;
        RECT 0.270 436.240 449.815 438.240 ;
        RECT 4.400 434.880 449.815 436.240 ;
        RECT 4.400 434.840 445.600 434.880 ;
        RECT 0.270 433.480 445.600 434.840 ;
        RECT 0.270 432.160 449.815 433.480 ;
        RECT 4.400 430.800 449.815 432.160 ;
        RECT 4.400 430.760 445.600 430.800 ;
        RECT 0.270 429.400 445.600 430.760 ;
        RECT 0.270 427.400 449.815 429.400 ;
        RECT 4.400 426.040 449.815 427.400 ;
        RECT 4.400 426.000 445.600 426.040 ;
        RECT 0.270 424.640 445.600 426.000 ;
        RECT 0.270 422.640 449.815 424.640 ;
        RECT 4.400 421.960 449.815 422.640 ;
        RECT 4.400 421.240 445.600 421.960 ;
        RECT 0.270 420.560 445.600 421.240 ;
        RECT 0.270 417.880 449.815 420.560 ;
        RECT 4.400 417.200 449.815 417.880 ;
        RECT 4.400 416.480 445.600 417.200 ;
        RECT 0.270 415.800 445.600 416.480 ;
        RECT 0.270 413.120 449.815 415.800 ;
        RECT 4.400 411.720 445.600 413.120 ;
        RECT 0.270 408.360 449.815 411.720 ;
        RECT 4.400 406.960 445.600 408.360 ;
        RECT 0.270 403.600 449.815 406.960 ;
        RECT 4.400 402.200 445.600 403.600 ;
        RECT 0.270 399.520 449.815 402.200 ;
        RECT 4.400 398.120 445.600 399.520 ;
        RECT 0.270 394.760 449.815 398.120 ;
        RECT 4.400 393.360 445.600 394.760 ;
        RECT 0.270 390.680 449.815 393.360 ;
        RECT 0.270 390.000 445.600 390.680 ;
        RECT 4.400 389.280 445.600 390.000 ;
        RECT 4.400 388.600 449.815 389.280 ;
        RECT 0.270 385.920 449.815 388.600 ;
        RECT 0.270 385.240 445.600 385.920 ;
        RECT 4.400 384.520 445.600 385.240 ;
        RECT 4.400 383.840 449.815 384.520 ;
        RECT 0.270 381.840 449.815 383.840 ;
        RECT 0.270 380.480 445.600 381.840 ;
        RECT 4.400 380.440 445.600 380.480 ;
        RECT 4.400 379.080 449.815 380.440 ;
        RECT 0.270 377.080 449.815 379.080 ;
        RECT 0.270 375.720 445.600 377.080 ;
        RECT 4.400 375.680 445.600 375.720 ;
        RECT 4.400 374.320 449.815 375.680 ;
        RECT 0.270 373.000 449.815 374.320 ;
        RECT 0.270 371.600 445.600 373.000 ;
        RECT 0.270 370.960 449.815 371.600 ;
        RECT 4.400 369.560 449.815 370.960 ;
        RECT 0.270 368.240 449.815 369.560 ;
        RECT 0.270 366.880 445.600 368.240 ;
        RECT 4.400 366.840 445.600 366.880 ;
        RECT 4.400 365.480 449.815 366.840 ;
        RECT 0.270 363.480 449.815 365.480 ;
        RECT 0.270 362.120 445.600 363.480 ;
        RECT 4.400 362.080 445.600 362.120 ;
        RECT 4.400 360.720 449.815 362.080 ;
        RECT 0.270 359.400 449.815 360.720 ;
        RECT 0.270 358.000 445.600 359.400 ;
        RECT 0.270 357.360 449.815 358.000 ;
        RECT 4.400 355.960 449.815 357.360 ;
        RECT 0.270 354.640 449.815 355.960 ;
        RECT 0.270 353.240 445.600 354.640 ;
        RECT 0.270 352.600 449.815 353.240 ;
        RECT 4.400 351.200 449.815 352.600 ;
        RECT 0.270 350.560 449.815 351.200 ;
        RECT 0.270 349.160 445.600 350.560 ;
        RECT 0.270 347.840 449.815 349.160 ;
        RECT 4.400 346.440 449.815 347.840 ;
        RECT 0.270 345.800 449.815 346.440 ;
        RECT 0.270 344.400 445.600 345.800 ;
        RECT 0.270 343.080 449.815 344.400 ;
        RECT 4.400 341.720 449.815 343.080 ;
        RECT 4.400 341.680 445.600 341.720 ;
        RECT 0.270 340.320 445.600 341.680 ;
        RECT 0.270 338.320 449.815 340.320 ;
        RECT 4.400 336.960 449.815 338.320 ;
        RECT 4.400 336.920 445.600 336.960 ;
        RECT 0.270 335.560 445.600 336.920 ;
        RECT 0.270 334.240 449.815 335.560 ;
        RECT 4.400 332.880 449.815 334.240 ;
        RECT 4.400 332.840 445.600 332.880 ;
        RECT 0.270 331.480 445.600 332.840 ;
        RECT 0.270 329.480 449.815 331.480 ;
        RECT 4.400 328.120 449.815 329.480 ;
        RECT 4.400 328.080 445.600 328.120 ;
        RECT 0.270 326.720 445.600 328.080 ;
        RECT 0.270 324.720 449.815 326.720 ;
        RECT 4.400 323.360 449.815 324.720 ;
        RECT 4.400 323.320 445.600 323.360 ;
        RECT 0.270 321.960 445.600 323.320 ;
        RECT 0.270 319.960 449.815 321.960 ;
        RECT 4.400 319.280 449.815 319.960 ;
        RECT 4.400 318.560 445.600 319.280 ;
        RECT 0.270 317.880 445.600 318.560 ;
        RECT 0.270 315.200 449.815 317.880 ;
        RECT 4.400 314.520 449.815 315.200 ;
        RECT 4.400 313.800 445.600 314.520 ;
        RECT 0.270 313.120 445.600 313.800 ;
        RECT 0.270 310.440 449.815 313.120 ;
        RECT 4.400 309.040 445.600 310.440 ;
        RECT 0.270 305.680 449.815 309.040 ;
        RECT 4.400 304.280 445.600 305.680 ;
        RECT 0.270 301.600 449.815 304.280 ;
        RECT 4.400 300.200 445.600 301.600 ;
        RECT 0.270 296.840 449.815 300.200 ;
        RECT 4.400 295.440 445.600 296.840 ;
        RECT 0.270 292.760 449.815 295.440 ;
        RECT 0.270 292.080 445.600 292.760 ;
        RECT 4.400 291.360 445.600 292.080 ;
        RECT 4.400 290.680 449.815 291.360 ;
        RECT 0.270 288.000 449.815 290.680 ;
        RECT 0.270 287.320 445.600 288.000 ;
        RECT 4.400 286.600 445.600 287.320 ;
        RECT 4.400 285.920 449.815 286.600 ;
        RECT 0.270 283.240 449.815 285.920 ;
        RECT 0.270 282.560 445.600 283.240 ;
        RECT 4.400 281.840 445.600 282.560 ;
        RECT 4.400 281.160 449.815 281.840 ;
        RECT 0.270 279.160 449.815 281.160 ;
        RECT 0.270 277.800 445.600 279.160 ;
        RECT 4.400 277.760 445.600 277.800 ;
        RECT 4.400 276.400 449.815 277.760 ;
        RECT 0.270 274.400 449.815 276.400 ;
        RECT 0.270 273.040 445.600 274.400 ;
        RECT 4.400 273.000 445.600 273.040 ;
        RECT 4.400 271.640 449.815 273.000 ;
        RECT 0.270 270.320 449.815 271.640 ;
        RECT 0.270 268.960 445.600 270.320 ;
        RECT 4.400 268.920 445.600 268.960 ;
        RECT 4.400 267.560 449.815 268.920 ;
        RECT 0.270 265.560 449.815 267.560 ;
        RECT 0.270 264.200 445.600 265.560 ;
        RECT 4.400 264.160 445.600 264.200 ;
        RECT 4.400 262.800 449.815 264.160 ;
        RECT 0.270 261.480 449.815 262.800 ;
        RECT 0.270 260.080 445.600 261.480 ;
        RECT 0.270 259.440 449.815 260.080 ;
        RECT 4.400 258.040 449.815 259.440 ;
        RECT 0.270 256.720 449.815 258.040 ;
        RECT 0.270 255.320 445.600 256.720 ;
        RECT 0.270 254.680 449.815 255.320 ;
        RECT 4.400 253.280 449.815 254.680 ;
        RECT 0.270 252.640 449.815 253.280 ;
        RECT 0.270 251.240 445.600 252.640 ;
        RECT 0.270 249.920 449.815 251.240 ;
        RECT 4.400 248.520 449.815 249.920 ;
        RECT 0.270 247.880 449.815 248.520 ;
        RECT 0.270 246.480 445.600 247.880 ;
        RECT 0.270 245.160 449.815 246.480 ;
        RECT 4.400 243.760 449.815 245.160 ;
        RECT 0.270 243.120 449.815 243.760 ;
        RECT 0.270 241.720 445.600 243.120 ;
        RECT 0.270 240.400 449.815 241.720 ;
        RECT 4.400 239.040 449.815 240.400 ;
        RECT 4.400 239.000 445.600 239.040 ;
        RECT 0.270 237.640 445.600 239.000 ;
        RECT 0.270 236.320 449.815 237.640 ;
        RECT 4.400 234.920 449.815 236.320 ;
        RECT 0.270 234.280 449.815 234.920 ;
        RECT 0.270 232.880 445.600 234.280 ;
        RECT 0.270 231.560 449.815 232.880 ;
        RECT 4.400 230.200 449.815 231.560 ;
        RECT 4.400 230.160 445.600 230.200 ;
        RECT 0.270 228.800 445.600 230.160 ;
        RECT 0.270 226.800 449.815 228.800 ;
        RECT 4.400 225.440 449.815 226.800 ;
        RECT 4.400 225.400 445.600 225.440 ;
        RECT 0.270 224.040 445.600 225.400 ;
        RECT 0.270 222.040 449.815 224.040 ;
        RECT 4.400 221.360 449.815 222.040 ;
        RECT 4.400 220.640 445.600 221.360 ;
        RECT 0.270 219.960 445.600 220.640 ;
        RECT 0.270 217.280 449.815 219.960 ;
        RECT 4.400 216.600 449.815 217.280 ;
        RECT 4.400 215.880 445.600 216.600 ;
        RECT 0.270 215.200 445.600 215.880 ;
        RECT 0.270 212.520 449.815 215.200 ;
        RECT 4.400 211.120 445.600 212.520 ;
        RECT 0.270 207.760 449.815 211.120 ;
        RECT 4.400 206.360 445.600 207.760 ;
        RECT 0.270 203.000 449.815 206.360 ;
        RECT 4.400 201.600 445.600 203.000 ;
        RECT 0.270 198.920 449.815 201.600 ;
        RECT 4.400 197.520 445.600 198.920 ;
        RECT 0.270 194.160 449.815 197.520 ;
        RECT 4.400 192.760 445.600 194.160 ;
        RECT 0.270 190.080 449.815 192.760 ;
        RECT 0.270 189.400 445.600 190.080 ;
        RECT 4.400 188.680 445.600 189.400 ;
        RECT 4.400 188.000 449.815 188.680 ;
        RECT 0.270 185.320 449.815 188.000 ;
        RECT 0.270 184.640 445.600 185.320 ;
        RECT 4.400 183.920 445.600 184.640 ;
        RECT 4.400 183.240 449.815 183.920 ;
        RECT 0.270 181.240 449.815 183.240 ;
        RECT 0.270 179.880 445.600 181.240 ;
        RECT 4.400 179.840 445.600 179.880 ;
        RECT 4.400 178.480 449.815 179.840 ;
        RECT 0.270 176.480 449.815 178.480 ;
        RECT 0.270 175.120 445.600 176.480 ;
        RECT 4.400 175.080 445.600 175.120 ;
        RECT 4.400 173.720 449.815 175.080 ;
        RECT 0.270 172.400 449.815 173.720 ;
        RECT 0.270 171.000 445.600 172.400 ;
        RECT 0.270 170.360 449.815 171.000 ;
        RECT 4.400 168.960 449.815 170.360 ;
        RECT 0.270 167.640 449.815 168.960 ;
        RECT 0.270 166.280 445.600 167.640 ;
        RECT 4.400 166.240 445.600 166.280 ;
        RECT 4.400 164.880 449.815 166.240 ;
        RECT 0.270 162.880 449.815 164.880 ;
        RECT 0.270 161.520 445.600 162.880 ;
        RECT 4.400 161.480 445.600 161.520 ;
        RECT 4.400 160.120 449.815 161.480 ;
        RECT 0.270 158.800 449.815 160.120 ;
        RECT 0.270 157.400 445.600 158.800 ;
        RECT 0.270 156.760 449.815 157.400 ;
        RECT 4.400 155.360 449.815 156.760 ;
        RECT 0.270 154.040 449.815 155.360 ;
        RECT 0.270 152.640 445.600 154.040 ;
        RECT 0.270 152.000 449.815 152.640 ;
        RECT 4.400 150.600 449.815 152.000 ;
        RECT 0.270 149.960 449.815 150.600 ;
        RECT 0.270 148.560 445.600 149.960 ;
        RECT 0.270 147.240 449.815 148.560 ;
        RECT 4.400 145.840 449.815 147.240 ;
        RECT 0.270 145.200 449.815 145.840 ;
        RECT 0.270 143.800 445.600 145.200 ;
        RECT 0.270 142.480 449.815 143.800 ;
        RECT 4.400 141.120 449.815 142.480 ;
        RECT 4.400 141.080 445.600 141.120 ;
        RECT 0.270 139.720 445.600 141.080 ;
        RECT 0.270 137.720 449.815 139.720 ;
        RECT 4.400 136.360 449.815 137.720 ;
        RECT 4.400 136.320 445.600 136.360 ;
        RECT 0.270 134.960 445.600 136.320 ;
        RECT 0.270 133.640 449.815 134.960 ;
        RECT 4.400 132.280 449.815 133.640 ;
        RECT 4.400 132.240 445.600 132.280 ;
        RECT 0.270 130.880 445.600 132.240 ;
        RECT 0.270 128.880 449.815 130.880 ;
        RECT 4.400 127.520 449.815 128.880 ;
        RECT 4.400 127.480 445.600 127.520 ;
        RECT 0.270 126.120 445.600 127.480 ;
        RECT 0.270 124.120 449.815 126.120 ;
        RECT 4.400 122.760 449.815 124.120 ;
        RECT 4.400 122.720 445.600 122.760 ;
        RECT 0.270 121.360 445.600 122.720 ;
        RECT 0.270 119.360 449.815 121.360 ;
        RECT 4.400 118.680 449.815 119.360 ;
        RECT 4.400 117.960 445.600 118.680 ;
        RECT 0.270 117.280 445.600 117.960 ;
        RECT 0.270 114.600 449.815 117.280 ;
        RECT 4.400 113.920 449.815 114.600 ;
        RECT 4.400 113.200 445.600 113.920 ;
        RECT 0.270 112.520 445.600 113.200 ;
        RECT 0.270 109.840 449.815 112.520 ;
        RECT 4.400 108.440 445.600 109.840 ;
        RECT 0.270 105.080 449.815 108.440 ;
        RECT 4.400 103.680 445.600 105.080 ;
        RECT 0.270 101.000 449.815 103.680 ;
        RECT 4.400 99.600 445.600 101.000 ;
        RECT 0.270 96.240 449.815 99.600 ;
        RECT 4.400 94.840 445.600 96.240 ;
        RECT 0.270 92.160 449.815 94.840 ;
        RECT 0.270 91.480 445.600 92.160 ;
        RECT 4.400 90.760 445.600 91.480 ;
        RECT 4.400 90.080 449.815 90.760 ;
        RECT 0.270 87.400 449.815 90.080 ;
        RECT 0.270 86.720 445.600 87.400 ;
        RECT 4.400 86.000 445.600 86.720 ;
        RECT 4.400 85.320 449.815 86.000 ;
        RECT 0.270 82.640 449.815 85.320 ;
        RECT 0.270 81.960 445.600 82.640 ;
        RECT 4.400 81.240 445.600 81.960 ;
        RECT 4.400 80.560 449.815 81.240 ;
        RECT 0.270 78.560 449.815 80.560 ;
        RECT 0.270 77.200 445.600 78.560 ;
        RECT 4.400 77.160 445.600 77.200 ;
        RECT 4.400 75.800 449.815 77.160 ;
        RECT 0.270 73.800 449.815 75.800 ;
        RECT 0.270 72.440 445.600 73.800 ;
        RECT 4.400 72.400 445.600 72.440 ;
        RECT 4.400 71.040 449.815 72.400 ;
        RECT 0.270 69.720 449.815 71.040 ;
        RECT 0.270 68.360 445.600 69.720 ;
        RECT 4.400 68.320 445.600 68.360 ;
        RECT 4.400 66.960 449.815 68.320 ;
        RECT 0.270 64.960 449.815 66.960 ;
        RECT 0.270 63.600 445.600 64.960 ;
        RECT 4.400 63.560 445.600 63.600 ;
        RECT 4.400 62.200 449.815 63.560 ;
        RECT 0.270 60.880 449.815 62.200 ;
        RECT 0.270 59.480 445.600 60.880 ;
        RECT 0.270 58.840 449.815 59.480 ;
        RECT 4.400 57.440 449.815 58.840 ;
        RECT 0.270 56.120 449.815 57.440 ;
        RECT 0.270 54.720 445.600 56.120 ;
        RECT 0.270 54.080 449.815 54.720 ;
        RECT 4.400 52.680 449.815 54.080 ;
        RECT 0.270 52.040 449.815 52.680 ;
        RECT 0.270 50.640 445.600 52.040 ;
        RECT 0.270 49.320 449.815 50.640 ;
        RECT 4.400 47.920 449.815 49.320 ;
        RECT 0.270 47.280 449.815 47.920 ;
        RECT 0.270 45.880 445.600 47.280 ;
        RECT 0.270 44.560 449.815 45.880 ;
        RECT 4.400 43.160 449.815 44.560 ;
        RECT 0.270 42.520 449.815 43.160 ;
        RECT 0.270 41.120 445.600 42.520 ;
        RECT 0.270 39.800 449.815 41.120 ;
        RECT 4.400 38.440 449.815 39.800 ;
        RECT 4.400 38.400 445.600 38.440 ;
        RECT 0.270 37.040 445.600 38.400 ;
        RECT 0.270 35.720 449.815 37.040 ;
        RECT 4.400 34.320 449.815 35.720 ;
        RECT 0.270 33.680 449.815 34.320 ;
        RECT 0.270 32.280 445.600 33.680 ;
        RECT 0.270 30.960 449.815 32.280 ;
        RECT 4.400 29.600 449.815 30.960 ;
        RECT 4.400 29.560 445.600 29.600 ;
        RECT 0.270 28.200 445.600 29.560 ;
        RECT 0.270 26.200 449.815 28.200 ;
        RECT 4.400 24.840 449.815 26.200 ;
        RECT 4.400 24.800 445.600 24.840 ;
        RECT 0.270 23.440 445.600 24.800 ;
        RECT 0.270 21.440 449.815 23.440 ;
        RECT 4.400 20.760 449.815 21.440 ;
        RECT 4.400 20.040 445.600 20.760 ;
        RECT 0.270 19.360 445.600 20.040 ;
        RECT 0.270 16.680 449.815 19.360 ;
        RECT 4.400 16.000 449.815 16.680 ;
        RECT 4.400 15.280 445.600 16.000 ;
        RECT 0.270 14.600 445.600 15.280 ;
        RECT 0.270 11.920 449.815 14.600 ;
        RECT 4.400 10.520 445.600 11.920 ;
        RECT 0.270 7.160 449.815 10.520 ;
        RECT 4.400 5.760 445.600 7.160 ;
        RECT 0.270 3.080 449.815 5.760 ;
        RECT 4.400 2.215 445.600 3.080 ;
      LAYER met4 ;
        RECT 0.295 11.735 20.640 883.825 ;
        RECT 23.040 11.735 97.440 883.825 ;
        RECT 99.840 11.735 174.240 883.825 ;
        RECT 176.640 11.735 251.040 883.825 ;
        RECT 253.440 11.735 327.840 883.825 ;
        RECT 330.240 11.735 404.640 883.825 ;
        RECT 407.040 11.735 449.585 883.825 ;
  END
END ExperiarCore
END LIBRARY

