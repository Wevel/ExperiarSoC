magic
tech sky130A
magscale 1 2
timestamp 1653062708
<< obsli1 >>
rect 1104 2159 158884 97393
<< obsm1 >>
rect 382 1232 159514 98320
<< metal2 >>
rect 386 99200 442 100000
rect 1214 99200 1270 100000
rect 2042 99200 2098 100000
rect 2870 99200 2926 100000
rect 3790 99200 3846 100000
rect 4618 99200 4674 100000
rect 5446 99200 5502 100000
rect 6366 99200 6422 100000
rect 7194 99200 7250 100000
rect 8022 99200 8078 100000
rect 8850 99200 8906 100000
rect 9770 99200 9826 100000
rect 10598 99200 10654 100000
rect 11426 99200 11482 100000
rect 12346 99200 12402 100000
rect 13174 99200 13230 100000
rect 14002 99200 14058 100000
rect 14922 99200 14978 100000
rect 15750 99200 15806 100000
rect 16578 99200 16634 100000
rect 17406 99200 17462 100000
rect 18326 99200 18382 100000
rect 19154 99200 19210 100000
rect 19982 99200 20038 100000
rect 20902 99200 20958 100000
rect 21730 99200 21786 100000
rect 22558 99200 22614 100000
rect 23478 99200 23534 100000
rect 24306 99200 24362 100000
rect 25134 99200 25190 100000
rect 25962 99200 26018 100000
rect 26882 99200 26938 100000
rect 27710 99200 27766 100000
rect 28538 99200 28594 100000
rect 29458 99200 29514 100000
rect 30286 99200 30342 100000
rect 31114 99200 31170 100000
rect 32034 99200 32090 100000
rect 32862 99200 32918 100000
rect 33690 99200 33746 100000
rect 34518 99200 34574 100000
rect 35438 99200 35494 100000
rect 36266 99200 36322 100000
rect 37094 99200 37150 100000
rect 38014 99200 38070 100000
rect 38842 99200 38898 100000
rect 39670 99200 39726 100000
rect 40590 99200 40646 100000
rect 41418 99200 41474 100000
rect 42246 99200 42302 100000
rect 43074 99200 43130 100000
rect 43994 99200 44050 100000
rect 44822 99200 44878 100000
rect 45650 99200 45706 100000
rect 46570 99200 46626 100000
rect 47398 99200 47454 100000
rect 48226 99200 48282 100000
rect 49146 99200 49202 100000
rect 49974 99200 50030 100000
rect 50802 99200 50858 100000
rect 51630 99200 51686 100000
rect 52550 99200 52606 100000
rect 53378 99200 53434 100000
rect 54206 99200 54262 100000
rect 55126 99200 55182 100000
rect 55954 99200 56010 100000
rect 56782 99200 56838 100000
rect 57702 99200 57758 100000
rect 58530 99200 58586 100000
rect 59358 99200 59414 100000
rect 60186 99200 60242 100000
rect 61106 99200 61162 100000
rect 61934 99200 61990 100000
rect 62762 99200 62818 100000
rect 63682 99200 63738 100000
rect 64510 99200 64566 100000
rect 65338 99200 65394 100000
rect 66258 99200 66314 100000
rect 67086 99200 67142 100000
rect 67914 99200 67970 100000
rect 68742 99200 68798 100000
rect 69662 99200 69718 100000
rect 70490 99200 70546 100000
rect 71318 99200 71374 100000
rect 72238 99200 72294 100000
rect 73066 99200 73122 100000
rect 73894 99200 73950 100000
rect 74814 99200 74870 100000
rect 75642 99200 75698 100000
rect 76470 99200 76526 100000
rect 77298 99200 77354 100000
rect 78218 99200 78274 100000
rect 79046 99200 79102 100000
rect 79874 99200 79930 100000
rect 80794 99200 80850 100000
rect 81622 99200 81678 100000
rect 82450 99200 82506 100000
rect 83370 99200 83426 100000
rect 84198 99200 84254 100000
rect 85026 99200 85082 100000
rect 85854 99200 85910 100000
rect 86774 99200 86830 100000
rect 87602 99200 87658 100000
rect 88430 99200 88486 100000
rect 89350 99200 89406 100000
rect 90178 99200 90234 100000
rect 91006 99200 91062 100000
rect 91926 99200 91982 100000
rect 92754 99200 92810 100000
rect 93582 99200 93638 100000
rect 94410 99200 94466 100000
rect 95330 99200 95386 100000
rect 96158 99200 96214 100000
rect 96986 99200 97042 100000
rect 97906 99200 97962 100000
rect 98734 99200 98790 100000
rect 99562 99200 99618 100000
rect 100482 99200 100538 100000
rect 101310 99200 101366 100000
rect 102138 99200 102194 100000
rect 102966 99200 103022 100000
rect 103886 99200 103942 100000
rect 104714 99200 104770 100000
rect 105542 99200 105598 100000
rect 106462 99200 106518 100000
rect 107290 99200 107346 100000
rect 108118 99200 108174 100000
rect 109038 99200 109094 100000
rect 109866 99200 109922 100000
rect 110694 99200 110750 100000
rect 111522 99200 111578 100000
rect 112442 99200 112498 100000
rect 113270 99200 113326 100000
rect 114098 99200 114154 100000
rect 115018 99200 115074 100000
rect 115846 99200 115902 100000
rect 116674 99200 116730 100000
rect 117594 99200 117650 100000
rect 118422 99200 118478 100000
rect 119250 99200 119306 100000
rect 120078 99200 120134 100000
rect 120998 99200 121054 100000
rect 121826 99200 121882 100000
rect 122654 99200 122710 100000
rect 123574 99200 123630 100000
rect 124402 99200 124458 100000
rect 125230 99200 125286 100000
rect 126150 99200 126206 100000
rect 126978 99200 127034 100000
rect 127806 99200 127862 100000
rect 128634 99200 128690 100000
rect 129554 99200 129610 100000
rect 130382 99200 130438 100000
rect 131210 99200 131266 100000
rect 132130 99200 132186 100000
rect 132958 99200 133014 100000
rect 133786 99200 133842 100000
rect 134706 99200 134762 100000
rect 135534 99200 135590 100000
rect 136362 99200 136418 100000
rect 137190 99200 137246 100000
rect 138110 99200 138166 100000
rect 138938 99200 138994 100000
rect 139766 99200 139822 100000
rect 140686 99200 140742 100000
rect 141514 99200 141570 100000
rect 142342 99200 142398 100000
rect 143262 99200 143318 100000
rect 144090 99200 144146 100000
rect 144918 99200 144974 100000
rect 145746 99200 145802 100000
rect 146666 99200 146722 100000
rect 147494 99200 147550 100000
rect 148322 99200 148378 100000
rect 149242 99200 149298 100000
rect 150070 99200 150126 100000
rect 150898 99200 150954 100000
rect 151818 99200 151874 100000
rect 152646 99200 152702 100000
rect 153474 99200 153530 100000
rect 154302 99200 154358 100000
rect 155222 99200 155278 100000
rect 156050 99200 156106 100000
rect 156878 99200 156934 100000
rect 157798 99200 157854 100000
rect 158626 99200 158682 100000
rect 159454 99200 159510 100000
rect 1950 0 2006 800
rect 5814 0 5870 800
rect 9678 0 9734 800
rect 13634 0 13690 800
rect 17498 0 17554 800
rect 21454 0 21510 800
rect 25318 0 25374 800
rect 29182 0 29238 800
rect 33138 0 33194 800
rect 37002 0 37058 800
rect 40958 0 41014 800
rect 44822 0 44878 800
rect 48686 0 48742 800
rect 52642 0 52698 800
rect 56506 0 56562 800
rect 60462 0 60518 800
rect 64326 0 64382 800
rect 68282 0 68338 800
rect 72146 0 72202 800
rect 76010 0 76066 800
rect 79966 0 80022 800
rect 83830 0 83886 800
rect 87786 0 87842 800
rect 91650 0 91706 800
rect 95514 0 95570 800
rect 99470 0 99526 800
rect 103334 0 103390 800
rect 107290 0 107346 800
rect 111154 0 111210 800
rect 115110 0 115166 800
rect 118974 0 119030 800
rect 122838 0 122894 800
rect 126794 0 126850 800
rect 130658 0 130714 800
rect 134614 0 134670 800
rect 138478 0 138534 800
rect 142342 0 142398 800
rect 146298 0 146354 800
rect 150162 0 150218 800
rect 154118 0 154174 800
rect 157982 0 158038 800
<< obsm2 >>
rect 498 99144 1158 99657
rect 1326 99144 1986 99657
rect 2154 99144 2814 99657
rect 2982 99144 3734 99657
rect 3902 99144 4562 99657
rect 4730 99144 5390 99657
rect 5558 99144 6310 99657
rect 6478 99144 7138 99657
rect 7306 99144 7966 99657
rect 8134 99144 8794 99657
rect 8962 99144 9714 99657
rect 9882 99144 10542 99657
rect 10710 99144 11370 99657
rect 11538 99144 12290 99657
rect 12458 99144 13118 99657
rect 13286 99144 13946 99657
rect 14114 99144 14866 99657
rect 15034 99144 15694 99657
rect 15862 99144 16522 99657
rect 16690 99144 17350 99657
rect 17518 99144 18270 99657
rect 18438 99144 19098 99657
rect 19266 99144 19926 99657
rect 20094 99144 20846 99657
rect 21014 99144 21674 99657
rect 21842 99144 22502 99657
rect 22670 99144 23422 99657
rect 23590 99144 24250 99657
rect 24418 99144 25078 99657
rect 25246 99144 25906 99657
rect 26074 99144 26826 99657
rect 26994 99144 27654 99657
rect 27822 99144 28482 99657
rect 28650 99144 29402 99657
rect 29570 99144 30230 99657
rect 30398 99144 31058 99657
rect 31226 99144 31978 99657
rect 32146 99144 32806 99657
rect 32974 99144 33634 99657
rect 33802 99144 34462 99657
rect 34630 99144 35382 99657
rect 35550 99144 36210 99657
rect 36378 99144 37038 99657
rect 37206 99144 37958 99657
rect 38126 99144 38786 99657
rect 38954 99144 39614 99657
rect 39782 99144 40534 99657
rect 40702 99144 41362 99657
rect 41530 99144 42190 99657
rect 42358 99144 43018 99657
rect 43186 99144 43938 99657
rect 44106 99144 44766 99657
rect 44934 99144 45594 99657
rect 45762 99144 46514 99657
rect 46682 99144 47342 99657
rect 47510 99144 48170 99657
rect 48338 99144 49090 99657
rect 49258 99144 49918 99657
rect 50086 99144 50746 99657
rect 50914 99144 51574 99657
rect 51742 99144 52494 99657
rect 52662 99144 53322 99657
rect 53490 99144 54150 99657
rect 54318 99144 55070 99657
rect 55238 99144 55898 99657
rect 56066 99144 56726 99657
rect 56894 99144 57646 99657
rect 57814 99144 58474 99657
rect 58642 99144 59302 99657
rect 59470 99144 60130 99657
rect 60298 99144 61050 99657
rect 61218 99144 61878 99657
rect 62046 99144 62706 99657
rect 62874 99144 63626 99657
rect 63794 99144 64454 99657
rect 64622 99144 65282 99657
rect 65450 99144 66202 99657
rect 66370 99144 67030 99657
rect 67198 99144 67858 99657
rect 68026 99144 68686 99657
rect 68854 99144 69606 99657
rect 69774 99144 70434 99657
rect 70602 99144 71262 99657
rect 71430 99144 72182 99657
rect 72350 99144 73010 99657
rect 73178 99144 73838 99657
rect 74006 99144 74758 99657
rect 74926 99144 75586 99657
rect 75754 99144 76414 99657
rect 76582 99144 77242 99657
rect 77410 99144 78162 99657
rect 78330 99144 78990 99657
rect 79158 99144 79818 99657
rect 79986 99144 80738 99657
rect 80906 99144 81566 99657
rect 81734 99144 82394 99657
rect 82562 99144 83314 99657
rect 83482 99144 84142 99657
rect 84310 99144 84970 99657
rect 85138 99144 85798 99657
rect 85966 99144 86718 99657
rect 86886 99144 87546 99657
rect 87714 99144 88374 99657
rect 88542 99144 89294 99657
rect 89462 99144 90122 99657
rect 90290 99144 90950 99657
rect 91118 99144 91870 99657
rect 92038 99144 92698 99657
rect 92866 99144 93526 99657
rect 93694 99144 94354 99657
rect 94522 99144 95274 99657
rect 95442 99144 96102 99657
rect 96270 99144 96930 99657
rect 97098 99144 97850 99657
rect 98018 99144 98678 99657
rect 98846 99144 99506 99657
rect 99674 99144 100426 99657
rect 100594 99144 101254 99657
rect 101422 99144 102082 99657
rect 102250 99144 102910 99657
rect 103078 99144 103830 99657
rect 103998 99144 104658 99657
rect 104826 99144 105486 99657
rect 105654 99144 106406 99657
rect 106574 99144 107234 99657
rect 107402 99144 108062 99657
rect 108230 99144 108982 99657
rect 109150 99144 109810 99657
rect 109978 99144 110638 99657
rect 110806 99144 111466 99657
rect 111634 99144 112386 99657
rect 112554 99144 113214 99657
rect 113382 99144 114042 99657
rect 114210 99144 114962 99657
rect 115130 99144 115790 99657
rect 115958 99144 116618 99657
rect 116786 99144 117538 99657
rect 117706 99144 118366 99657
rect 118534 99144 119194 99657
rect 119362 99144 120022 99657
rect 120190 99144 120942 99657
rect 121110 99144 121770 99657
rect 121938 99144 122598 99657
rect 122766 99144 123518 99657
rect 123686 99144 124346 99657
rect 124514 99144 125174 99657
rect 125342 99144 126094 99657
rect 126262 99144 126922 99657
rect 127090 99144 127750 99657
rect 127918 99144 128578 99657
rect 128746 99144 129498 99657
rect 129666 99144 130326 99657
rect 130494 99144 131154 99657
rect 131322 99144 132074 99657
rect 132242 99144 132902 99657
rect 133070 99144 133730 99657
rect 133898 99144 134650 99657
rect 134818 99144 135478 99657
rect 135646 99144 136306 99657
rect 136474 99144 137134 99657
rect 137302 99144 138054 99657
rect 138222 99144 138882 99657
rect 139050 99144 139710 99657
rect 139878 99144 140630 99657
rect 140798 99144 141458 99657
rect 141626 99144 142286 99657
rect 142454 99144 143206 99657
rect 143374 99144 144034 99657
rect 144202 99144 144862 99657
rect 145030 99144 145690 99657
rect 145858 99144 146610 99657
rect 146778 99144 147438 99657
rect 147606 99144 148266 99657
rect 148434 99144 149186 99657
rect 149354 99144 150014 99657
rect 150182 99144 150842 99657
rect 151010 99144 151762 99657
rect 151930 99144 152590 99657
rect 152758 99144 153418 99657
rect 153586 99144 154246 99657
rect 154414 99144 155166 99657
rect 155334 99144 155994 99657
rect 156162 99144 156822 99657
rect 156990 99144 157742 99657
rect 157910 99144 158570 99657
rect 158738 99144 159398 99657
rect 388 856 159508 99144
rect 388 167 1894 856
rect 2062 167 5758 856
rect 5926 167 9622 856
rect 9790 167 13578 856
rect 13746 167 17442 856
rect 17610 167 21398 856
rect 21566 167 25262 856
rect 25430 167 29126 856
rect 29294 167 33082 856
rect 33250 167 36946 856
rect 37114 167 40902 856
rect 41070 167 44766 856
rect 44934 167 48630 856
rect 48798 167 52586 856
rect 52754 167 56450 856
rect 56618 167 60406 856
rect 60574 167 64270 856
rect 64438 167 68226 856
rect 68394 167 72090 856
rect 72258 167 75954 856
rect 76122 167 79910 856
rect 80078 167 83774 856
rect 83942 167 87730 856
rect 87898 167 91594 856
rect 91762 167 95458 856
rect 95626 167 99414 856
rect 99582 167 103278 856
rect 103446 167 107234 856
rect 107402 167 111098 856
rect 111266 167 115054 856
rect 115222 167 118918 856
rect 119086 167 122782 856
rect 122950 167 126738 856
rect 126906 167 130602 856
rect 130770 167 134558 856
rect 134726 167 138422 856
rect 138590 167 142286 856
rect 142454 167 146242 856
rect 146410 167 150106 856
rect 150274 167 154062 856
rect 154230 167 157926 856
rect 158094 167 159508 856
<< metal3 >>
rect 159200 99560 160000 99680
rect 0 99016 800 99136
rect 159200 99016 160000 99136
rect 159200 98608 160000 98728
rect 159200 98064 160000 98184
rect 159200 97520 160000 97640
rect 0 97248 800 97368
rect 159200 97112 160000 97232
rect 159200 96568 160000 96688
rect 159200 96160 160000 96280
rect 0 95480 800 95600
rect 159200 95616 160000 95736
rect 159200 95072 160000 95192
rect 159200 94664 160000 94784
rect 159200 94120 160000 94240
rect 0 93712 800 93832
rect 159200 93712 160000 93832
rect 159200 93168 160000 93288
rect 159200 92624 160000 92744
rect 159200 92216 160000 92336
rect 0 91944 800 92064
rect 159200 91672 160000 91792
rect 159200 91264 160000 91384
rect 159200 90720 160000 90840
rect 0 90176 800 90296
rect 159200 90176 160000 90296
rect 159200 89768 160000 89888
rect 159200 89224 160000 89344
rect 159200 88816 160000 88936
rect 0 88408 800 88528
rect 159200 88272 160000 88392
rect 159200 87728 160000 87848
rect 159200 87320 160000 87440
rect 0 86640 800 86760
rect 159200 86776 160000 86896
rect 159200 86368 160000 86488
rect 159200 85824 160000 85944
rect 159200 85280 160000 85400
rect 0 84872 800 84992
rect 159200 84872 160000 84992
rect 159200 84328 160000 84448
rect 159200 83920 160000 84040
rect 0 83240 800 83360
rect 159200 83376 160000 83496
rect 159200 82832 160000 82952
rect 159200 82424 160000 82544
rect 159200 81880 160000 82000
rect 0 81472 800 81592
rect 159200 81472 160000 81592
rect 159200 80928 160000 81048
rect 159200 80384 160000 80504
rect 159200 79976 160000 80096
rect 0 79704 800 79824
rect 159200 79432 160000 79552
rect 159200 79024 160000 79144
rect 159200 78480 160000 78600
rect 0 77936 800 78056
rect 159200 77936 160000 78056
rect 159200 77528 160000 77648
rect 159200 76984 160000 77104
rect 159200 76576 160000 76696
rect 0 76168 800 76288
rect 159200 76032 160000 76152
rect 159200 75488 160000 75608
rect 159200 75080 160000 75200
rect 0 74400 800 74520
rect 159200 74536 160000 74656
rect 159200 74128 160000 74248
rect 159200 73584 160000 73704
rect 159200 73040 160000 73160
rect 0 72632 800 72752
rect 159200 72632 160000 72752
rect 159200 72088 160000 72208
rect 159200 71680 160000 71800
rect 159200 71136 160000 71256
rect 0 70864 800 70984
rect 159200 70592 160000 70712
rect 159200 70184 160000 70304
rect 159200 69640 160000 69760
rect 0 69096 800 69216
rect 159200 69232 160000 69352
rect 159200 68688 160000 68808
rect 159200 68144 160000 68264
rect 159200 67736 160000 67856
rect 0 67464 800 67584
rect 159200 67192 160000 67312
rect 159200 66784 160000 66904
rect 159200 66240 160000 66360
rect 0 65696 800 65816
rect 159200 65696 160000 65816
rect 159200 65288 160000 65408
rect 159200 64744 160000 64864
rect 159200 64200 160000 64320
rect 0 63928 800 64048
rect 159200 63792 160000 63912
rect 159200 63248 160000 63368
rect 159200 62840 160000 62960
rect 0 62160 800 62280
rect 159200 62296 160000 62416
rect 159200 61752 160000 61872
rect 159200 61344 160000 61464
rect 159200 60800 160000 60920
rect 0 60392 800 60512
rect 159200 60392 160000 60512
rect 159200 59848 160000 59968
rect 159200 59304 160000 59424
rect 159200 58896 160000 59016
rect 0 58624 800 58744
rect 159200 58352 160000 58472
rect 159200 57944 160000 58064
rect 159200 57400 160000 57520
rect 0 56856 800 56976
rect 159200 56856 160000 56976
rect 159200 56448 160000 56568
rect 159200 55904 160000 56024
rect 159200 55496 160000 55616
rect 0 55088 800 55208
rect 159200 54952 160000 55072
rect 159200 54408 160000 54528
rect 159200 54000 160000 54120
rect 0 53320 800 53440
rect 159200 53456 160000 53576
rect 159200 53048 160000 53168
rect 159200 52504 160000 52624
rect 159200 51960 160000 52080
rect 0 51552 800 51672
rect 159200 51552 160000 51672
rect 159200 51008 160000 51128
rect 159200 50600 160000 50720
rect 0 49920 800 50040
rect 159200 50056 160000 50176
rect 159200 49512 160000 49632
rect 159200 49104 160000 49224
rect 159200 48560 160000 48680
rect 0 48152 800 48272
rect 159200 48152 160000 48272
rect 159200 47608 160000 47728
rect 159200 47064 160000 47184
rect 159200 46656 160000 46776
rect 0 46384 800 46504
rect 159200 46112 160000 46232
rect 159200 45704 160000 45824
rect 159200 45160 160000 45280
rect 0 44616 800 44736
rect 159200 44616 160000 44736
rect 159200 44208 160000 44328
rect 159200 43664 160000 43784
rect 159200 43256 160000 43376
rect 0 42848 800 42968
rect 159200 42712 160000 42832
rect 159200 42168 160000 42288
rect 159200 41760 160000 41880
rect 0 41080 800 41200
rect 159200 41216 160000 41336
rect 159200 40808 160000 40928
rect 159200 40264 160000 40384
rect 159200 39720 160000 39840
rect 0 39312 800 39432
rect 159200 39312 160000 39432
rect 159200 38768 160000 38888
rect 159200 38360 160000 38480
rect 159200 37816 160000 37936
rect 0 37544 800 37664
rect 159200 37272 160000 37392
rect 159200 36864 160000 36984
rect 159200 36320 160000 36440
rect 0 35776 800 35896
rect 159200 35912 160000 36032
rect 159200 35368 160000 35488
rect 159200 34824 160000 34944
rect 159200 34416 160000 34536
rect 0 34144 800 34264
rect 159200 33872 160000 33992
rect 159200 33464 160000 33584
rect 159200 32920 160000 33040
rect 0 32376 800 32496
rect 159200 32376 160000 32496
rect 159200 31968 160000 32088
rect 159200 31424 160000 31544
rect 159200 30880 160000 31000
rect 0 30608 800 30728
rect 159200 30472 160000 30592
rect 159200 29928 160000 30048
rect 159200 29520 160000 29640
rect 0 28840 800 28960
rect 159200 28976 160000 29096
rect 159200 28432 160000 28552
rect 159200 28024 160000 28144
rect 159200 27480 160000 27600
rect 0 27072 800 27192
rect 159200 27072 160000 27192
rect 159200 26528 160000 26648
rect 159200 25984 160000 26104
rect 159200 25576 160000 25696
rect 0 25304 800 25424
rect 159200 25032 160000 25152
rect 159200 24624 160000 24744
rect 159200 24080 160000 24200
rect 0 23536 800 23656
rect 159200 23536 160000 23656
rect 159200 23128 160000 23248
rect 159200 22584 160000 22704
rect 159200 22176 160000 22296
rect 0 21768 800 21888
rect 159200 21632 160000 21752
rect 159200 21088 160000 21208
rect 159200 20680 160000 20800
rect 0 20000 800 20120
rect 159200 20136 160000 20256
rect 159200 19728 160000 19848
rect 159200 19184 160000 19304
rect 159200 18640 160000 18760
rect 0 18232 800 18352
rect 159200 18232 160000 18352
rect 159200 17688 160000 17808
rect 159200 17280 160000 17400
rect 0 16600 800 16720
rect 159200 16736 160000 16856
rect 159200 16192 160000 16312
rect 159200 15784 160000 15904
rect 159200 15240 160000 15360
rect 0 14832 800 14952
rect 159200 14832 160000 14952
rect 159200 14288 160000 14408
rect 159200 13744 160000 13864
rect 159200 13336 160000 13456
rect 0 13064 800 13184
rect 159200 12792 160000 12912
rect 159200 12384 160000 12504
rect 159200 11840 160000 11960
rect 0 11296 800 11416
rect 159200 11296 160000 11416
rect 159200 10888 160000 11008
rect 159200 10344 160000 10464
rect 159200 9936 160000 10056
rect 0 9528 800 9648
rect 159200 9392 160000 9512
rect 159200 8848 160000 8968
rect 159200 8440 160000 8560
rect 0 7760 800 7880
rect 159200 7896 160000 8016
rect 159200 7488 160000 7608
rect 159200 6944 160000 7064
rect 159200 6400 160000 6520
rect 0 5992 800 6112
rect 159200 5992 160000 6112
rect 159200 5448 160000 5568
rect 159200 5040 160000 5160
rect 159200 4496 160000 4616
rect 0 4224 800 4344
rect 159200 3952 160000 4072
rect 159200 3544 160000 3664
rect 159200 3000 160000 3120
rect 0 2456 800 2576
rect 159200 2592 160000 2712
rect 159200 2048 160000 2168
rect 159200 1504 160000 1624
rect 159200 1096 160000 1216
rect 0 824 800 944
rect 159200 552 160000 672
rect 159200 144 160000 264
<< obsm3 >>
rect 800 99480 159120 99653
rect 800 99216 159200 99480
rect 880 98936 159120 99216
rect 800 98808 159200 98936
rect 800 98528 159120 98808
rect 800 98264 159200 98528
rect 800 97984 159120 98264
rect 800 97720 159200 97984
rect 800 97448 159120 97720
rect 880 97440 159120 97448
rect 880 97312 159200 97440
rect 880 97168 159120 97312
rect 800 97032 159120 97168
rect 800 96768 159200 97032
rect 800 96488 159120 96768
rect 800 96360 159200 96488
rect 800 96080 159120 96360
rect 800 95816 159200 96080
rect 800 95680 159120 95816
rect 880 95536 159120 95680
rect 880 95400 159200 95536
rect 800 95272 159200 95400
rect 800 94992 159120 95272
rect 800 94864 159200 94992
rect 800 94584 159120 94864
rect 800 94320 159200 94584
rect 800 94040 159120 94320
rect 800 93912 159200 94040
rect 880 93632 159120 93912
rect 800 93368 159200 93632
rect 800 93088 159120 93368
rect 800 92824 159200 93088
rect 800 92544 159120 92824
rect 800 92416 159200 92544
rect 800 92144 159120 92416
rect 880 92136 159120 92144
rect 880 91872 159200 92136
rect 880 91864 159120 91872
rect 800 91592 159120 91864
rect 800 91464 159200 91592
rect 800 91184 159120 91464
rect 800 90920 159200 91184
rect 800 90640 159120 90920
rect 800 90376 159200 90640
rect 880 90096 159120 90376
rect 800 89968 159200 90096
rect 800 89688 159120 89968
rect 800 89424 159200 89688
rect 800 89144 159120 89424
rect 800 89016 159200 89144
rect 800 88736 159120 89016
rect 800 88608 159200 88736
rect 880 88472 159200 88608
rect 880 88328 159120 88472
rect 800 88192 159120 88328
rect 800 87928 159200 88192
rect 800 87648 159120 87928
rect 800 87520 159200 87648
rect 800 87240 159120 87520
rect 800 86976 159200 87240
rect 800 86840 159120 86976
rect 880 86696 159120 86840
rect 880 86568 159200 86696
rect 880 86560 159120 86568
rect 800 86288 159120 86560
rect 800 86024 159200 86288
rect 800 85744 159120 86024
rect 800 85480 159200 85744
rect 800 85200 159120 85480
rect 800 85072 159200 85200
rect 880 84792 159120 85072
rect 800 84528 159200 84792
rect 800 84248 159120 84528
rect 800 84120 159200 84248
rect 800 83840 159120 84120
rect 800 83576 159200 83840
rect 800 83440 159120 83576
rect 880 83296 159120 83440
rect 880 83160 159200 83296
rect 800 83032 159200 83160
rect 800 82752 159120 83032
rect 800 82624 159200 82752
rect 800 82344 159120 82624
rect 800 82080 159200 82344
rect 800 81800 159120 82080
rect 800 81672 159200 81800
rect 880 81392 159120 81672
rect 800 81128 159200 81392
rect 800 80848 159120 81128
rect 800 80584 159200 80848
rect 800 80304 159120 80584
rect 800 80176 159200 80304
rect 800 79904 159120 80176
rect 880 79896 159120 79904
rect 880 79632 159200 79896
rect 880 79624 159120 79632
rect 800 79352 159120 79624
rect 800 79224 159200 79352
rect 800 78944 159120 79224
rect 800 78680 159200 78944
rect 800 78400 159120 78680
rect 800 78136 159200 78400
rect 880 77856 159120 78136
rect 800 77728 159200 77856
rect 800 77448 159120 77728
rect 800 77184 159200 77448
rect 800 76904 159120 77184
rect 800 76776 159200 76904
rect 800 76496 159120 76776
rect 800 76368 159200 76496
rect 880 76232 159200 76368
rect 880 76088 159120 76232
rect 800 75952 159120 76088
rect 800 75688 159200 75952
rect 800 75408 159120 75688
rect 800 75280 159200 75408
rect 800 75000 159120 75280
rect 800 74736 159200 75000
rect 800 74600 159120 74736
rect 880 74456 159120 74600
rect 880 74328 159200 74456
rect 880 74320 159120 74328
rect 800 74048 159120 74320
rect 800 73784 159200 74048
rect 800 73504 159120 73784
rect 800 73240 159200 73504
rect 800 72960 159120 73240
rect 800 72832 159200 72960
rect 880 72552 159120 72832
rect 800 72288 159200 72552
rect 800 72008 159120 72288
rect 800 71880 159200 72008
rect 800 71600 159120 71880
rect 800 71336 159200 71600
rect 800 71064 159120 71336
rect 880 71056 159120 71064
rect 880 70792 159200 71056
rect 880 70784 159120 70792
rect 800 70512 159120 70784
rect 800 70384 159200 70512
rect 800 70104 159120 70384
rect 800 69840 159200 70104
rect 800 69560 159120 69840
rect 800 69432 159200 69560
rect 800 69296 159120 69432
rect 880 69152 159120 69296
rect 880 69016 159200 69152
rect 800 68888 159200 69016
rect 800 68608 159120 68888
rect 800 68344 159200 68608
rect 800 68064 159120 68344
rect 800 67936 159200 68064
rect 800 67664 159120 67936
rect 880 67656 159120 67664
rect 880 67392 159200 67656
rect 880 67384 159120 67392
rect 800 67112 159120 67384
rect 800 66984 159200 67112
rect 800 66704 159120 66984
rect 800 66440 159200 66704
rect 800 66160 159120 66440
rect 800 65896 159200 66160
rect 880 65616 159120 65896
rect 800 65488 159200 65616
rect 800 65208 159120 65488
rect 800 64944 159200 65208
rect 800 64664 159120 64944
rect 800 64400 159200 64664
rect 800 64128 159120 64400
rect 880 64120 159120 64128
rect 880 63992 159200 64120
rect 880 63848 159120 63992
rect 800 63712 159120 63848
rect 800 63448 159200 63712
rect 800 63168 159120 63448
rect 800 63040 159200 63168
rect 800 62760 159120 63040
rect 800 62496 159200 62760
rect 800 62360 159120 62496
rect 880 62216 159120 62360
rect 880 62080 159200 62216
rect 800 61952 159200 62080
rect 800 61672 159120 61952
rect 800 61544 159200 61672
rect 800 61264 159120 61544
rect 800 61000 159200 61264
rect 800 60720 159120 61000
rect 800 60592 159200 60720
rect 880 60312 159120 60592
rect 800 60048 159200 60312
rect 800 59768 159120 60048
rect 800 59504 159200 59768
rect 800 59224 159120 59504
rect 800 59096 159200 59224
rect 800 58824 159120 59096
rect 880 58816 159120 58824
rect 880 58552 159200 58816
rect 880 58544 159120 58552
rect 800 58272 159120 58544
rect 800 58144 159200 58272
rect 800 57864 159120 58144
rect 800 57600 159200 57864
rect 800 57320 159120 57600
rect 800 57056 159200 57320
rect 880 56776 159120 57056
rect 800 56648 159200 56776
rect 800 56368 159120 56648
rect 800 56104 159200 56368
rect 800 55824 159120 56104
rect 800 55696 159200 55824
rect 800 55416 159120 55696
rect 800 55288 159200 55416
rect 880 55152 159200 55288
rect 880 55008 159120 55152
rect 800 54872 159120 55008
rect 800 54608 159200 54872
rect 800 54328 159120 54608
rect 800 54200 159200 54328
rect 800 53920 159120 54200
rect 800 53656 159200 53920
rect 800 53520 159120 53656
rect 880 53376 159120 53520
rect 880 53248 159200 53376
rect 880 53240 159120 53248
rect 800 52968 159120 53240
rect 800 52704 159200 52968
rect 800 52424 159120 52704
rect 800 52160 159200 52424
rect 800 51880 159120 52160
rect 800 51752 159200 51880
rect 880 51472 159120 51752
rect 800 51208 159200 51472
rect 800 50928 159120 51208
rect 800 50800 159200 50928
rect 800 50520 159120 50800
rect 800 50256 159200 50520
rect 800 50120 159120 50256
rect 880 49976 159120 50120
rect 880 49840 159200 49976
rect 800 49712 159200 49840
rect 800 49432 159120 49712
rect 800 49304 159200 49432
rect 800 49024 159120 49304
rect 800 48760 159200 49024
rect 800 48480 159120 48760
rect 800 48352 159200 48480
rect 880 48072 159120 48352
rect 800 47808 159200 48072
rect 800 47528 159120 47808
rect 800 47264 159200 47528
rect 800 46984 159120 47264
rect 800 46856 159200 46984
rect 800 46584 159120 46856
rect 880 46576 159120 46584
rect 880 46312 159200 46576
rect 880 46304 159120 46312
rect 800 46032 159120 46304
rect 800 45904 159200 46032
rect 800 45624 159120 45904
rect 800 45360 159200 45624
rect 800 45080 159120 45360
rect 800 44816 159200 45080
rect 880 44536 159120 44816
rect 800 44408 159200 44536
rect 800 44128 159120 44408
rect 800 43864 159200 44128
rect 800 43584 159120 43864
rect 800 43456 159200 43584
rect 800 43176 159120 43456
rect 800 43048 159200 43176
rect 880 42912 159200 43048
rect 880 42768 159120 42912
rect 800 42632 159120 42768
rect 800 42368 159200 42632
rect 800 42088 159120 42368
rect 800 41960 159200 42088
rect 800 41680 159120 41960
rect 800 41416 159200 41680
rect 800 41280 159120 41416
rect 880 41136 159120 41280
rect 880 41008 159200 41136
rect 880 41000 159120 41008
rect 800 40728 159120 41000
rect 800 40464 159200 40728
rect 800 40184 159120 40464
rect 800 39920 159200 40184
rect 800 39640 159120 39920
rect 800 39512 159200 39640
rect 880 39232 159120 39512
rect 800 38968 159200 39232
rect 800 38688 159120 38968
rect 800 38560 159200 38688
rect 800 38280 159120 38560
rect 800 38016 159200 38280
rect 800 37744 159120 38016
rect 880 37736 159120 37744
rect 880 37472 159200 37736
rect 880 37464 159120 37472
rect 800 37192 159120 37464
rect 800 37064 159200 37192
rect 800 36784 159120 37064
rect 800 36520 159200 36784
rect 800 36240 159120 36520
rect 800 36112 159200 36240
rect 800 35976 159120 36112
rect 880 35832 159120 35976
rect 880 35696 159200 35832
rect 800 35568 159200 35696
rect 800 35288 159120 35568
rect 800 35024 159200 35288
rect 800 34744 159120 35024
rect 800 34616 159200 34744
rect 800 34344 159120 34616
rect 880 34336 159120 34344
rect 880 34072 159200 34336
rect 880 34064 159120 34072
rect 800 33792 159120 34064
rect 800 33664 159200 33792
rect 800 33384 159120 33664
rect 800 33120 159200 33384
rect 800 32840 159120 33120
rect 800 32576 159200 32840
rect 880 32296 159120 32576
rect 800 32168 159200 32296
rect 800 31888 159120 32168
rect 800 31624 159200 31888
rect 800 31344 159120 31624
rect 800 31080 159200 31344
rect 800 30808 159120 31080
rect 880 30800 159120 30808
rect 880 30672 159200 30800
rect 880 30528 159120 30672
rect 800 30392 159120 30528
rect 800 30128 159200 30392
rect 800 29848 159120 30128
rect 800 29720 159200 29848
rect 800 29440 159120 29720
rect 800 29176 159200 29440
rect 800 29040 159120 29176
rect 880 28896 159120 29040
rect 880 28760 159200 28896
rect 800 28632 159200 28760
rect 800 28352 159120 28632
rect 800 28224 159200 28352
rect 800 27944 159120 28224
rect 800 27680 159200 27944
rect 800 27400 159120 27680
rect 800 27272 159200 27400
rect 880 26992 159120 27272
rect 800 26728 159200 26992
rect 800 26448 159120 26728
rect 800 26184 159200 26448
rect 800 25904 159120 26184
rect 800 25776 159200 25904
rect 800 25504 159120 25776
rect 880 25496 159120 25504
rect 880 25232 159200 25496
rect 880 25224 159120 25232
rect 800 24952 159120 25224
rect 800 24824 159200 24952
rect 800 24544 159120 24824
rect 800 24280 159200 24544
rect 800 24000 159120 24280
rect 800 23736 159200 24000
rect 880 23456 159120 23736
rect 800 23328 159200 23456
rect 800 23048 159120 23328
rect 800 22784 159200 23048
rect 800 22504 159120 22784
rect 800 22376 159200 22504
rect 800 22096 159120 22376
rect 800 21968 159200 22096
rect 880 21832 159200 21968
rect 880 21688 159120 21832
rect 800 21552 159120 21688
rect 800 21288 159200 21552
rect 800 21008 159120 21288
rect 800 20880 159200 21008
rect 800 20600 159120 20880
rect 800 20336 159200 20600
rect 800 20200 159120 20336
rect 880 20056 159120 20200
rect 880 19928 159200 20056
rect 880 19920 159120 19928
rect 800 19648 159120 19920
rect 800 19384 159200 19648
rect 800 19104 159120 19384
rect 800 18840 159200 19104
rect 800 18560 159120 18840
rect 800 18432 159200 18560
rect 880 18152 159120 18432
rect 800 17888 159200 18152
rect 800 17608 159120 17888
rect 800 17480 159200 17608
rect 800 17200 159120 17480
rect 800 16936 159200 17200
rect 800 16800 159120 16936
rect 880 16656 159120 16800
rect 880 16520 159200 16656
rect 800 16392 159200 16520
rect 800 16112 159120 16392
rect 800 15984 159200 16112
rect 800 15704 159120 15984
rect 800 15440 159200 15704
rect 800 15160 159120 15440
rect 800 15032 159200 15160
rect 880 14752 159120 15032
rect 800 14488 159200 14752
rect 800 14208 159120 14488
rect 800 13944 159200 14208
rect 800 13664 159120 13944
rect 800 13536 159200 13664
rect 800 13264 159120 13536
rect 880 13256 159120 13264
rect 880 12992 159200 13256
rect 880 12984 159120 12992
rect 800 12712 159120 12984
rect 800 12584 159200 12712
rect 800 12304 159120 12584
rect 800 12040 159200 12304
rect 800 11760 159120 12040
rect 800 11496 159200 11760
rect 880 11216 159120 11496
rect 800 11088 159200 11216
rect 800 10808 159120 11088
rect 800 10544 159200 10808
rect 800 10264 159120 10544
rect 800 10136 159200 10264
rect 800 9856 159120 10136
rect 800 9728 159200 9856
rect 880 9592 159200 9728
rect 880 9448 159120 9592
rect 800 9312 159120 9448
rect 800 9048 159200 9312
rect 800 8768 159120 9048
rect 800 8640 159200 8768
rect 800 8360 159120 8640
rect 800 8096 159200 8360
rect 800 7960 159120 8096
rect 880 7816 159120 7960
rect 880 7688 159200 7816
rect 880 7680 159120 7688
rect 800 7408 159120 7680
rect 800 7144 159200 7408
rect 800 6864 159120 7144
rect 800 6600 159200 6864
rect 800 6320 159120 6600
rect 800 6192 159200 6320
rect 880 5912 159120 6192
rect 800 5648 159200 5912
rect 800 5368 159120 5648
rect 800 5240 159200 5368
rect 800 4960 159120 5240
rect 800 4696 159200 4960
rect 800 4424 159120 4696
rect 880 4416 159120 4424
rect 880 4152 159200 4416
rect 880 4144 159120 4152
rect 800 3872 159120 4144
rect 800 3744 159200 3872
rect 800 3464 159120 3744
rect 800 3200 159200 3464
rect 800 2920 159120 3200
rect 800 2792 159200 2920
rect 800 2656 159120 2792
rect 880 2512 159120 2656
rect 880 2376 159200 2512
rect 800 2248 159200 2376
rect 800 1968 159120 2248
rect 800 1704 159200 1968
rect 800 1424 159120 1704
rect 800 1296 159200 1424
rect 800 1024 159120 1296
rect 880 1016 159120 1024
rect 880 752 159200 1016
rect 880 744 159120 752
rect 800 472 159120 744
rect 800 344 159200 472
rect 800 171 159120 344
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
rect 111728 2128 112048 97424
rect 127088 2128 127408 97424
rect 142448 2128 142768 97424
rect 157808 2128 158128 97424
<< obsm4 >>
rect 156275 57019 157077 94349
<< labels >>
rlabel metal2 s 5446 99200 5502 100000 6 addr0[0]
port 1 nsew signal output
rlabel metal2 s 6366 99200 6422 100000 6 addr0[1]
port 2 nsew signal output
rlabel metal2 s 7194 99200 7250 100000 6 addr0[2]
port 3 nsew signal output
rlabel metal2 s 8022 99200 8078 100000 6 addr0[3]
port 4 nsew signal output
rlabel metal2 s 8850 99200 8906 100000 6 addr0[4]
port 5 nsew signal output
rlabel metal2 s 9770 99200 9826 100000 6 addr0[5]
port 6 nsew signal output
rlabel metal2 s 10598 99200 10654 100000 6 addr0[6]
port 7 nsew signal output
rlabel metal2 s 11426 99200 11482 100000 6 addr0[7]
port 8 nsew signal output
rlabel metal2 s 12346 99200 12402 100000 6 addr0[8]
port 9 nsew signal output
rlabel metal2 s 96158 99200 96214 100000 6 addr1[0]
port 10 nsew signal output
rlabel metal2 s 96986 99200 97042 100000 6 addr1[1]
port 11 nsew signal output
rlabel metal2 s 97906 99200 97962 100000 6 addr1[2]
port 12 nsew signal output
rlabel metal2 s 98734 99200 98790 100000 6 addr1[3]
port 13 nsew signal output
rlabel metal2 s 99562 99200 99618 100000 6 addr1[4]
port 14 nsew signal output
rlabel metal2 s 100482 99200 100538 100000 6 addr1[5]
port 15 nsew signal output
rlabel metal2 s 101310 99200 101366 100000 6 addr1[6]
port 16 nsew signal output
rlabel metal2 s 102138 99200 102194 100000 6 addr1[7]
port 17 nsew signal output
rlabel metal2 s 102966 99200 103022 100000 6 addr1[8]
port 18 nsew signal output
rlabel metal2 s 386 99200 442 100000 6 clk0
port 19 nsew signal output
rlabel metal2 s 95330 99200 95386 100000 6 clk1
port 20 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 159200 1096 160000 1216 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 159200 3952 160000 4072 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 159200 20680 160000 20800 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 159200 22176 160000 22296 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 159200 23536 160000 23656 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 159200 25032 160000 25152 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 159200 26528 160000 26648 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 159200 28024 160000 28144 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 159200 29520 160000 29640 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 159200 30880 160000 31000 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 159200 32376 160000 32496 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 159200 33872 160000 33992 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 159200 5992 160000 6112 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 159200 35368 160000 35488 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 159200 36864 160000 36984 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 159200 38360 160000 38480 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 159200 39720 160000 39840 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 159200 41216 160000 41336 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 159200 42712 160000 42832 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 159200 44208 160000 44328 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 159200 45704 160000 45824 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 159200 7896 160000 8016 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 159200 9936 160000 10056 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 159200 11840 160000 11960 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 159200 13336 160000 13456 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 159200 14832 160000 14952 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 159200 16192 160000 16312 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 159200 17688 160000 17808 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 159200 19184 160000 19304 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 159200 1504 160000 1624 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 159200 4496 160000 4616 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 159200 21088 160000 21208 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 159200 22584 160000 22704 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 159200 24080 160000 24200 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 159200 25576 160000 25696 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 159200 27072 160000 27192 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 159200 28432 160000 28552 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 159200 29928 160000 30048 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 159200 31424 160000 31544 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 159200 32920 160000 33040 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 159200 34416 160000 34536 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 159200 6400 160000 6520 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 159200 35912 160000 36032 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 159200 37272 160000 37392 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 159200 38768 160000 38888 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 159200 40264 160000 40384 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 159200 41760 160000 41880 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 159200 43256 160000 43376 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 159200 44616 160000 44736 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 159200 46112 160000 46232 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 159200 47064 160000 47184 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 159200 48152 160000 48272 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 159200 8440 160000 8560 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 159200 49104 160000 49224 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 159200 50056 160000 50176 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 159200 10344 160000 10464 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 159200 12384 160000 12504 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 159200 13744 160000 13864 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 159200 15240 160000 15360 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 159200 16736 160000 16856 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 159200 18232 160000 18352 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 159200 19728 160000 19848 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 159200 5040 160000 5160 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 159200 21632 160000 21752 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 159200 23128 160000 23248 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 159200 24624 160000 24744 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 159200 25984 160000 26104 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 159200 27480 160000 27600 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 159200 28976 160000 29096 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 159200 30472 160000 30592 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 159200 31968 160000 32088 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 159200 33464 160000 33584 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 159200 34824 160000 34944 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 159200 6944 160000 7064 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 159200 36320 160000 36440 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 159200 37816 160000 37936 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 159200 39312 160000 39432 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 159200 40808 160000 40928 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 159200 42168 160000 42288 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 159200 43664 160000 43784 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 159200 45160 160000 45280 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 159200 46656 160000 46776 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 159200 47608 160000 47728 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 159200 48560 160000 48680 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 159200 8848 160000 8968 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 159200 49512 160000 49632 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 159200 50600 160000 50720 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 159200 10888 160000 11008 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 159200 12792 160000 12912 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 159200 14288 160000 14408 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 159200 15784 160000 15904 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 159200 17280 160000 17400 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 159200 18640 160000 18760 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 159200 20136 160000 20256 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 159200 2048 160000 2168 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 159200 5448 160000 5568 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 159200 7488 160000 7608 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 159200 9392 160000 9512 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 159200 11296 160000 11416 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 159200 2592 160000 2712 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 159200 3000 160000 3120 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 159200 3544 160000 3664 6 core_wb_we_o
port 130 nsew signal output
rlabel metal2 s 158626 99200 158682 100000 6 csb0[0]
port 131 nsew signal output
rlabel metal2 s 159454 99200 159510 100000 6 csb0[1]
port 132 nsew signal output
rlabel metal2 s 157982 0 158038 800 6 csb1[0]
port 133 nsew signal output
rlabel metal3 s 159200 99560 160000 99680 6 csb1[1]
port 134 nsew signal output
rlabel metal2 s 13174 99200 13230 100000 6 din0[0]
port 135 nsew signal output
rlabel metal2 s 21730 99200 21786 100000 6 din0[10]
port 136 nsew signal output
rlabel metal2 s 22558 99200 22614 100000 6 din0[11]
port 137 nsew signal output
rlabel metal2 s 23478 99200 23534 100000 6 din0[12]
port 138 nsew signal output
rlabel metal2 s 24306 99200 24362 100000 6 din0[13]
port 139 nsew signal output
rlabel metal2 s 25134 99200 25190 100000 6 din0[14]
port 140 nsew signal output
rlabel metal2 s 25962 99200 26018 100000 6 din0[15]
port 141 nsew signal output
rlabel metal2 s 26882 99200 26938 100000 6 din0[16]
port 142 nsew signal output
rlabel metal2 s 27710 99200 27766 100000 6 din0[17]
port 143 nsew signal output
rlabel metal2 s 28538 99200 28594 100000 6 din0[18]
port 144 nsew signal output
rlabel metal2 s 29458 99200 29514 100000 6 din0[19]
port 145 nsew signal output
rlabel metal2 s 14002 99200 14058 100000 6 din0[1]
port 146 nsew signal output
rlabel metal2 s 30286 99200 30342 100000 6 din0[20]
port 147 nsew signal output
rlabel metal2 s 31114 99200 31170 100000 6 din0[21]
port 148 nsew signal output
rlabel metal2 s 32034 99200 32090 100000 6 din0[22]
port 149 nsew signal output
rlabel metal2 s 32862 99200 32918 100000 6 din0[23]
port 150 nsew signal output
rlabel metal2 s 33690 99200 33746 100000 6 din0[24]
port 151 nsew signal output
rlabel metal2 s 34518 99200 34574 100000 6 din0[25]
port 152 nsew signal output
rlabel metal2 s 35438 99200 35494 100000 6 din0[26]
port 153 nsew signal output
rlabel metal2 s 36266 99200 36322 100000 6 din0[27]
port 154 nsew signal output
rlabel metal2 s 37094 99200 37150 100000 6 din0[28]
port 155 nsew signal output
rlabel metal2 s 38014 99200 38070 100000 6 din0[29]
port 156 nsew signal output
rlabel metal2 s 14922 99200 14978 100000 6 din0[2]
port 157 nsew signal output
rlabel metal2 s 38842 99200 38898 100000 6 din0[30]
port 158 nsew signal output
rlabel metal2 s 39670 99200 39726 100000 6 din0[31]
port 159 nsew signal output
rlabel metal2 s 15750 99200 15806 100000 6 din0[3]
port 160 nsew signal output
rlabel metal2 s 16578 99200 16634 100000 6 din0[4]
port 161 nsew signal output
rlabel metal2 s 17406 99200 17462 100000 6 din0[5]
port 162 nsew signal output
rlabel metal2 s 18326 99200 18382 100000 6 din0[6]
port 163 nsew signal output
rlabel metal2 s 19154 99200 19210 100000 6 din0[7]
port 164 nsew signal output
rlabel metal2 s 19982 99200 20038 100000 6 din0[8]
port 165 nsew signal output
rlabel metal2 s 20902 99200 20958 100000 6 din0[9]
port 166 nsew signal output
rlabel metal2 s 40590 99200 40646 100000 6 dout0[0]
port 167 nsew signal input
rlabel metal2 s 49146 99200 49202 100000 6 dout0[10]
port 168 nsew signal input
rlabel metal2 s 49974 99200 50030 100000 6 dout0[11]
port 169 nsew signal input
rlabel metal2 s 50802 99200 50858 100000 6 dout0[12]
port 170 nsew signal input
rlabel metal2 s 51630 99200 51686 100000 6 dout0[13]
port 171 nsew signal input
rlabel metal2 s 52550 99200 52606 100000 6 dout0[14]
port 172 nsew signal input
rlabel metal2 s 53378 99200 53434 100000 6 dout0[15]
port 173 nsew signal input
rlabel metal2 s 54206 99200 54262 100000 6 dout0[16]
port 174 nsew signal input
rlabel metal2 s 55126 99200 55182 100000 6 dout0[17]
port 175 nsew signal input
rlabel metal2 s 55954 99200 56010 100000 6 dout0[18]
port 176 nsew signal input
rlabel metal2 s 56782 99200 56838 100000 6 dout0[19]
port 177 nsew signal input
rlabel metal2 s 41418 99200 41474 100000 6 dout0[1]
port 178 nsew signal input
rlabel metal2 s 57702 99200 57758 100000 6 dout0[20]
port 179 nsew signal input
rlabel metal2 s 58530 99200 58586 100000 6 dout0[21]
port 180 nsew signal input
rlabel metal2 s 59358 99200 59414 100000 6 dout0[22]
port 181 nsew signal input
rlabel metal2 s 60186 99200 60242 100000 6 dout0[23]
port 182 nsew signal input
rlabel metal2 s 61106 99200 61162 100000 6 dout0[24]
port 183 nsew signal input
rlabel metal2 s 61934 99200 61990 100000 6 dout0[25]
port 184 nsew signal input
rlabel metal2 s 62762 99200 62818 100000 6 dout0[26]
port 185 nsew signal input
rlabel metal2 s 63682 99200 63738 100000 6 dout0[27]
port 186 nsew signal input
rlabel metal2 s 64510 99200 64566 100000 6 dout0[28]
port 187 nsew signal input
rlabel metal2 s 65338 99200 65394 100000 6 dout0[29]
port 188 nsew signal input
rlabel metal2 s 42246 99200 42302 100000 6 dout0[2]
port 189 nsew signal input
rlabel metal2 s 66258 99200 66314 100000 6 dout0[30]
port 190 nsew signal input
rlabel metal2 s 67086 99200 67142 100000 6 dout0[31]
port 191 nsew signal input
rlabel metal2 s 67914 99200 67970 100000 6 dout0[32]
port 192 nsew signal input
rlabel metal2 s 68742 99200 68798 100000 6 dout0[33]
port 193 nsew signal input
rlabel metal2 s 69662 99200 69718 100000 6 dout0[34]
port 194 nsew signal input
rlabel metal2 s 70490 99200 70546 100000 6 dout0[35]
port 195 nsew signal input
rlabel metal2 s 71318 99200 71374 100000 6 dout0[36]
port 196 nsew signal input
rlabel metal2 s 72238 99200 72294 100000 6 dout0[37]
port 197 nsew signal input
rlabel metal2 s 73066 99200 73122 100000 6 dout0[38]
port 198 nsew signal input
rlabel metal2 s 73894 99200 73950 100000 6 dout0[39]
port 199 nsew signal input
rlabel metal2 s 43074 99200 43130 100000 6 dout0[3]
port 200 nsew signal input
rlabel metal2 s 74814 99200 74870 100000 6 dout0[40]
port 201 nsew signal input
rlabel metal2 s 75642 99200 75698 100000 6 dout0[41]
port 202 nsew signal input
rlabel metal2 s 76470 99200 76526 100000 6 dout0[42]
port 203 nsew signal input
rlabel metal2 s 77298 99200 77354 100000 6 dout0[43]
port 204 nsew signal input
rlabel metal2 s 78218 99200 78274 100000 6 dout0[44]
port 205 nsew signal input
rlabel metal2 s 79046 99200 79102 100000 6 dout0[45]
port 206 nsew signal input
rlabel metal2 s 79874 99200 79930 100000 6 dout0[46]
port 207 nsew signal input
rlabel metal2 s 80794 99200 80850 100000 6 dout0[47]
port 208 nsew signal input
rlabel metal2 s 81622 99200 81678 100000 6 dout0[48]
port 209 nsew signal input
rlabel metal2 s 82450 99200 82506 100000 6 dout0[49]
port 210 nsew signal input
rlabel metal2 s 43994 99200 44050 100000 6 dout0[4]
port 211 nsew signal input
rlabel metal2 s 83370 99200 83426 100000 6 dout0[50]
port 212 nsew signal input
rlabel metal2 s 84198 99200 84254 100000 6 dout0[51]
port 213 nsew signal input
rlabel metal2 s 85026 99200 85082 100000 6 dout0[52]
port 214 nsew signal input
rlabel metal2 s 85854 99200 85910 100000 6 dout0[53]
port 215 nsew signal input
rlabel metal2 s 86774 99200 86830 100000 6 dout0[54]
port 216 nsew signal input
rlabel metal2 s 87602 99200 87658 100000 6 dout0[55]
port 217 nsew signal input
rlabel metal2 s 88430 99200 88486 100000 6 dout0[56]
port 218 nsew signal input
rlabel metal2 s 89350 99200 89406 100000 6 dout0[57]
port 219 nsew signal input
rlabel metal2 s 90178 99200 90234 100000 6 dout0[58]
port 220 nsew signal input
rlabel metal2 s 91006 99200 91062 100000 6 dout0[59]
port 221 nsew signal input
rlabel metal2 s 44822 99200 44878 100000 6 dout0[5]
port 222 nsew signal input
rlabel metal2 s 91926 99200 91982 100000 6 dout0[60]
port 223 nsew signal input
rlabel metal2 s 92754 99200 92810 100000 6 dout0[61]
port 224 nsew signal input
rlabel metal2 s 93582 99200 93638 100000 6 dout0[62]
port 225 nsew signal input
rlabel metal2 s 94410 99200 94466 100000 6 dout0[63]
port 226 nsew signal input
rlabel metal2 s 45650 99200 45706 100000 6 dout0[6]
port 227 nsew signal input
rlabel metal2 s 46570 99200 46626 100000 6 dout0[7]
port 228 nsew signal input
rlabel metal2 s 47398 99200 47454 100000 6 dout0[8]
port 229 nsew signal input
rlabel metal2 s 48226 99200 48282 100000 6 dout0[9]
port 230 nsew signal input
rlabel metal2 s 103886 99200 103942 100000 6 dout1[0]
port 231 nsew signal input
rlabel metal2 s 112442 99200 112498 100000 6 dout1[10]
port 232 nsew signal input
rlabel metal2 s 113270 99200 113326 100000 6 dout1[11]
port 233 nsew signal input
rlabel metal2 s 114098 99200 114154 100000 6 dout1[12]
port 234 nsew signal input
rlabel metal2 s 115018 99200 115074 100000 6 dout1[13]
port 235 nsew signal input
rlabel metal2 s 115846 99200 115902 100000 6 dout1[14]
port 236 nsew signal input
rlabel metal2 s 116674 99200 116730 100000 6 dout1[15]
port 237 nsew signal input
rlabel metal2 s 117594 99200 117650 100000 6 dout1[16]
port 238 nsew signal input
rlabel metal2 s 118422 99200 118478 100000 6 dout1[17]
port 239 nsew signal input
rlabel metal2 s 119250 99200 119306 100000 6 dout1[18]
port 240 nsew signal input
rlabel metal2 s 120078 99200 120134 100000 6 dout1[19]
port 241 nsew signal input
rlabel metal2 s 104714 99200 104770 100000 6 dout1[1]
port 242 nsew signal input
rlabel metal2 s 120998 99200 121054 100000 6 dout1[20]
port 243 nsew signal input
rlabel metal2 s 121826 99200 121882 100000 6 dout1[21]
port 244 nsew signal input
rlabel metal2 s 122654 99200 122710 100000 6 dout1[22]
port 245 nsew signal input
rlabel metal2 s 123574 99200 123630 100000 6 dout1[23]
port 246 nsew signal input
rlabel metal2 s 124402 99200 124458 100000 6 dout1[24]
port 247 nsew signal input
rlabel metal2 s 125230 99200 125286 100000 6 dout1[25]
port 248 nsew signal input
rlabel metal2 s 126150 99200 126206 100000 6 dout1[26]
port 249 nsew signal input
rlabel metal2 s 126978 99200 127034 100000 6 dout1[27]
port 250 nsew signal input
rlabel metal2 s 127806 99200 127862 100000 6 dout1[28]
port 251 nsew signal input
rlabel metal2 s 128634 99200 128690 100000 6 dout1[29]
port 252 nsew signal input
rlabel metal2 s 105542 99200 105598 100000 6 dout1[2]
port 253 nsew signal input
rlabel metal2 s 129554 99200 129610 100000 6 dout1[30]
port 254 nsew signal input
rlabel metal2 s 130382 99200 130438 100000 6 dout1[31]
port 255 nsew signal input
rlabel metal2 s 131210 99200 131266 100000 6 dout1[32]
port 256 nsew signal input
rlabel metal2 s 132130 99200 132186 100000 6 dout1[33]
port 257 nsew signal input
rlabel metal2 s 132958 99200 133014 100000 6 dout1[34]
port 258 nsew signal input
rlabel metal2 s 133786 99200 133842 100000 6 dout1[35]
port 259 nsew signal input
rlabel metal2 s 134706 99200 134762 100000 6 dout1[36]
port 260 nsew signal input
rlabel metal2 s 135534 99200 135590 100000 6 dout1[37]
port 261 nsew signal input
rlabel metal2 s 136362 99200 136418 100000 6 dout1[38]
port 262 nsew signal input
rlabel metal2 s 137190 99200 137246 100000 6 dout1[39]
port 263 nsew signal input
rlabel metal2 s 106462 99200 106518 100000 6 dout1[3]
port 264 nsew signal input
rlabel metal2 s 138110 99200 138166 100000 6 dout1[40]
port 265 nsew signal input
rlabel metal2 s 138938 99200 138994 100000 6 dout1[41]
port 266 nsew signal input
rlabel metal2 s 139766 99200 139822 100000 6 dout1[42]
port 267 nsew signal input
rlabel metal2 s 140686 99200 140742 100000 6 dout1[43]
port 268 nsew signal input
rlabel metal2 s 141514 99200 141570 100000 6 dout1[44]
port 269 nsew signal input
rlabel metal2 s 142342 99200 142398 100000 6 dout1[45]
port 270 nsew signal input
rlabel metal2 s 143262 99200 143318 100000 6 dout1[46]
port 271 nsew signal input
rlabel metal2 s 144090 99200 144146 100000 6 dout1[47]
port 272 nsew signal input
rlabel metal2 s 144918 99200 144974 100000 6 dout1[48]
port 273 nsew signal input
rlabel metal2 s 145746 99200 145802 100000 6 dout1[49]
port 274 nsew signal input
rlabel metal2 s 107290 99200 107346 100000 6 dout1[4]
port 275 nsew signal input
rlabel metal2 s 146666 99200 146722 100000 6 dout1[50]
port 276 nsew signal input
rlabel metal2 s 147494 99200 147550 100000 6 dout1[51]
port 277 nsew signal input
rlabel metal2 s 148322 99200 148378 100000 6 dout1[52]
port 278 nsew signal input
rlabel metal2 s 149242 99200 149298 100000 6 dout1[53]
port 279 nsew signal input
rlabel metal2 s 150070 99200 150126 100000 6 dout1[54]
port 280 nsew signal input
rlabel metal2 s 150898 99200 150954 100000 6 dout1[55]
port 281 nsew signal input
rlabel metal2 s 151818 99200 151874 100000 6 dout1[56]
port 282 nsew signal input
rlabel metal2 s 152646 99200 152702 100000 6 dout1[57]
port 283 nsew signal input
rlabel metal2 s 153474 99200 153530 100000 6 dout1[58]
port 284 nsew signal input
rlabel metal2 s 154302 99200 154358 100000 6 dout1[59]
port 285 nsew signal input
rlabel metal2 s 108118 99200 108174 100000 6 dout1[5]
port 286 nsew signal input
rlabel metal2 s 155222 99200 155278 100000 6 dout1[60]
port 287 nsew signal input
rlabel metal2 s 156050 99200 156106 100000 6 dout1[61]
port 288 nsew signal input
rlabel metal2 s 156878 99200 156934 100000 6 dout1[62]
port 289 nsew signal input
rlabel metal2 s 157798 99200 157854 100000 6 dout1[63]
port 290 nsew signal input
rlabel metal2 s 109038 99200 109094 100000 6 dout1[6]
port 291 nsew signal input
rlabel metal2 s 109866 99200 109922 100000 6 dout1[7]
port 292 nsew signal input
rlabel metal2 s 110694 99200 110750 100000 6 dout1[8]
port 293 nsew signal input
rlabel metal2 s 111522 99200 111578 100000 6 dout1[9]
port 294 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 jtag_tck
port 295 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 jtag_tdi
port 296 nsew signal input
rlabel metal3 s 159200 99016 160000 99136 6 jtag_tdo
port 297 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 jtag_tms
port 298 nsew signal input
rlabel metal3 s 159200 51008 160000 51128 6 localMemory_wb_ack_o
port 299 nsew signal output
rlabel metal3 s 159200 54000 160000 54120 6 localMemory_wb_adr_i[0]
port 300 nsew signal input
rlabel metal3 s 159200 70592 160000 70712 6 localMemory_wb_adr_i[10]
port 301 nsew signal input
rlabel metal3 s 159200 72088 160000 72208 6 localMemory_wb_adr_i[11]
port 302 nsew signal input
rlabel metal3 s 159200 73584 160000 73704 6 localMemory_wb_adr_i[12]
port 303 nsew signal input
rlabel metal3 s 159200 75080 160000 75200 6 localMemory_wb_adr_i[13]
port 304 nsew signal input
rlabel metal3 s 159200 76576 160000 76696 6 localMemory_wb_adr_i[14]
port 305 nsew signal input
rlabel metal3 s 159200 77936 160000 78056 6 localMemory_wb_adr_i[15]
port 306 nsew signal input
rlabel metal3 s 159200 79432 160000 79552 6 localMemory_wb_adr_i[16]
port 307 nsew signal input
rlabel metal3 s 159200 80928 160000 81048 6 localMemory_wb_adr_i[17]
port 308 nsew signal input
rlabel metal3 s 159200 82424 160000 82544 6 localMemory_wb_adr_i[18]
port 309 nsew signal input
rlabel metal3 s 159200 83920 160000 84040 6 localMemory_wb_adr_i[19]
port 310 nsew signal input
rlabel metal3 s 159200 55904 160000 56024 6 localMemory_wb_adr_i[1]
port 311 nsew signal input
rlabel metal3 s 159200 85280 160000 85400 6 localMemory_wb_adr_i[20]
port 312 nsew signal input
rlabel metal3 s 159200 86776 160000 86896 6 localMemory_wb_adr_i[21]
port 313 nsew signal input
rlabel metal3 s 159200 88272 160000 88392 6 localMemory_wb_adr_i[22]
port 314 nsew signal input
rlabel metal3 s 159200 89768 160000 89888 6 localMemory_wb_adr_i[23]
port 315 nsew signal input
rlabel metal3 s 159200 57944 160000 58064 6 localMemory_wb_adr_i[2]
port 316 nsew signal input
rlabel metal3 s 159200 59848 160000 59968 6 localMemory_wb_adr_i[3]
port 317 nsew signal input
rlabel metal3 s 159200 61752 160000 61872 6 localMemory_wb_adr_i[4]
port 318 nsew signal input
rlabel metal3 s 159200 63248 160000 63368 6 localMemory_wb_adr_i[5]
port 319 nsew signal input
rlabel metal3 s 159200 64744 160000 64864 6 localMemory_wb_adr_i[6]
port 320 nsew signal input
rlabel metal3 s 159200 66240 160000 66360 6 localMemory_wb_adr_i[7]
port 321 nsew signal input
rlabel metal3 s 159200 67736 160000 67856 6 localMemory_wb_adr_i[8]
port 322 nsew signal input
rlabel metal3 s 159200 69232 160000 69352 6 localMemory_wb_adr_i[9]
port 323 nsew signal input
rlabel metal3 s 159200 51552 160000 51672 6 localMemory_wb_cyc_i
port 324 nsew signal input
rlabel metal3 s 159200 54408 160000 54528 6 localMemory_wb_data_i[0]
port 325 nsew signal input
rlabel metal3 s 159200 71136 160000 71256 6 localMemory_wb_data_i[10]
port 326 nsew signal input
rlabel metal3 s 159200 72632 160000 72752 6 localMemory_wb_data_i[11]
port 327 nsew signal input
rlabel metal3 s 159200 74128 160000 74248 6 localMemory_wb_data_i[12]
port 328 nsew signal input
rlabel metal3 s 159200 75488 160000 75608 6 localMemory_wb_data_i[13]
port 329 nsew signal input
rlabel metal3 s 159200 76984 160000 77104 6 localMemory_wb_data_i[14]
port 330 nsew signal input
rlabel metal3 s 159200 78480 160000 78600 6 localMemory_wb_data_i[15]
port 331 nsew signal input
rlabel metal3 s 159200 79976 160000 80096 6 localMemory_wb_data_i[16]
port 332 nsew signal input
rlabel metal3 s 159200 81472 160000 81592 6 localMemory_wb_data_i[17]
port 333 nsew signal input
rlabel metal3 s 159200 82832 160000 82952 6 localMemory_wb_data_i[18]
port 334 nsew signal input
rlabel metal3 s 159200 84328 160000 84448 6 localMemory_wb_data_i[19]
port 335 nsew signal input
rlabel metal3 s 159200 56448 160000 56568 6 localMemory_wb_data_i[1]
port 336 nsew signal input
rlabel metal3 s 159200 85824 160000 85944 6 localMemory_wb_data_i[20]
port 337 nsew signal input
rlabel metal3 s 159200 87320 160000 87440 6 localMemory_wb_data_i[21]
port 338 nsew signal input
rlabel metal3 s 159200 88816 160000 88936 6 localMemory_wb_data_i[22]
port 339 nsew signal input
rlabel metal3 s 159200 90176 160000 90296 6 localMemory_wb_data_i[23]
port 340 nsew signal input
rlabel metal3 s 159200 91264 160000 91384 6 localMemory_wb_data_i[24]
port 341 nsew signal input
rlabel metal3 s 159200 92216 160000 92336 6 localMemory_wb_data_i[25]
port 342 nsew signal input
rlabel metal3 s 159200 93168 160000 93288 6 localMemory_wb_data_i[26]
port 343 nsew signal input
rlabel metal3 s 159200 94120 160000 94240 6 localMemory_wb_data_i[27]
port 344 nsew signal input
rlabel metal3 s 159200 95072 160000 95192 6 localMemory_wb_data_i[28]
port 345 nsew signal input
rlabel metal3 s 159200 96160 160000 96280 6 localMemory_wb_data_i[29]
port 346 nsew signal input
rlabel metal3 s 159200 58352 160000 58472 6 localMemory_wb_data_i[2]
port 347 nsew signal input
rlabel metal3 s 159200 97112 160000 97232 6 localMemory_wb_data_i[30]
port 348 nsew signal input
rlabel metal3 s 159200 98064 160000 98184 6 localMemory_wb_data_i[31]
port 349 nsew signal input
rlabel metal3 s 159200 60392 160000 60512 6 localMemory_wb_data_i[3]
port 350 nsew signal input
rlabel metal3 s 159200 62296 160000 62416 6 localMemory_wb_data_i[4]
port 351 nsew signal input
rlabel metal3 s 159200 63792 160000 63912 6 localMemory_wb_data_i[5]
port 352 nsew signal input
rlabel metal3 s 159200 65288 160000 65408 6 localMemory_wb_data_i[6]
port 353 nsew signal input
rlabel metal3 s 159200 66784 160000 66904 6 localMemory_wb_data_i[7]
port 354 nsew signal input
rlabel metal3 s 159200 68144 160000 68264 6 localMemory_wb_data_i[8]
port 355 nsew signal input
rlabel metal3 s 159200 69640 160000 69760 6 localMemory_wb_data_i[9]
port 356 nsew signal input
rlabel metal3 s 159200 54952 160000 55072 6 localMemory_wb_data_o[0]
port 357 nsew signal output
rlabel metal3 s 159200 71680 160000 71800 6 localMemory_wb_data_o[10]
port 358 nsew signal output
rlabel metal3 s 159200 73040 160000 73160 6 localMemory_wb_data_o[11]
port 359 nsew signal output
rlabel metal3 s 159200 74536 160000 74656 6 localMemory_wb_data_o[12]
port 360 nsew signal output
rlabel metal3 s 159200 76032 160000 76152 6 localMemory_wb_data_o[13]
port 361 nsew signal output
rlabel metal3 s 159200 77528 160000 77648 6 localMemory_wb_data_o[14]
port 362 nsew signal output
rlabel metal3 s 159200 79024 160000 79144 6 localMemory_wb_data_o[15]
port 363 nsew signal output
rlabel metal3 s 159200 80384 160000 80504 6 localMemory_wb_data_o[16]
port 364 nsew signal output
rlabel metal3 s 159200 81880 160000 82000 6 localMemory_wb_data_o[17]
port 365 nsew signal output
rlabel metal3 s 159200 83376 160000 83496 6 localMemory_wb_data_o[18]
port 366 nsew signal output
rlabel metal3 s 159200 84872 160000 84992 6 localMemory_wb_data_o[19]
port 367 nsew signal output
rlabel metal3 s 159200 56856 160000 56976 6 localMemory_wb_data_o[1]
port 368 nsew signal output
rlabel metal3 s 159200 86368 160000 86488 6 localMemory_wb_data_o[20]
port 369 nsew signal output
rlabel metal3 s 159200 87728 160000 87848 6 localMemory_wb_data_o[21]
port 370 nsew signal output
rlabel metal3 s 159200 89224 160000 89344 6 localMemory_wb_data_o[22]
port 371 nsew signal output
rlabel metal3 s 159200 90720 160000 90840 6 localMemory_wb_data_o[23]
port 372 nsew signal output
rlabel metal3 s 159200 91672 160000 91792 6 localMemory_wb_data_o[24]
port 373 nsew signal output
rlabel metal3 s 159200 92624 160000 92744 6 localMemory_wb_data_o[25]
port 374 nsew signal output
rlabel metal3 s 159200 93712 160000 93832 6 localMemory_wb_data_o[26]
port 375 nsew signal output
rlabel metal3 s 159200 94664 160000 94784 6 localMemory_wb_data_o[27]
port 376 nsew signal output
rlabel metal3 s 159200 95616 160000 95736 6 localMemory_wb_data_o[28]
port 377 nsew signal output
rlabel metal3 s 159200 96568 160000 96688 6 localMemory_wb_data_o[29]
port 378 nsew signal output
rlabel metal3 s 159200 58896 160000 59016 6 localMemory_wb_data_o[2]
port 379 nsew signal output
rlabel metal3 s 159200 97520 160000 97640 6 localMemory_wb_data_o[30]
port 380 nsew signal output
rlabel metal3 s 159200 98608 160000 98728 6 localMemory_wb_data_o[31]
port 381 nsew signal output
rlabel metal3 s 159200 60800 160000 60920 6 localMemory_wb_data_o[3]
port 382 nsew signal output
rlabel metal3 s 159200 62840 160000 62960 6 localMemory_wb_data_o[4]
port 383 nsew signal output
rlabel metal3 s 159200 64200 160000 64320 6 localMemory_wb_data_o[5]
port 384 nsew signal output
rlabel metal3 s 159200 65696 160000 65816 6 localMemory_wb_data_o[6]
port 385 nsew signal output
rlabel metal3 s 159200 67192 160000 67312 6 localMemory_wb_data_o[7]
port 386 nsew signal output
rlabel metal3 s 159200 68688 160000 68808 6 localMemory_wb_data_o[8]
port 387 nsew signal output
rlabel metal3 s 159200 70184 160000 70304 6 localMemory_wb_data_o[9]
port 388 nsew signal output
rlabel metal3 s 159200 51960 160000 52080 6 localMemory_wb_error_o
port 389 nsew signal output
rlabel metal3 s 159200 55496 160000 55616 6 localMemory_wb_sel_i[0]
port 390 nsew signal input
rlabel metal3 s 159200 57400 160000 57520 6 localMemory_wb_sel_i[1]
port 391 nsew signal input
rlabel metal3 s 159200 59304 160000 59424 6 localMemory_wb_sel_i[2]
port 392 nsew signal input
rlabel metal3 s 159200 61344 160000 61464 6 localMemory_wb_sel_i[3]
port 393 nsew signal input
rlabel metal3 s 159200 52504 160000 52624 6 localMemory_wb_stall_o
port 394 nsew signal output
rlabel metal3 s 159200 53048 160000 53168 6 localMemory_wb_stb_i
port 395 nsew signal input
rlabel metal3 s 159200 53456 160000 53576 6 localMemory_wb_we_i
port 396 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 manufacturerID[0]
port 397 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 manufacturerID[10]
port 398 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 manufacturerID[1]
port 399 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 manufacturerID[2]
port 400 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 manufacturerID[3]
port 401 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 manufacturerID[4]
port 402 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 manufacturerID[5]
port 403 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 manufacturerID[6]
port 404 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 manufacturerID[7]
port 405 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 manufacturerID[8]
port 406 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 manufacturerID[9]
port 407 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 partID[0]
port 408 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 partID[10]
port 409 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 partID[11]
port 410 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 partID[12]
port 411 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 partID[13]
port 412 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 partID[14]
port 413 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 partID[15]
port 414 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 partID[1]
port 415 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 partID[2]
port 416 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 partID[3]
port 417 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 partID[4]
port 418 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 partID[5]
port 419 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 partID[6]
port 420 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 partID[7]
port 421 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 partID[8]
port 422 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 partID[9]
port 423 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 probe_errorCode[0]
port 424 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 probe_errorCode[1]
port 425 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 probe_errorCode[2]
port 426 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 probe_errorCode[3]
port 427 nsew signal output
rlabel metal3 s 0 824 800 944 6 probe_isBranch
port 428 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 probe_isCompressed
port 429 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 probe_isLoad
port 430 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 probe_isStore
port 431 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 probe_jtagInstruction[0]
port 432 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 probe_jtagInstruction[1]
port 433 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 probe_jtagInstruction[2]
port 434 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 probe_jtagInstruction[3]
port 435 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 probe_jtagInstruction[4]
port 436 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 probe_opcode[0]
port 437 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 probe_opcode[1]
port 438 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 probe_opcode[2]
port 439 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 probe_opcode[3]
port 440 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 probe_opcode[4]
port 441 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 probe_opcode[5]
port 442 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 probe_opcode[6]
port 443 nsew signal output
rlabel metal3 s 0 14832 800 14952 6 probe_programCounter[0]
port 444 nsew signal output
rlabel metal3 s 0 58624 800 58744 6 probe_programCounter[10]
port 445 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 probe_programCounter[11]
port 446 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 probe_programCounter[12]
port 447 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 probe_programCounter[13]
port 448 nsew signal output
rlabel metal3 s 0 65696 800 65816 6 probe_programCounter[14]
port 449 nsew signal output
rlabel metal3 s 0 67464 800 67584 6 probe_programCounter[15]
port 450 nsew signal output
rlabel metal3 s 0 69096 800 69216 6 probe_programCounter[16]
port 451 nsew signal output
rlabel metal3 s 0 70864 800 70984 6 probe_programCounter[17]
port 452 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 probe_programCounter[18]
port 453 nsew signal output
rlabel metal3 s 0 74400 800 74520 6 probe_programCounter[19]
port 454 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 probe_programCounter[1]
port 455 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 probe_programCounter[20]
port 456 nsew signal output
rlabel metal3 s 0 77936 800 78056 6 probe_programCounter[21]
port 457 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 probe_programCounter[22]
port 458 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 probe_programCounter[23]
port 459 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 probe_programCounter[24]
port 460 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 probe_programCounter[25]
port 461 nsew signal output
rlabel metal3 s 0 86640 800 86760 6 probe_programCounter[26]
port 462 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 probe_programCounter[27]
port 463 nsew signal output
rlabel metal3 s 0 90176 800 90296 6 probe_programCounter[28]
port 464 nsew signal output
rlabel metal3 s 0 91944 800 92064 6 probe_programCounter[29]
port 465 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 probe_programCounter[2]
port 466 nsew signal output
rlabel metal3 s 0 93712 800 93832 6 probe_programCounter[30]
port 467 nsew signal output
rlabel metal3 s 0 95480 800 95600 6 probe_programCounter[31]
port 468 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 probe_programCounter[3]
port 469 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 probe_programCounter[4]
port 470 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 probe_programCounter[5]
port 471 nsew signal output
rlabel metal3 s 0 51552 800 51672 6 probe_programCounter[6]
port 472 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 probe_programCounter[7]
port 473 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 probe_programCounter[8]
port 474 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 probe_programCounter[9]
port 475 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 probe_state[0]
port 476 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 probe_state[1]
port 477 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 probe_takeBranch
port 478 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal2 s 138478 0 138534 800 6 versionID[0]
port 480 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 versionID[1]
port 481 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 versionID[2]
port 482 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 versionID[3]
port 483 nsew signal input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal3 s 159200 144 160000 264 6 wb_clk_i
port 485 nsew signal input
rlabel metal3 s 159200 552 160000 672 6 wb_rst_i
port 486 nsew signal input
rlabel metal2 s 1214 99200 1270 100000 6 web0
port 487 nsew signal output
rlabel metal2 s 2042 99200 2098 100000 6 wmask0[0]
port 488 nsew signal output
rlabel metal2 s 2870 99200 2926 100000 6 wmask0[1]
port 489 nsew signal output
rlabel metal2 s 3790 99200 3846 100000 6 wmask0[2]
port 490 nsew signal output
rlabel metal2 s 4618 99200 4674 100000 6 wmask0[3]
port 491 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 160000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7028258
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/ExperiarCore/results/signoff/ExperiarCore.magic.gds
string GDS_START 492612
<< end >>

