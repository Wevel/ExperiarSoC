magic
tech sky130A
magscale 1 2
timestamp 1652907394
<< obsli1 >>
rect 1104 2159 158884 97393
<< obsm1 >>
rect 382 1572 159514 98048
<< metal2 >>
rect 386 99200 442 100000
rect 1214 99200 1270 100000
rect 2042 99200 2098 100000
rect 2962 99200 3018 100000
rect 3790 99200 3846 100000
rect 4618 99200 4674 100000
rect 5538 99200 5594 100000
rect 6366 99200 6422 100000
rect 7194 99200 7250 100000
rect 8114 99200 8170 100000
rect 8942 99200 8998 100000
rect 9770 99200 9826 100000
rect 10690 99200 10746 100000
rect 11518 99200 11574 100000
rect 12346 99200 12402 100000
rect 13266 99200 13322 100000
rect 14094 99200 14150 100000
rect 14922 99200 14978 100000
rect 15842 99200 15898 100000
rect 16670 99200 16726 100000
rect 17498 99200 17554 100000
rect 18418 99200 18474 100000
rect 19246 99200 19302 100000
rect 20166 99200 20222 100000
rect 20994 99200 21050 100000
rect 21822 99200 21878 100000
rect 22742 99200 22798 100000
rect 23570 99200 23626 100000
rect 24398 99200 24454 100000
rect 25318 99200 25374 100000
rect 26146 99200 26202 100000
rect 26974 99200 27030 100000
rect 27894 99200 27950 100000
rect 28722 99200 28778 100000
rect 29550 99200 29606 100000
rect 30470 99200 30526 100000
rect 31298 99200 31354 100000
rect 32126 99200 32182 100000
rect 33046 99200 33102 100000
rect 33874 99200 33930 100000
rect 34702 99200 34758 100000
rect 35622 99200 35678 100000
rect 36450 99200 36506 100000
rect 37370 99200 37426 100000
rect 38198 99200 38254 100000
rect 39026 99200 39082 100000
rect 39946 99200 40002 100000
rect 40774 99200 40830 100000
rect 41602 99200 41658 100000
rect 42522 99200 42578 100000
rect 43350 99200 43406 100000
rect 44178 99200 44234 100000
rect 45098 99200 45154 100000
rect 45926 99200 45982 100000
rect 46754 99200 46810 100000
rect 47674 99200 47730 100000
rect 48502 99200 48558 100000
rect 49330 99200 49386 100000
rect 50250 99200 50306 100000
rect 51078 99200 51134 100000
rect 51906 99200 51962 100000
rect 52826 99200 52882 100000
rect 53654 99200 53710 100000
rect 54574 99200 54630 100000
rect 55402 99200 55458 100000
rect 56230 99200 56286 100000
rect 57150 99200 57206 100000
rect 57978 99200 58034 100000
rect 58806 99200 58862 100000
rect 59726 99200 59782 100000
rect 60554 99200 60610 100000
rect 61382 99200 61438 100000
rect 62302 99200 62358 100000
rect 63130 99200 63186 100000
rect 63958 99200 64014 100000
rect 64878 99200 64934 100000
rect 65706 99200 65762 100000
rect 66534 99200 66590 100000
rect 67454 99200 67510 100000
rect 68282 99200 68338 100000
rect 69110 99200 69166 100000
rect 70030 99200 70086 100000
rect 70858 99200 70914 100000
rect 71778 99200 71834 100000
rect 72606 99200 72662 100000
rect 73434 99200 73490 100000
rect 74354 99200 74410 100000
rect 75182 99200 75238 100000
rect 76010 99200 76066 100000
rect 76930 99200 76986 100000
rect 77758 99200 77814 100000
rect 78586 99200 78642 100000
rect 79506 99200 79562 100000
rect 80334 99200 80390 100000
rect 81162 99200 81218 100000
rect 82082 99200 82138 100000
rect 82910 99200 82966 100000
rect 83738 99200 83794 100000
rect 84658 99200 84714 100000
rect 85486 99200 85542 100000
rect 86314 99200 86370 100000
rect 87234 99200 87290 100000
rect 88062 99200 88118 100000
rect 88890 99200 88946 100000
rect 89810 99200 89866 100000
rect 90638 99200 90694 100000
rect 91558 99200 91614 100000
rect 92386 99200 92442 100000
rect 93214 99200 93270 100000
rect 94134 99200 94190 100000
rect 94962 99200 95018 100000
rect 95790 99200 95846 100000
rect 96710 99200 96766 100000
rect 97538 99200 97594 100000
rect 98366 99200 98422 100000
rect 99286 99200 99342 100000
rect 100114 99200 100170 100000
rect 100942 99200 100998 100000
rect 101862 99200 101918 100000
rect 102690 99200 102746 100000
rect 103518 99200 103574 100000
rect 104438 99200 104494 100000
rect 105266 99200 105322 100000
rect 106094 99200 106150 100000
rect 107014 99200 107070 100000
rect 107842 99200 107898 100000
rect 108762 99200 108818 100000
rect 109590 99200 109646 100000
rect 110418 99200 110474 100000
rect 111338 99200 111394 100000
rect 112166 99200 112222 100000
rect 112994 99200 113050 100000
rect 113914 99200 113970 100000
rect 114742 99200 114798 100000
rect 115570 99200 115626 100000
rect 116490 99200 116546 100000
rect 117318 99200 117374 100000
rect 118146 99200 118202 100000
rect 119066 99200 119122 100000
rect 119894 99200 119950 100000
rect 120722 99200 120778 100000
rect 121642 99200 121698 100000
rect 122470 99200 122526 100000
rect 123298 99200 123354 100000
rect 124218 99200 124274 100000
rect 125046 99200 125102 100000
rect 125966 99200 126022 100000
rect 126794 99200 126850 100000
rect 127622 99200 127678 100000
rect 128542 99200 128598 100000
rect 129370 99200 129426 100000
rect 130198 99200 130254 100000
rect 131118 99200 131174 100000
rect 131946 99200 132002 100000
rect 132774 99200 132830 100000
rect 133694 99200 133750 100000
rect 134522 99200 134578 100000
rect 135350 99200 135406 100000
rect 136270 99200 136326 100000
rect 137098 99200 137154 100000
rect 137926 99200 137982 100000
rect 138846 99200 138902 100000
rect 139674 99200 139730 100000
rect 140502 99200 140558 100000
rect 141422 99200 141478 100000
rect 142250 99200 142306 100000
rect 143170 99200 143226 100000
rect 143998 99200 144054 100000
rect 144826 99200 144882 100000
rect 145746 99200 145802 100000
rect 146574 99200 146630 100000
rect 147402 99200 147458 100000
rect 148322 99200 148378 100000
rect 149150 99200 149206 100000
rect 149978 99200 150034 100000
rect 150898 99200 150954 100000
rect 151726 99200 151782 100000
rect 152554 99200 152610 100000
rect 153474 99200 153530 100000
rect 154302 99200 154358 100000
rect 155130 99200 155186 100000
rect 156050 99200 156106 100000
rect 156878 99200 156934 100000
rect 157706 99200 157762 100000
rect 158626 99200 158682 100000
rect 159454 99200 159510 100000
rect 1950 0 2006 800
rect 5906 0 5962 800
rect 9862 0 9918 800
rect 13910 0 13966 800
rect 17866 0 17922 800
rect 21914 0 21970 800
rect 25870 0 25926 800
rect 29918 0 29974 800
rect 33874 0 33930 800
rect 37922 0 37978 800
rect 41878 0 41934 800
rect 45926 0 45982 800
rect 49882 0 49938 800
rect 53930 0 53986 800
rect 57886 0 57942 800
rect 61934 0 61990 800
rect 65890 0 65946 800
rect 69938 0 69994 800
rect 73894 0 73950 800
rect 77942 0 77998 800
rect 81898 0 81954 800
rect 85854 0 85910 800
rect 89902 0 89958 800
rect 93858 0 93914 800
rect 97906 0 97962 800
rect 101862 0 101918 800
rect 105910 0 105966 800
rect 109866 0 109922 800
rect 113914 0 113970 800
rect 117870 0 117926 800
rect 121918 0 121974 800
rect 125874 0 125930 800
rect 129922 0 129978 800
rect 133878 0 133934 800
rect 137926 0 137982 800
rect 141882 0 141938 800
rect 145930 0 145986 800
rect 149886 0 149942 800
rect 153934 0 153990 800
rect 157890 0 157946 800
<< obsm2 >>
rect 498 99144 1158 99657
rect 1326 99144 1986 99657
rect 2154 99144 2906 99657
rect 3074 99144 3734 99657
rect 3902 99144 4562 99657
rect 4730 99144 5482 99657
rect 5650 99144 6310 99657
rect 6478 99144 7138 99657
rect 7306 99144 8058 99657
rect 8226 99144 8886 99657
rect 9054 99144 9714 99657
rect 9882 99144 10634 99657
rect 10802 99144 11462 99657
rect 11630 99144 12290 99657
rect 12458 99144 13210 99657
rect 13378 99144 14038 99657
rect 14206 99144 14866 99657
rect 15034 99144 15786 99657
rect 15954 99144 16614 99657
rect 16782 99144 17442 99657
rect 17610 99144 18362 99657
rect 18530 99144 19190 99657
rect 19358 99144 20110 99657
rect 20278 99144 20938 99657
rect 21106 99144 21766 99657
rect 21934 99144 22686 99657
rect 22854 99144 23514 99657
rect 23682 99144 24342 99657
rect 24510 99144 25262 99657
rect 25430 99144 26090 99657
rect 26258 99144 26918 99657
rect 27086 99144 27838 99657
rect 28006 99144 28666 99657
rect 28834 99144 29494 99657
rect 29662 99144 30414 99657
rect 30582 99144 31242 99657
rect 31410 99144 32070 99657
rect 32238 99144 32990 99657
rect 33158 99144 33818 99657
rect 33986 99144 34646 99657
rect 34814 99144 35566 99657
rect 35734 99144 36394 99657
rect 36562 99144 37314 99657
rect 37482 99144 38142 99657
rect 38310 99144 38970 99657
rect 39138 99144 39890 99657
rect 40058 99144 40718 99657
rect 40886 99144 41546 99657
rect 41714 99144 42466 99657
rect 42634 99144 43294 99657
rect 43462 99144 44122 99657
rect 44290 99144 45042 99657
rect 45210 99144 45870 99657
rect 46038 99144 46698 99657
rect 46866 99144 47618 99657
rect 47786 99144 48446 99657
rect 48614 99144 49274 99657
rect 49442 99144 50194 99657
rect 50362 99144 51022 99657
rect 51190 99144 51850 99657
rect 52018 99144 52770 99657
rect 52938 99144 53598 99657
rect 53766 99144 54518 99657
rect 54686 99144 55346 99657
rect 55514 99144 56174 99657
rect 56342 99144 57094 99657
rect 57262 99144 57922 99657
rect 58090 99144 58750 99657
rect 58918 99144 59670 99657
rect 59838 99144 60498 99657
rect 60666 99144 61326 99657
rect 61494 99144 62246 99657
rect 62414 99144 63074 99657
rect 63242 99144 63902 99657
rect 64070 99144 64822 99657
rect 64990 99144 65650 99657
rect 65818 99144 66478 99657
rect 66646 99144 67398 99657
rect 67566 99144 68226 99657
rect 68394 99144 69054 99657
rect 69222 99144 69974 99657
rect 70142 99144 70802 99657
rect 70970 99144 71722 99657
rect 71890 99144 72550 99657
rect 72718 99144 73378 99657
rect 73546 99144 74298 99657
rect 74466 99144 75126 99657
rect 75294 99144 75954 99657
rect 76122 99144 76874 99657
rect 77042 99144 77702 99657
rect 77870 99144 78530 99657
rect 78698 99144 79450 99657
rect 79618 99144 80278 99657
rect 80446 99144 81106 99657
rect 81274 99144 82026 99657
rect 82194 99144 82854 99657
rect 83022 99144 83682 99657
rect 83850 99144 84602 99657
rect 84770 99144 85430 99657
rect 85598 99144 86258 99657
rect 86426 99144 87178 99657
rect 87346 99144 88006 99657
rect 88174 99144 88834 99657
rect 89002 99144 89754 99657
rect 89922 99144 90582 99657
rect 90750 99144 91502 99657
rect 91670 99144 92330 99657
rect 92498 99144 93158 99657
rect 93326 99144 94078 99657
rect 94246 99144 94906 99657
rect 95074 99144 95734 99657
rect 95902 99144 96654 99657
rect 96822 99144 97482 99657
rect 97650 99144 98310 99657
rect 98478 99144 99230 99657
rect 99398 99144 100058 99657
rect 100226 99144 100886 99657
rect 101054 99144 101806 99657
rect 101974 99144 102634 99657
rect 102802 99144 103462 99657
rect 103630 99144 104382 99657
rect 104550 99144 105210 99657
rect 105378 99144 106038 99657
rect 106206 99144 106958 99657
rect 107126 99144 107786 99657
rect 107954 99144 108706 99657
rect 108874 99144 109534 99657
rect 109702 99144 110362 99657
rect 110530 99144 111282 99657
rect 111450 99144 112110 99657
rect 112278 99144 112938 99657
rect 113106 99144 113858 99657
rect 114026 99144 114686 99657
rect 114854 99144 115514 99657
rect 115682 99144 116434 99657
rect 116602 99144 117262 99657
rect 117430 99144 118090 99657
rect 118258 99144 119010 99657
rect 119178 99144 119838 99657
rect 120006 99144 120666 99657
rect 120834 99144 121586 99657
rect 121754 99144 122414 99657
rect 122582 99144 123242 99657
rect 123410 99144 124162 99657
rect 124330 99144 124990 99657
rect 125158 99144 125910 99657
rect 126078 99144 126738 99657
rect 126906 99144 127566 99657
rect 127734 99144 128486 99657
rect 128654 99144 129314 99657
rect 129482 99144 130142 99657
rect 130310 99144 131062 99657
rect 131230 99144 131890 99657
rect 132058 99144 132718 99657
rect 132886 99144 133638 99657
rect 133806 99144 134466 99657
rect 134634 99144 135294 99657
rect 135462 99144 136214 99657
rect 136382 99144 137042 99657
rect 137210 99144 137870 99657
rect 138038 99144 138790 99657
rect 138958 99144 139618 99657
rect 139786 99144 140446 99657
rect 140614 99144 141366 99657
rect 141534 99144 142194 99657
rect 142362 99144 143114 99657
rect 143282 99144 143942 99657
rect 144110 99144 144770 99657
rect 144938 99144 145690 99657
rect 145858 99144 146518 99657
rect 146686 99144 147346 99657
rect 147514 99144 148266 99657
rect 148434 99144 149094 99657
rect 149262 99144 149922 99657
rect 150090 99144 150842 99657
rect 151010 99144 151670 99657
rect 151838 99144 152498 99657
rect 152666 99144 153418 99657
rect 153586 99144 154246 99657
rect 154414 99144 155074 99657
rect 155242 99144 155994 99657
rect 156162 99144 156822 99657
rect 156990 99144 157650 99657
rect 157818 99144 158570 99657
rect 158738 99144 159398 99657
rect 388 856 159508 99144
rect 388 575 1894 856
rect 2062 575 5850 856
rect 6018 575 9806 856
rect 9974 575 13854 856
rect 14022 575 17810 856
rect 17978 575 21858 856
rect 22026 575 25814 856
rect 25982 575 29862 856
rect 30030 575 33818 856
rect 33986 575 37866 856
rect 38034 575 41822 856
rect 41990 575 45870 856
rect 46038 575 49826 856
rect 49994 575 53874 856
rect 54042 575 57830 856
rect 57998 575 61878 856
rect 62046 575 65834 856
rect 66002 575 69882 856
rect 70050 575 73838 856
rect 74006 575 77886 856
rect 78054 575 81842 856
rect 82010 575 85798 856
rect 85966 575 89846 856
rect 90014 575 93802 856
rect 93970 575 97850 856
rect 98018 575 101806 856
rect 101974 575 105854 856
rect 106022 575 109810 856
rect 109978 575 113858 856
rect 114026 575 117814 856
rect 117982 575 121862 856
rect 122030 575 125818 856
rect 125986 575 129866 856
rect 130034 575 133822 856
rect 133990 575 137870 856
rect 138038 575 141826 856
rect 141994 575 145874 856
rect 146042 575 149830 856
rect 149998 575 153878 856
rect 154046 575 157834 856
rect 158002 575 159508 856
<< metal3 >>
rect 159200 99560 160000 99680
rect 0 98880 800 99000
rect 159200 99016 160000 99136
rect 159200 98608 160000 98728
rect 159200 98064 160000 98184
rect 159200 97656 160000 97776
rect 0 97112 800 97232
rect 159200 97112 160000 97232
rect 159200 96704 160000 96824
rect 159200 96160 160000 96280
rect 159200 95752 160000 95872
rect 0 95344 800 95464
rect 159200 95208 160000 95328
rect 159200 94664 160000 94784
rect 159200 94256 160000 94376
rect 0 93576 800 93696
rect 159200 93712 160000 93832
rect 159200 93304 160000 93424
rect 159200 92760 160000 92880
rect 159200 92352 160000 92472
rect 0 91808 800 91928
rect 159200 91808 160000 91928
rect 159200 91400 160000 91520
rect 159200 90856 160000 90976
rect 159200 90312 160000 90432
rect 0 90040 800 90160
rect 159200 89904 160000 90024
rect 159200 89360 160000 89480
rect 159200 88952 160000 89072
rect 0 88272 800 88392
rect 159200 88408 160000 88528
rect 159200 88000 160000 88120
rect 159200 87456 160000 87576
rect 159200 87048 160000 87168
rect 0 86504 800 86624
rect 159200 86504 160000 86624
rect 159200 86096 160000 86216
rect 159200 85552 160000 85672
rect 159200 85008 160000 85128
rect 0 84600 800 84720
rect 159200 84600 160000 84720
rect 159200 84056 160000 84176
rect 159200 83648 160000 83768
rect 159200 83104 160000 83224
rect 0 82832 800 82952
rect 159200 82696 160000 82816
rect 159200 82152 160000 82272
rect 159200 81744 160000 81864
rect 0 81064 800 81184
rect 159200 81200 160000 81320
rect 159200 80656 160000 80776
rect 159200 80248 160000 80368
rect 159200 79704 160000 79824
rect 0 79296 800 79416
rect 159200 79296 160000 79416
rect 159200 78752 160000 78872
rect 159200 78344 160000 78464
rect 159200 77800 160000 77920
rect 0 77528 800 77648
rect 159200 77392 160000 77512
rect 159200 76848 160000 76968
rect 159200 76440 160000 76560
rect 0 75760 800 75880
rect 159200 75896 160000 76016
rect 159200 75352 160000 75472
rect 159200 74944 160000 75064
rect 159200 74400 160000 74520
rect 0 73992 800 74112
rect 159200 73992 160000 74112
rect 159200 73448 160000 73568
rect 159200 73040 160000 73160
rect 159200 72496 160000 72616
rect 0 72224 800 72344
rect 159200 72088 160000 72208
rect 159200 71544 160000 71664
rect 159200 71000 160000 71120
rect 159200 70592 160000 70712
rect 0 70320 800 70440
rect 159200 70048 160000 70168
rect 159200 69640 160000 69760
rect 159200 69096 160000 69216
rect 0 68552 800 68672
rect 159200 68688 160000 68808
rect 159200 68144 160000 68264
rect 159200 67736 160000 67856
rect 159200 67192 160000 67312
rect 0 66784 800 66904
rect 159200 66784 160000 66904
rect 159200 66240 160000 66360
rect 159200 65696 160000 65816
rect 159200 65288 160000 65408
rect 0 65016 800 65136
rect 159200 64744 160000 64864
rect 159200 64336 160000 64456
rect 159200 63792 160000 63912
rect 0 63248 800 63368
rect 159200 63384 160000 63504
rect 159200 62840 160000 62960
rect 159200 62432 160000 62552
rect 159200 61888 160000 62008
rect 0 61480 800 61600
rect 159200 61344 160000 61464
rect 159200 60936 160000 61056
rect 159200 60392 160000 60512
rect 159200 59984 160000 60104
rect 0 59712 800 59832
rect 159200 59440 160000 59560
rect 159200 59032 160000 59152
rect 159200 58488 160000 58608
rect 0 57944 800 58064
rect 159200 58080 160000 58200
rect 159200 57536 160000 57656
rect 159200 56992 160000 57112
rect 159200 56584 160000 56704
rect 0 56040 800 56160
rect 159200 56040 160000 56160
rect 159200 55632 160000 55752
rect 159200 55088 160000 55208
rect 159200 54680 160000 54800
rect 0 54272 800 54392
rect 159200 54136 160000 54256
rect 159200 53728 160000 53848
rect 159200 53184 160000 53304
rect 159200 52776 160000 52896
rect 0 52504 800 52624
rect 159200 52232 160000 52352
rect 159200 51688 160000 51808
rect 159200 51280 160000 51400
rect 0 50736 800 50856
rect 159200 50736 160000 50856
rect 159200 50328 160000 50448
rect 159200 49784 160000 49904
rect 159200 49376 160000 49496
rect 0 48968 800 49088
rect 159200 48832 160000 48952
rect 159200 48424 160000 48544
rect 159200 47880 160000 48000
rect 0 47200 800 47320
rect 159200 47336 160000 47456
rect 159200 46928 160000 47048
rect 159200 46384 160000 46504
rect 159200 45976 160000 46096
rect 0 45432 800 45552
rect 159200 45432 160000 45552
rect 159200 45024 160000 45144
rect 159200 44480 160000 44600
rect 159200 44072 160000 44192
rect 0 43664 800 43784
rect 159200 43528 160000 43648
rect 159200 43120 160000 43240
rect 159200 42576 160000 42696
rect 159200 42032 160000 42152
rect 0 41760 800 41880
rect 159200 41624 160000 41744
rect 159200 41080 160000 41200
rect 159200 40672 160000 40792
rect 0 39992 800 40112
rect 159200 40128 160000 40248
rect 159200 39720 160000 39840
rect 159200 39176 160000 39296
rect 159200 38768 160000 38888
rect 0 38224 800 38344
rect 159200 38224 160000 38344
rect 159200 37680 160000 37800
rect 159200 37272 160000 37392
rect 159200 36728 160000 36848
rect 0 36456 800 36576
rect 159200 36320 160000 36440
rect 159200 35776 160000 35896
rect 159200 35368 160000 35488
rect 0 34688 800 34808
rect 159200 34824 160000 34944
rect 159200 34416 160000 34536
rect 159200 33872 160000 33992
rect 159200 33464 160000 33584
rect 0 32920 800 33040
rect 159200 32920 160000 33040
rect 159200 32376 160000 32496
rect 159200 31968 160000 32088
rect 159200 31424 160000 31544
rect 0 31152 800 31272
rect 159200 31016 160000 31136
rect 159200 30472 160000 30592
rect 159200 30064 160000 30184
rect 0 29384 800 29504
rect 159200 29520 160000 29640
rect 159200 29112 160000 29232
rect 159200 28568 160000 28688
rect 159200 28024 160000 28144
rect 0 27480 800 27600
rect 159200 27616 160000 27736
rect 159200 27072 160000 27192
rect 159200 26664 160000 26784
rect 159200 26120 160000 26240
rect 0 25712 800 25832
rect 159200 25712 160000 25832
rect 159200 25168 160000 25288
rect 159200 24760 160000 24880
rect 159200 24216 160000 24336
rect 0 23944 800 24064
rect 159200 23672 160000 23792
rect 159200 23264 160000 23384
rect 159200 22720 160000 22840
rect 0 22176 800 22296
rect 159200 22312 160000 22432
rect 159200 21768 160000 21888
rect 159200 21360 160000 21480
rect 159200 20816 160000 20936
rect 0 20408 800 20528
rect 159200 20408 160000 20528
rect 159200 19864 160000 19984
rect 159200 19456 160000 19576
rect 159200 18912 160000 19032
rect 0 18640 800 18760
rect 159200 18368 160000 18488
rect 159200 17960 160000 18080
rect 159200 17416 160000 17536
rect 0 16872 800 16992
rect 159200 17008 160000 17128
rect 159200 16464 160000 16584
rect 159200 16056 160000 16176
rect 159200 15512 160000 15632
rect 0 15104 800 15224
rect 159200 15104 160000 15224
rect 159200 14560 160000 14680
rect 159200 14016 160000 14136
rect 159200 13608 160000 13728
rect 0 13200 800 13320
rect 159200 13064 160000 13184
rect 159200 12656 160000 12776
rect 159200 12112 160000 12232
rect 159200 11704 160000 11824
rect 0 11432 800 11552
rect 159200 11160 160000 11280
rect 159200 10752 160000 10872
rect 159200 10208 160000 10328
rect 0 9664 800 9784
rect 159200 9800 160000 9920
rect 159200 9256 160000 9376
rect 159200 8712 160000 8832
rect 159200 8304 160000 8424
rect 0 7896 800 8016
rect 159200 7760 160000 7880
rect 159200 7352 160000 7472
rect 159200 6808 160000 6928
rect 159200 6400 160000 6520
rect 0 6128 800 6248
rect 159200 5856 160000 5976
rect 159200 5448 160000 5568
rect 159200 4904 160000 5024
rect 0 4360 800 4480
rect 159200 4360 160000 4480
rect 159200 3952 160000 4072
rect 159200 3408 160000 3528
rect 159200 3000 160000 3120
rect 0 2592 800 2712
rect 159200 2456 160000 2576
rect 159200 2048 160000 2168
rect 159200 1504 160000 1624
rect 159200 1096 160000 1216
rect 0 824 800 944
rect 159200 552 160000 672
rect 159200 144 160000 264
<< obsm3 >>
rect 800 99480 159120 99653
rect 800 99216 159200 99480
rect 800 99080 159120 99216
rect 880 98936 159120 99080
rect 880 98808 159200 98936
rect 880 98800 159120 98808
rect 800 98528 159120 98800
rect 800 98264 159200 98528
rect 800 97984 159120 98264
rect 800 97856 159200 97984
rect 800 97576 159120 97856
rect 800 97312 159200 97576
rect 880 97032 159120 97312
rect 800 96904 159200 97032
rect 800 96624 159120 96904
rect 800 96360 159200 96624
rect 800 96080 159120 96360
rect 800 95952 159200 96080
rect 800 95672 159120 95952
rect 800 95544 159200 95672
rect 880 95408 159200 95544
rect 880 95264 159120 95408
rect 800 95128 159120 95264
rect 800 94864 159200 95128
rect 800 94584 159120 94864
rect 800 94456 159200 94584
rect 800 94176 159120 94456
rect 800 93912 159200 94176
rect 800 93776 159120 93912
rect 880 93632 159120 93776
rect 880 93504 159200 93632
rect 880 93496 159120 93504
rect 800 93224 159120 93496
rect 800 92960 159200 93224
rect 800 92680 159120 92960
rect 800 92552 159200 92680
rect 800 92272 159120 92552
rect 800 92008 159200 92272
rect 880 91728 159120 92008
rect 800 91600 159200 91728
rect 800 91320 159120 91600
rect 800 91056 159200 91320
rect 800 90776 159120 91056
rect 800 90512 159200 90776
rect 800 90240 159120 90512
rect 880 90232 159120 90240
rect 880 90104 159200 90232
rect 880 89960 159120 90104
rect 800 89824 159120 89960
rect 800 89560 159200 89824
rect 800 89280 159120 89560
rect 800 89152 159200 89280
rect 800 88872 159120 89152
rect 800 88608 159200 88872
rect 800 88472 159120 88608
rect 880 88328 159120 88472
rect 880 88200 159200 88328
rect 880 88192 159120 88200
rect 800 87920 159120 88192
rect 800 87656 159200 87920
rect 800 87376 159120 87656
rect 800 87248 159200 87376
rect 800 86968 159120 87248
rect 800 86704 159200 86968
rect 880 86424 159120 86704
rect 800 86296 159200 86424
rect 800 86016 159120 86296
rect 800 85752 159200 86016
rect 800 85472 159120 85752
rect 800 85208 159200 85472
rect 800 84928 159120 85208
rect 800 84800 159200 84928
rect 880 84520 159120 84800
rect 800 84256 159200 84520
rect 800 83976 159120 84256
rect 800 83848 159200 83976
rect 800 83568 159120 83848
rect 800 83304 159200 83568
rect 800 83032 159120 83304
rect 880 83024 159120 83032
rect 880 82896 159200 83024
rect 880 82752 159120 82896
rect 800 82616 159120 82752
rect 800 82352 159200 82616
rect 800 82072 159120 82352
rect 800 81944 159200 82072
rect 800 81664 159120 81944
rect 800 81400 159200 81664
rect 800 81264 159120 81400
rect 880 81120 159120 81264
rect 880 80984 159200 81120
rect 800 80856 159200 80984
rect 800 80576 159120 80856
rect 800 80448 159200 80576
rect 800 80168 159120 80448
rect 800 79904 159200 80168
rect 800 79624 159120 79904
rect 800 79496 159200 79624
rect 880 79216 159120 79496
rect 800 78952 159200 79216
rect 800 78672 159120 78952
rect 800 78544 159200 78672
rect 800 78264 159120 78544
rect 800 78000 159200 78264
rect 800 77728 159120 78000
rect 880 77720 159120 77728
rect 880 77592 159200 77720
rect 880 77448 159120 77592
rect 800 77312 159120 77448
rect 800 77048 159200 77312
rect 800 76768 159120 77048
rect 800 76640 159200 76768
rect 800 76360 159120 76640
rect 800 76096 159200 76360
rect 800 75960 159120 76096
rect 880 75816 159120 75960
rect 880 75680 159200 75816
rect 800 75552 159200 75680
rect 800 75272 159120 75552
rect 800 75144 159200 75272
rect 800 74864 159120 75144
rect 800 74600 159200 74864
rect 800 74320 159120 74600
rect 800 74192 159200 74320
rect 880 73912 159120 74192
rect 800 73648 159200 73912
rect 800 73368 159120 73648
rect 800 73240 159200 73368
rect 800 72960 159120 73240
rect 800 72696 159200 72960
rect 800 72424 159120 72696
rect 880 72416 159120 72424
rect 880 72288 159200 72416
rect 880 72144 159120 72288
rect 800 72008 159120 72144
rect 800 71744 159200 72008
rect 800 71464 159120 71744
rect 800 71200 159200 71464
rect 800 70920 159120 71200
rect 800 70792 159200 70920
rect 800 70520 159120 70792
rect 880 70512 159120 70520
rect 880 70248 159200 70512
rect 880 70240 159120 70248
rect 800 69968 159120 70240
rect 800 69840 159200 69968
rect 800 69560 159120 69840
rect 800 69296 159200 69560
rect 800 69016 159120 69296
rect 800 68888 159200 69016
rect 800 68752 159120 68888
rect 880 68608 159120 68752
rect 880 68472 159200 68608
rect 800 68344 159200 68472
rect 800 68064 159120 68344
rect 800 67936 159200 68064
rect 800 67656 159120 67936
rect 800 67392 159200 67656
rect 800 67112 159120 67392
rect 800 66984 159200 67112
rect 880 66704 159120 66984
rect 800 66440 159200 66704
rect 800 66160 159120 66440
rect 800 65896 159200 66160
rect 800 65616 159120 65896
rect 800 65488 159200 65616
rect 800 65216 159120 65488
rect 880 65208 159120 65216
rect 880 64944 159200 65208
rect 880 64936 159120 64944
rect 800 64664 159120 64936
rect 800 64536 159200 64664
rect 800 64256 159120 64536
rect 800 63992 159200 64256
rect 800 63712 159120 63992
rect 800 63584 159200 63712
rect 800 63448 159120 63584
rect 880 63304 159120 63448
rect 880 63168 159200 63304
rect 800 63040 159200 63168
rect 800 62760 159120 63040
rect 800 62632 159200 62760
rect 800 62352 159120 62632
rect 800 62088 159200 62352
rect 800 61808 159120 62088
rect 800 61680 159200 61808
rect 880 61544 159200 61680
rect 880 61400 159120 61544
rect 800 61264 159120 61400
rect 800 61136 159200 61264
rect 800 60856 159120 61136
rect 800 60592 159200 60856
rect 800 60312 159120 60592
rect 800 60184 159200 60312
rect 800 59912 159120 60184
rect 880 59904 159120 59912
rect 880 59640 159200 59904
rect 880 59632 159120 59640
rect 800 59360 159120 59632
rect 800 59232 159200 59360
rect 800 58952 159120 59232
rect 800 58688 159200 58952
rect 800 58408 159120 58688
rect 800 58280 159200 58408
rect 800 58144 159120 58280
rect 880 58000 159120 58144
rect 880 57864 159200 58000
rect 800 57736 159200 57864
rect 800 57456 159120 57736
rect 800 57192 159200 57456
rect 800 56912 159120 57192
rect 800 56784 159200 56912
rect 800 56504 159120 56784
rect 800 56240 159200 56504
rect 880 55960 159120 56240
rect 800 55832 159200 55960
rect 800 55552 159120 55832
rect 800 55288 159200 55552
rect 800 55008 159120 55288
rect 800 54880 159200 55008
rect 800 54600 159120 54880
rect 800 54472 159200 54600
rect 880 54336 159200 54472
rect 880 54192 159120 54336
rect 800 54056 159120 54192
rect 800 53928 159200 54056
rect 800 53648 159120 53928
rect 800 53384 159200 53648
rect 800 53104 159120 53384
rect 800 52976 159200 53104
rect 800 52704 159120 52976
rect 880 52696 159120 52704
rect 880 52432 159200 52696
rect 880 52424 159120 52432
rect 800 52152 159120 52424
rect 800 51888 159200 52152
rect 800 51608 159120 51888
rect 800 51480 159200 51608
rect 800 51200 159120 51480
rect 800 50936 159200 51200
rect 880 50656 159120 50936
rect 800 50528 159200 50656
rect 800 50248 159120 50528
rect 800 49984 159200 50248
rect 800 49704 159120 49984
rect 800 49576 159200 49704
rect 800 49296 159120 49576
rect 800 49168 159200 49296
rect 880 49032 159200 49168
rect 880 48888 159120 49032
rect 800 48752 159120 48888
rect 800 48624 159200 48752
rect 800 48344 159120 48624
rect 800 48080 159200 48344
rect 800 47800 159120 48080
rect 800 47536 159200 47800
rect 800 47400 159120 47536
rect 880 47256 159120 47400
rect 880 47128 159200 47256
rect 880 47120 159120 47128
rect 800 46848 159120 47120
rect 800 46584 159200 46848
rect 800 46304 159120 46584
rect 800 46176 159200 46304
rect 800 45896 159120 46176
rect 800 45632 159200 45896
rect 880 45352 159120 45632
rect 800 45224 159200 45352
rect 800 44944 159120 45224
rect 800 44680 159200 44944
rect 800 44400 159120 44680
rect 800 44272 159200 44400
rect 800 43992 159120 44272
rect 800 43864 159200 43992
rect 880 43728 159200 43864
rect 880 43584 159120 43728
rect 800 43448 159120 43584
rect 800 43320 159200 43448
rect 800 43040 159120 43320
rect 800 42776 159200 43040
rect 800 42496 159120 42776
rect 800 42232 159200 42496
rect 800 41960 159120 42232
rect 880 41952 159120 41960
rect 880 41824 159200 41952
rect 880 41680 159120 41824
rect 800 41544 159120 41680
rect 800 41280 159200 41544
rect 800 41000 159120 41280
rect 800 40872 159200 41000
rect 800 40592 159120 40872
rect 800 40328 159200 40592
rect 800 40192 159120 40328
rect 880 40048 159120 40192
rect 880 39920 159200 40048
rect 880 39912 159120 39920
rect 800 39640 159120 39912
rect 800 39376 159200 39640
rect 800 39096 159120 39376
rect 800 38968 159200 39096
rect 800 38688 159120 38968
rect 800 38424 159200 38688
rect 880 38144 159120 38424
rect 800 37880 159200 38144
rect 800 37600 159120 37880
rect 800 37472 159200 37600
rect 800 37192 159120 37472
rect 800 36928 159200 37192
rect 800 36656 159120 36928
rect 880 36648 159120 36656
rect 880 36520 159200 36648
rect 880 36376 159120 36520
rect 800 36240 159120 36376
rect 800 35976 159200 36240
rect 800 35696 159120 35976
rect 800 35568 159200 35696
rect 800 35288 159120 35568
rect 800 35024 159200 35288
rect 800 34888 159120 35024
rect 880 34744 159120 34888
rect 880 34616 159200 34744
rect 880 34608 159120 34616
rect 800 34336 159120 34608
rect 800 34072 159200 34336
rect 800 33792 159120 34072
rect 800 33664 159200 33792
rect 800 33384 159120 33664
rect 800 33120 159200 33384
rect 880 32840 159120 33120
rect 800 32576 159200 32840
rect 800 32296 159120 32576
rect 800 32168 159200 32296
rect 800 31888 159120 32168
rect 800 31624 159200 31888
rect 800 31352 159120 31624
rect 880 31344 159120 31352
rect 880 31216 159200 31344
rect 880 31072 159120 31216
rect 800 30936 159120 31072
rect 800 30672 159200 30936
rect 800 30392 159120 30672
rect 800 30264 159200 30392
rect 800 29984 159120 30264
rect 800 29720 159200 29984
rect 800 29584 159120 29720
rect 880 29440 159120 29584
rect 880 29312 159200 29440
rect 880 29304 159120 29312
rect 800 29032 159120 29304
rect 800 28768 159200 29032
rect 800 28488 159120 28768
rect 800 28224 159200 28488
rect 800 27944 159120 28224
rect 800 27816 159200 27944
rect 800 27680 159120 27816
rect 880 27536 159120 27680
rect 880 27400 159200 27536
rect 800 27272 159200 27400
rect 800 26992 159120 27272
rect 800 26864 159200 26992
rect 800 26584 159120 26864
rect 800 26320 159200 26584
rect 800 26040 159120 26320
rect 800 25912 159200 26040
rect 880 25632 159120 25912
rect 800 25368 159200 25632
rect 800 25088 159120 25368
rect 800 24960 159200 25088
rect 800 24680 159120 24960
rect 800 24416 159200 24680
rect 800 24144 159120 24416
rect 880 24136 159120 24144
rect 880 23872 159200 24136
rect 880 23864 159120 23872
rect 800 23592 159120 23864
rect 800 23464 159200 23592
rect 800 23184 159120 23464
rect 800 22920 159200 23184
rect 800 22640 159120 22920
rect 800 22512 159200 22640
rect 800 22376 159120 22512
rect 880 22232 159120 22376
rect 880 22096 159200 22232
rect 800 21968 159200 22096
rect 800 21688 159120 21968
rect 800 21560 159200 21688
rect 800 21280 159120 21560
rect 800 21016 159200 21280
rect 800 20736 159120 21016
rect 800 20608 159200 20736
rect 880 20328 159120 20608
rect 800 20064 159200 20328
rect 800 19784 159120 20064
rect 800 19656 159200 19784
rect 800 19376 159120 19656
rect 800 19112 159200 19376
rect 800 18840 159120 19112
rect 880 18832 159120 18840
rect 880 18568 159200 18832
rect 880 18560 159120 18568
rect 800 18288 159120 18560
rect 800 18160 159200 18288
rect 800 17880 159120 18160
rect 800 17616 159200 17880
rect 800 17336 159120 17616
rect 800 17208 159200 17336
rect 800 17072 159120 17208
rect 880 16928 159120 17072
rect 880 16792 159200 16928
rect 800 16664 159200 16792
rect 800 16384 159120 16664
rect 800 16256 159200 16384
rect 800 15976 159120 16256
rect 800 15712 159200 15976
rect 800 15432 159120 15712
rect 800 15304 159200 15432
rect 880 15024 159120 15304
rect 800 14760 159200 15024
rect 800 14480 159120 14760
rect 800 14216 159200 14480
rect 800 13936 159120 14216
rect 800 13808 159200 13936
rect 800 13528 159120 13808
rect 800 13400 159200 13528
rect 880 13264 159200 13400
rect 880 13120 159120 13264
rect 800 12984 159120 13120
rect 800 12856 159200 12984
rect 800 12576 159120 12856
rect 800 12312 159200 12576
rect 800 12032 159120 12312
rect 800 11904 159200 12032
rect 800 11632 159120 11904
rect 880 11624 159120 11632
rect 880 11360 159200 11624
rect 880 11352 159120 11360
rect 800 11080 159120 11352
rect 800 10952 159200 11080
rect 800 10672 159120 10952
rect 800 10408 159200 10672
rect 800 10128 159120 10408
rect 800 10000 159200 10128
rect 800 9864 159120 10000
rect 880 9720 159120 9864
rect 880 9584 159200 9720
rect 800 9456 159200 9584
rect 800 9176 159120 9456
rect 800 8912 159200 9176
rect 800 8632 159120 8912
rect 800 8504 159200 8632
rect 800 8224 159120 8504
rect 800 8096 159200 8224
rect 880 7960 159200 8096
rect 880 7816 159120 7960
rect 800 7680 159120 7816
rect 800 7552 159200 7680
rect 800 7272 159120 7552
rect 800 7008 159200 7272
rect 800 6728 159120 7008
rect 800 6600 159200 6728
rect 800 6328 159120 6600
rect 880 6320 159120 6328
rect 880 6056 159200 6320
rect 880 6048 159120 6056
rect 800 5776 159120 6048
rect 800 5648 159200 5776
rect 800 5368 159120 5648
rect 800 5104 159200 5368
rect 800 4824 159120 5104
rect 800 4560 159200 4824
rect 880 4280 159120 4560
rect 800 4152 159200 4280
rect 800 3872 159120 4152
rect 800 3608 159200 3872
rect 800 3328 159120 3608
rect 800 3200 159200 3328
rect 800 2920 159120 3200
rect 800 2792 159200 2920
rect 880 2656 159200 2792
rect 880 2512 159120 2656
rect 800 2376 159120 2512
rect 800 2248 159200 2376
rect 800 1968 159120 2248
rect 800 1704 159200 1968
rect 800 1424 159120 1704
rect 800 1296 159200 1424
rect 800 1024 159120 1296
rect 880 1016 159120 1024
rect 880 752 159200 1016
rect 880 744 159120 752
rect 800 472 159120 744
rect 800 344 159200 472
rect 800 64 159120 344
rect 800 36 159200 64
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
rect 111728 2128 112048 97424
rect 127088 2128 127408 97424
rect 142448 2128 142768 97424
rect 157808 2128 158128 97424
<< obsm4 >>
rect 22323 97504 157261 97885
rect 22323 2048 34848 97504
rect 35328 2048 50208 97504
rect 50688 2048 65568 97504
rect 66048 2048 80928 97504
rect 81408 2048 96288 97504
rect 96768 2048 111648 97504
rect 112128 2048 127008 97504
rect 127488 2048 142368 97504
rect 142848 2048 157261 97504
rect 22323 35 157261 2048
<< labels >>
rlabel metal2 s 5538 99200 5594 100000 6 addr0[0]
port 1 nsew signal output
rlabel metal2 s 6366 99200 6422 100000 6 addr0[1]
port 2 nsew signal output
rlabel metal2 s 7194 99200 7250 100000 6 addr0[2]
port 3 nsew signal output
rlabel metal2 s 8114 99200 8170 100000 6 addr0[3]
port 4 nsew signal output
rlabel metal2 s 8942 99200 8998 100000 6 addr0[4]
port 5 nsew signal output
rlabel metal2 s 9770 99200 9826 100000 6 addr0[5]
port 6 nsew signal output
rlabel metal2 s 10690 99200 10746 100000 6 addr0[6]
port 7 nsew signal output
rlabel metal2 s 11518 99200 11574 100000 6 addr0[7]
port 8 nsew signal output
rlabel metal2 s 12346 99200 12402 100000 6 addr0[8]
port 9 nsew signal output
rlabel metal2 s 96710 99200 96766 100000 6 addr1[0]
port 10 nsew signal output
rlabel metal2 s 97538 99200 97594 100000 6 addr1[1]
port 11 nsew signal output
rlabel metal2 s 98366 99200 98422 100000 6 addr1[2]
port 12 nsew signal output
rlabel metal2 s 99286 99200 99342 100000 6 addr1[3]
port 13 nsew signal output
rlabel metal2 s 100114 99200 100170 100000 6 addr1[4]
port 14 nsew signal output
rlabel metal2 s 100942 99200 100998 100000 6 addr1[5]
port 15 nsew signal output
rlabel metal2 s 101862 99200 101918 100000 6 addr1[6]
port 16 nsew signal output
rlabel metal2 s 102690 99200 102746 100000 6 addr1[7]
port 17 nsew signal output
rlabel metal2 s 103518 99200 103574 100000 6 addr1[8]
port 18 nsew signal output
rlabel metal2 s 386 99200 442 100000 6 clk0
port 19 nsew signal output
rlabel metal2 s 95790 99200 95846 100000 6 clk1
port 20 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 coreIndex[0]
port 21 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 coreIndex[1]
port 22 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 coreIndex[2]
port 23 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 coreIndex[3]
port 24 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 coreIndex[4]
port 25 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 coreIndex[5]
port 26 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 coreIndex[6]
port 27 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 coreIndex[7]
port 28 nsew signal input
rlabel metal3 s 159200 1096 160000 1216 6 core_wb_ack_i
port 29 nsew signal input
rlabel metal3 s 159200 3952 160000 4072 6 core_wb_adr_o[0]
port 30 nsew signal output
rlabel metal3 s 159200 20408 160000 20528 6 core_wb_adr_o[10]
port 31 nsew signal output
rlabel metal3 s 159200 21768 160000 21888 6 core_wb_adr_o[11]
port 32 nsew signal output
rlabel metal3 s 159200 23264 160000 23384 6 core_wb_adr_o[12]
port 33 nsew signal output
rlabel metal3 s 159200 24760 160000 24880 6 core_wb_adr_o[13]
port 34 nsew signal output
rlabel metal3 s 159200 26120 160000 26240 6 core_wb_adr_o[14]
port 35 nsew signal output
rlabel metal3 s 159200 27616 160000 27736 6 core_wb_adr_o[15]
port 36 nsew signal output
rlabel metal3 s 159200 29112 160000 29232 6 core_wb_adr_o[16]
port 37 nsew signal output
rlabel metal3 s 159200 30472 160000 30592 6 core_wb_adr_o[17]
port 38 nsew signal output
rlabel metal3 s 159200 31968 160000 32088 6 core_wb_adr_o[18]
port 39 nsew signal output
rlabel metal3 s 159200 33464 160000 33584 6 core_wb_adr_o[19]
port 40 nsew signal output
rlabel metal3 s 159200 5856 160000 5976 6 core_wb_adr_o[1]
port 41 nsew signal output
rlabel metal3 s 159200 34824 160000 34944 6 core_wb_adr_o[20]
port 42 nsew signal output
rlabel metal3 s 159200 36320 160000 36440 6 core_wb_adr_o[21]
port 43 nsew signal output
rlabel metal3 s 159200 37680 160000 37800 6 core_wb_adr_o[22]
port 44 nsew signal output
rlabel metal3 s 159200 39176 160000 39296 6 core_wb_adr_o[23]
port 45 nsew signal output
rlabel metal3 s 159200 40672 160000 40792 6 core_wb_adr_o[24]
port 46 nsew signal output
rlabel metal3 s 159200 42032 160000 42152 6 core_wb_adr_o[25]
port 47 nsew signal output
rlabel metal3 s 159200 43528 160000 43648 6 core_wb_adr_o[26]
port 48 nsew signal output
rlabel metal3 s 159200 45024 160000 45144 6 core_wb_adr_o[27]
port 49 nsew signal output
rlabel metal3 s 159200 7760 160000 7880 6 core_wb_adr_o[2]
port 50 nsew signal output
rlabel metal3 s 159200 9800 160000 9920 6 core_wb_adr_o[3]
port 51 nsew signal output
rlabel metal3 s 159200 11704 160000 11824 6 core_wb_adr_o[4]
port 52 nsew signal output
rlabel metal3 s 159200 13064 160000 13184 6 core_wb_adr_o[5]
port 53 nsew signal output
rlabel metal3 s 159200 14560 160000 14680 6 core_wb_adr_o[6]
port 54 nsew signal output
rlabel metal3 s 159200 16056 160000 16176 6 core_wb_adr_o[7]
port 55 nsew signal output
rlabel metal3 s 159200 17416 160000 17536 6 core_wb_adr_o[8]
port 56 nsew signal output
rlabel metal3 s 159200 18912 160000 19032 6 core_wb_adr_o[9]
port 57 nsew signal output
rlabel metal3 s 159200 1504 160000 1624 6 core_wb_cyc_o
port 58 nsew signal output
rlabel metal3 s 159200 4360 160000 4480 6 core_wb_data_i[0]
port 59 nsew signal input
rlabel metal3 s 159200 20816 160000 20936 6 core_wb_data_i[10]
port 60 nsew signal input
rlabel metal3 s 159200 22312 160000 22432 6 core_wb_data_i[11]
port 61 nsew signal input
rlabel metal3 s 159200 23672 160000 23792 6 core_wb_data_i[12]
port 62 nsew signal input
rlabel metal3 s 159200 25168 160000 25288 6 core_wb_data_i[13]
port 63 nsew signal input
rlabel metal3 s 159200 26664 160000 26784 6 core_wb_data_i[14]
port 64 nsew signal input
rlabel metal3 s 159200 28024 160000 28144 6 core_wb_data_i[15]
port 65 nsew signal input
rlabel metal3 s 159200 29520 160000 29640 6 core_wb_data_i[16]
port 66 nsew signal input
rlabel metal3 s 159200 31016 160000 31136 6 core_wb_data_i[17]
port 67 nsew signal input
rlabel metal3 s 159200 32376 160000 32496 6 core_wb_data_i[18]
port 68 nsew signal input
rlabel metal3 s 159200 33872 160000 33992 6 core_wb_data_i[19]
port 69 nsew signal input
rlabel metal3 s 159200 6400 160000 6520 6 core_wb_data_i[1]
port 70 nsew signal input
rlabel metal3 s 159200 35368 160000 35488 6 core_wb_data_i[20]
port 71 nsew signal input
rlabel metal3 s 159200 36728 160000 36848 6 core_wb_data_i[21]
port 72 nsew signal input
rlabel metal3 s 159200 38224 160000 38344 6 core_wb_data_i[22]
port 73 nsew signal input
rlabel metal3 s 159200 39720 160000 39840 6 core_wb_data_i[23]
port 74 nsew signal input
rlabel metal3 s 159200 41080 160000 41200 6 core_wb_data_i[24]
port 75 nsew signal input
rlabel metal3 s 159200 42576 160000 42696 6 core_wb_data_i[25]
port 76 nsew signal input
rlabel metal3 s 159200 44072 160000 44192 6 core_wb_data_i[26]
port 77 nsew signal input
rlabel metal3 s 159200 45432 160000 45552 6 core_wb_data_i[27]
port 78 nsew signal input
rlabel metal3 s 159200 46384 160000 46504 6 core_wb_data_i[28]
port 79 nsew signal input
rlabel metal3 s 159200 47336 160000 47456 6 core_wb_data_i[29]
port 80 nsew signal input
rlabel metal3 s 159200 8304 160000 8424 6 core_wb_data_i[2]
port 81 nsew signal input
rlabel metal3 s 159200 48424 160000 48544 6 core_wb_data_i[30]
port 82 nsew signal input
rlabel metal3 s 159200 49376 160000 49496 6 core_wb_data_i[31]
port 83 nsew signal input
rlabel metal3 s 159200 10208 160000 10328 6 core_wb_data_i[3]
port 84 nsew signal input
rlabel metal3 s 159200 12112 160000 12232 6 core_wb_data_i[4]
port 85 nsew signal input
rlabel metal3 s 159200 13608 160000 13728 6 core_wb_data_i[5]
port 86 nsew signal input
rlabel metal3 s 159200 15104 160000 15224 6 core_wb_data_i[6]
port 87 nsew signal input
rlabel metal3 s 159200 16464 160000 16584 6 core_wb_data_i[7]
port 88 nsew signal input
rlabel metal3 s 159200 17960 160000 18080 6 core_wb_data_i[8]
port 89 nsew signal input
rlabel metal3 s 159200 19456 160000 19576 6 core_wb_data_i[9]
port 90 nsew signal input
rlabel metal3 s 159200 4904 160000 5024 6 core_wb_data_o[0]
port 91 nsew signal output
rlabel metal3 s 159200 21360 160000 21480 6 core_wb_data_o[10]
port 92 nsew signal output
rlabel metal3 s 159200 22720 160000 22840 6 core_wb_data_o[11]
port 93 nsew signal output
rlabel metal3 s 159200 24216 160000 24336 6 core_wb_data_o[12]
port 94 nsew signal output
rlabel metal3 s 159200 25712 160000 25832 6 core_wb_data_o[13]
port 95 nsew signal output
rlabel metal3 s 159200 27072 160000 27192 6 core_wb_data_o[14]
port 96 nsew signal output
rlabel metal3 s 159200 28568 160000 28688 6 core_wb_data_o[15]
port 97 nsew signal output
rlabel metal3 s 159200 30064 160000 30184 6 core_wb_data_o[16]
port 98 nsew signal output
rlabel metal3 s 159200 31424 160000 31544 6 core_wb_data_o[17]
port 99 nsew signal output
rlabel metal3 s 159200 32920 160000 33040 6 core_wb_data_o[18]
port 100 nsew signal output
rlabel metal3 s 159200 34416 160000 34536 6 core_wb_data_o[19]
port 101 nsew signal output
rlabel metal3 s 159200 6808 160000 6928 6 core_wb_data_o[1]
port 102 nsew signal output
rlabel metal3 s 159200 35776 160000 35896 6 core_wb_data_o[20]
port 103 nsew signal output
rlabel metal3 s 159200 37272 160000 37392 6 core_wb_data_o[21]
port 104 nsew signal output
rlabel metal3 s 159200 38768 160000 38888 6 core_wb_data_o[22]
port 105 nsew signal output
rlabel metal3 s 159200 40128 160000 40248 6 core_wb_data_o[23]
port 106 nsew signal output
rlabel metal3 s 159200 41624 160000 41744 6 core_wb_data_o[24]
port 107 nsew signal output
rlabel metal3 s 159200 43120 160000 43240 6 core_wb_data_o[25]
port 108 nsew signal output
rlabel metal3 s 159200 44480 160000 44600 6 core_wb_data_o[26]
port 109 nsew signal output
rlabel metal3 s 159200 45976 160000 46096 6 core_wb_data_o[27]
port 110 nsew signal output
rlabel metal3 s 159200 46928 160000 47048 6 core_wb_data_o[28]
port 111 nsew signal output
rlabel metal3 s 159200 47880 160000 48000 6 core_wb_data_o[29]
port 112 nsew signal output
rlabel metal3 s 159200 8712 160000 8832 6 core_wb_data_o[2]
port 113 nsew signal output
rlabel metal3 s 159200 48832 160000 48952 6 core_wb_data_o[30]
port 114 nsew signal output
rlabel metal3 s 159200 49784 160000 49904 6 core_wb_data_o[31]
port 115 nsew signal output
rlabel metal3 s 159200 10752 160000 10872 6 core_wb_data_o[3]
port 116 nsew signal output
rlabel metal3 s 159200 12656 160000 12776 6 core_wb_data_o[4]
port 117 nsew signal output
rlabel metal3 s 159200 14016 160000 14136 6 core_wb_data_o[5]
port 118 nsew signal output
rlabel metal3 s 159200 15512 160000 15632 6 core_wb_data_o[6]
port 119 nsew signal output
rlabel metal3 s 159200 17008 160000 17128 6 core_wb_data_o[7]
port 120 nsew signal output
rlabel metal3 s 159200 18368 160000 18488 6 core_wb_data_o[8]
port 121 nsew signal output
rlabel metal3 s 159200 19864 160000 19984 6 core_wb_data_o[9]
port 122 nsew signal output
rlabel metal3 s 159200 2048 160000 2168 6 core_wb_error_i
port 123 nsew signal input
rlabel metal3 s 159200 5448 160000 5568 6 core_wb_sel_o[0]
port 124 nsew signal output
rlabel metal3 s 159200 7352 160000 7472 6 core_wb_sel_o[1]
port 125 nsew signal output
rlabel metal3 s 159200 9256 160000 9376 6 core_wb_sel_o[2]
port 126 nsew signal output
rlabel metal3 s 159200 11160 160000 11280 6 core_wb_sel_o[3]
port 127 nsew signal output
rlabel metal3 s 159200 2456 160000 2576 6 core_wb_stall_i
port 128 nsew signal input
rlabel metal3 s 159200 3000 160000 3120 6 core_wb_stb_o
port 129 nsew signal output
rlabel metal3 s 159200 3408 160000 3528 6 core_wb_we_o
port 130 nsew signal output
rlabel metal3 s 159200 98608 160000 98728 6 csb0[0]
port 131 nsew signal output
rlabel metal3 s 159200 99016 160000 99136 6 csb0[1]
port 132 nsew signal output
rlabel metal3 s 0 98880 800 99000 6 csb1[0]
port 133 nsew signal output
rlabel metal3 s 159200 99560 160000 99680 6 csb1[1]
port 134 nsew signal output
rlabel metal2 s 13266 99200 13322 100000 6 din0[0]
port 135 nsew signal output
rlabel metal2 s 21822 99200 21878 100000 6 din0[10]
port 136 nsew signal output
rlabel metal2 s 22742 99200 22798 100000 6 din0[11]
port 137 nsew signal output
rlabel metal2 s 23570 99200 23626 100000 6 din0[12]
port 138 nsew signal output
rlabel metal2 s 24398 99200 24454 100000 6 din0[13]
port 139 nsew signal output
rlabel metal2 s 25318 99200 25374 100000 6 din0[14]
port 140 nsew signal output
rlabel metal2 s 26146 99200 26202 100000 6 din0[15]
port 141 nsew signal output
rlabel metal2 s 26974 99200 27030 100000 6 din0[16]
port 142 nsew signal output
rlabel metal2 s 27894 99200 27950 100000 6 din0[17]
port 143 nsew signal output
rlabel metal2 s 28722 99200 28778 100000 6 din0[18]
port 144 nsew signal output
rlabel metal2 s 29550 99200 29606 100000 6 din0[19]
port 145 nsew signal output
rlabel metal2 s 14094 99200 14150 100000 6 din0[1]
port 146 nsew signal output
rlabel metal2 s 30470 99200 30526 100000 6 din0[20]
port 147 nsew signal output
rlabel metal2 s 31298 99200 31354 100000 6 din0[21]
port 148 nsew signal output
rlabel metal2 s 32126 99200 32182 100000 6 din0[22]
port 149 nsew signal output
rlabel metal2 s 33046 99200 33102 100000 6 din0[23]
port 150 nsew signal output
rlabel metal2 s 33874 99200 33930 100000 6 din0[24]
port 151 nsew signal output
rlabel metal2 s 34702 99200 34758 100000 6 din0[25]
port 152 nsew signal output
rlabel metal2 s 35622 99200 35678 100000 6 din0[26]
port 153 nsew signal output
rlabel metal2 s 36450 99200 36506 100000 6 din0[27]
port 154 nsew signal output
rlabel metal2 s 37370 99200 37426 100000 6 din0[28]
port 155 nsew signal output
rlabel metal2 s 38198 99200 38254 100000 6 din0[29]
port 156 nsew signal output
rlabel metal2 s 14922 99200 14978 100000 6 din0[2]
port 157 nsew signal output
rlabel metal2 s 39026 99200 39082 100000 6 din0[30]
port 158 nsew signal output
rlabel metal2 s 39946 99200 40002 100000 6 din0[31]
port 159 nsew signal output
rlabel metal2 s 15842 99200 15898 100000 6 din0[3]
port 160 nsew signal output
rlabel metal2 s 16670 99200 16726 100000 6 din0[4]
port 161 nsew signal output
rlabel metal2 s 17498 99200 17554 100000 6 din0[5]
port 162 nsew signal output
rlabel metal2 s 18418 99200 18474 100000 6 din0[6]
port 163 nsew signal output
rlabel metal2 s 19246 99200 19302 100000 6 din0[7]
port 164 nsew signal output
rlabel metal2 s 20166 99200 20222 100000 6 din0[8]
port 165 nsew signal output
rlabel metal2 s 20994 99200 21050 100000 6 din0[9]
port 166 nsew signal output
rlabel metal2 s 40774 99200 40830 100000 6 dout0[0]
port 167 nsew signal input
rlabel metal2 s 49330 99200 49386 100000 6 dout0[10]
port 168 nsew signal input
rlabel metal2 s 50250 99200 50306 100000 6 dout0[11]
port 169 nsew signal input
rlabel metal2 s 51078 99200 51134 100000 6 dout0[12]
port 170 nsew signal input
rlabel metal2 s 51906 99200 51962 100000 6 dout0[13]
port 171 nsew signal input
rlabel metal2 s 52826 99200 52882 100000 6 dout0[14]
port 172 nsew signal input
rlabel metal2 s 53654 99200 53710 100000 6 dout0[15]
port 173 nsew signal input
rlabel metal2 s 54574 99200 54630 100000 6 dout0[16]
port 174 nsew signal input
rlabel metal2 s 55402 99200 55458 100000 6 dout0[17]
port 175 nsew signal input
rlabel metal2 s 56230 99200 56286 100000 6 dout0[18]
port 176 nsew signal input
rlabel metal2 s 57150 99200 57206 100000 6 dout0[19]
port 177 nsew signal input
rlabel metal2 s 41602 99200 41658 100000 6 dout0[1]
port 178 nsew signal input
rlabel metal2 s 57978 99200 58034 100000 6 dout0[20]
port 179 nsew signal input
rlabel metal2 s 58806 99200 58862 100000 6 dout0[21]
port 180 nsew signal input
rlabel metal2 s 59726 99200 59782 100000 6 dout0[22]
port 181 nsew signal input
rlabel metal2 s 60554 99200 60610 100000 6 dout0[23]
port 182 nsew signal input
rlabel metal2 s 61382 99200 61438 100000 6 dout0[24]
port 183 nsew signal input
rlabel metal2 s 62302 99200 62358 100000 6 dout0[25]
port 184 nsew signal input
rlabel metal2 s 63130 99200 63186 100000 6 dout0[26]
port 185 nsew signal input
rlabel metal2 s 63958 99200 64014 100000 6 dout0[27]
port 186 nsew signal input
rlabel metal2 s 64878 99200 64934 100000 6 dout0[28]
port 187 nsew signal input
rlabel metal2 s 65706 99200 65762 100000 6 dout0[29]
port 188 nsew signal input
rlabel metal2 s 42522 99200 42578 100000 6 dout0[2]
port 189 nsew signal input
rlabel metal2 s 66534 99200 66590 100000 6 dout0[30]
port 190 nsew signal input
rlabel metal2 s 67454 99200 67510 100000 6 dout0[31]
port 191 nsew signal input
rlabel metal2 s 68282 99200 68338 100000 6 dout0[32]
port 192 nsew signal input
rlabel metal2 s 69110 99200 69166 100000 6 dout0[33]
port 193 nsew signal input
rlabel metal2 s 70030 99200 70086 100000 6 dout0[34]
port 194 nsew signal input
rlabel metal2 s 70858 99200 70914 100000 6 dout0[35]
port 195 nsew signal input
rlabel metal2 s 71778 99200 71834 100000 6 dout0[36]
port 196 nsew signal input
rlabel metal2 s 72606 99200 72662 100000 6 dout0[37]
port 197 nsew signal input
rlabel metal2 s 73434 99200 73490 100000 6 dout0[38]
port 198 nsew signal input
rlabel metal2 s 74354 99200 74410 100000 6 dout0[39]
port 199 nsew signal input
rlabel metal2 s 43350 99200 43406 100000 6 dout0[3]
port 200 nsew signal input
rlabel metal2 s 75182 99200 75238 100000 6 dout0[40]
port 201 nsew signal input
rlabel metal2 s 76010 99200 76066 100000 6 dout0[41]
port 202 nsew signal input
rlabel metal2 s 76930 99200 76986 100000 6 dout0[42]
port 203 nsew signal input
rlabel metal2 s 77758 99200 77814 100000 6 dout0[43]
port 204 nsew signal input
rlabel metal2 s 78586 99200 78642 100000 6 dout0[44]
port 205 nsew signal input
rlabel metal2 s 79506 99200 79562 100000 6 dout0[45]
port 206 nsew signal input
rlabel metal2 s 80334 99200 80390 100000 6 dout0[46]
port 207 nsew signal input
rlabel metal2 s 81162 99200 81218 100000 6 dout0[47]
port 208 nsew signal input
rlabel metal2 s 82082 99200 82138 100000 6 dout0[48]
port 209 nsew signal input
rlabel metal2 s 82910 99200 82966 100000 6 dout0[49]
port 210 nsew signal input
rlabel metal2 s 44178 99200 44234 100000 6 dout0[4]
port 211 nsew signal input
rlabel metal2 s 83738 99200 83794 100000 6 dout0[50]
port 212 nsew signal input
rlabel metal2 s 84658 99200 84714 100000 6 dout0[51]
port 213 nsew signal input
rlabel metal2 s 85486 99200 85542 100000 6 dout0[52]
port 214 nsew signal input
rlabel metal2 s 86314 99200 86370 100000 6 dout0[53]
port 215 nsew signal input
rlabel metal2 s 87234 99200 87290 100000 6 dout0[54]
port 216 nsew signal input
rlabel metal2 s 88062 99200 88118 100000 6 dout0[55]
port 217 nsew signal input
rlabel metal2 s 88890 99200 88946 100000 6 dout0[56]
port 218 nsew signal input
rlabel metal2 s 89810 99200 89866 100000 6 dout0[57]
port 219 nsew signal input
rlabel metal2 s 90638 99200 90694 100000 6 dout0[58]
port 220 nsew signal input
rlabel metal2 s 91558 99200 91614 100000 6 dout0[59]
port 221 nsew signal input
rlabel metal2 s 45098 99200 45154 100000 6 dout0[5]
port 222 nsew signal input
rlabel metal2 s 92386 99200 92442 100000 6 dout0[60]
port 223 nsew signal input
rlabel metal2 s 93214 99200 93270 100000 6 dout0[61]
port 224 nsew signal input
rlabel metal2 s 94134 99200 94190 100000 6 dout0[62]
port 225 nsew signal input
rlabel metal2 s 94962 99200 95018 100000 6 dout0[63]
port 226 nsew signal input
rlabel metal2 s 45926 99200 45982 100000 6 dout0[6]
port 227 nsew signal input
rlabel metal2 s 46754 99200 46810 100000 6 dout0[7]
port 228 nsew signal input
rlabel metal2 s 47674 99200 47730 100000 6 dout0[8]
port 229 nsew signal input
rlabel metal2 s 48502 99200 48558 100000 6 dout0[9]
port 230 nsew signal input
rlabel metal2 s 104438 99200 104494 100000 6 dout1[0]
port 231 nsew signal input
rlabel metal2 s 112994 99200 113050 100000 6 dout1[10]
port 232 nsew signal input
rlabel metal2 s 113914 99200 113970 100000 6 dout1[11]
port 233 nsew signal input
rlabel metal2 s 114742 99200 114798 100000 6 dout1[12]
port 234 nsew signal input
rlabel metal2 s 115570 99200 115626 100000 6 dout1[13]
port 235 nsew signal input
rlabel metal2 s 116490 99200 116546 100000 6 dout1[14]
port 236 nsew signal input
rlabel metal2 s 117318 99200 117374 100000 6 dout1[15]
port 237 nsew signal input
rlabel metal2 s 118146 99200 118202 100000 6 dout1[16]
port 238 nsew signal input
rlabel metal2 s 119066 99200 119122 100000 6 dout1[17]
port 239 nsew signal input
rlabel metal2 s 119894 99200 119950 100000 6 dout1[18]
port 240 nsew signal input
rlabel metal2 s 120722 99200 120778 100000 6 dout1[19]
port 241 nsew signal input
rlabel metal2 s 105266 99200 105322 100000 6 dout1[1]
port 242 nsew signal input
rlabel metal2 s 121642 99200 121698 100000 6 dout1[20]
port 243 nsew signal input
rlabel metal2 s 122470 99200 122526 100000 6 dout1[21]
port 244 nsew signal input
rlabel metal2 s 123298 99200 123354 100000 6 dout1[22]
port 245 nsew signal input
rlabel metal2 s 124218 99200 124274 100000 6 dout1[23]
port 246 nsew signal input
rlabel metal2 s 125046 99200 125102 100000 6 dout1[24]
port 247 nsew signal input
rlabel metal2 s 125966 99200 126022 100000 6 dout1[25]
port 248 nsew signal input
rlabel metal2 s 126794 99200 126850 100000 6 dout1[26]
port 249 nsew signal input
rlabel metal2 s 127622 99200 127678 100000 6 dout1[27]
port 250 nsew signal input
rlabel metal2 s 128542 99200 128598 100000 6 dout1[28]
port 251 nsew signal input
rlabel metal2 s 129370 99200 129426 100000 6 dout1[29]
port 252 nsew signal input
rlabel metal2 s 106094 99200 106150 100000 6 dout1[2]
port 253 nsew signal input
rlabel metal2 s 130198 99200 130254 100000 6 dout1[30]
port 254 nsew signal input
rlabel metal2 s 131118 99200 131174 100000 6 dout1[31]
port 255 nsew signal input
rlabel metal2 s 131946 99200 132002 100000 6 dout1[32]
port 256 nsew signal input
rlabel metal2 s 132774 99200 132830 100000 6 dout1[33]
port 257 nsew signal input
rlabel metal2 s 133694 99200 133750 100000 6 dout1[34]
port 258 nsew signal input
rlabel metal2 s 134522 99200 134578 100000 6 dout1[35]
port 259 nsew signal input
rlabel metal2 s 135350 99200 135406 100000 6 dout1[36]
port 260 nsew signal input
rlabel metal2 s 136270 99200 136326 100000 6 dout1[37]
port 261 nsew signal input
rlabel metal2 s 137098 99200 137154 100000 6 dout1[38]
port 262 nsew signal input
rlabel metal2 s 137926 99200 137982 100000 6 dout1[39]
port 263 nsew signal input
rlabel metal2 s 107014 99200 107070 100000 6 dout1[3]
port 264 nsew signal input
rlabel metal2 s 138846 99200 138902 100000 6 dout1[40]
port 265 nsew signal input
rlabel metal2 s 139674 99200 139730 100000 6 dout1[41]
port 266 nsew signal input
rlabel metal2 s 140502 99200 140558 100000 6 dout1[42]
port 267 nsew signal input
rlabel metal2 s 141422 99200 141478 100000 6 dout1[43]
port 268 nsew signal input
rlabel metal2 s 142250 99200 142306 100000 6 dout1[44]
port 269 nsew signal input
rlabel metal2 s 143170 99200 143226 100000 6 dout1[45]
port 270 nsew signal input
rlabel metal2 s 143998 99200 144054 100000 6 dout1[46]
port 271 nsew signal input
rlabel metal2 s 144826 99200 144882 100000 6 dout1[47]
port 272 nsew signal input
rlabel metal2 s 145746 99200 145802 100000 6 dout1[48]
port 273 nsew signal input
rlabel metal2 s 146574 99200 146630 100000 6 dout1[49]
port 274 nsew signal input
rlabel metal2 s 107842 99200 107898 100000 6 dout1[4]
port 275 nsew signal input
rlabel metal2 s 147402 99200 147458 100000 6 dout1[50]
port 276 nsew signal input
rlabel metal2 s 148322 99200 148378 100000 6 dout1[51]
port 277 nsew signal input
rlabel metal2 s 149150 99200 149206 100000 6 dout1[52]
port 278 nsew signal input
rlabel metal2 s 149978 99200 150034 100000 6 dout1[53]
port 279 nsew signal input
rlabel metal2 s 150898 99200 150954 100000 6 dout1[54]
port 280 nsew signal input
rlabel metal2 s 151726 99200 151782 100000 6 dout1[55]
port 281 nsew signal input
rlabel metal2 s 152554 99200 152610 100000 6 dout1[56]
port 282 nsew signal input
rlabel metal2 s 153474 99200 153530 100000 6 dout1[57]
port 283 nsew signal input
rlabel metal2 s 154302 99200 154358 100000 6 dout1[58]
port 284 nsew signal input
rlabel metal2 s 155130 99200 155186 100000 6 dout1[59]
port 285 nsew signal input
rlabel metal2 s 108762 99200 108818 100000 6 dout1[5]
port 286 nsew signal input
rlabel metal2 s 156050 99200 156106 100000 6 dout1[60]
port 287 nsew signal input
rlabel metal2 s 156878 99200 156934 100000 6 dout1[61]
port 288 nsew signal input
rlabel metal2 s 157706 99200 157762 100000 6 dout1[62]
port 289 nsew signal input
rlabel metal2 s 158626 99200 158682 100000 6 dout1[63]
port 290 nsew signal input
rlabel metal2 s 109590 99200 109646 100000 6 dout1[6]
port 291 nsew signal input
rlabel metal2 s 110418 99200 110474 100000 6 dout1[7]
port 292 nsew signal input
rlabel metal2 s 111338 99200 111394 100000 6 dout1[8]
port 293 nsew signal input
rlabel metal2 s 112166 99200 112222 100000 6 dout1[9]
port 294 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 jtag_tck
port 295 nsew signal input
rlabel metal2 s 159454 99200 159510 100000 6 jtag_tdi
port 296 nsew signal input
rlabel metal3 s 159200 97656 160000 97776 6 jtag_tdo
port 297 nsew signal output
rlabel metal3 s 159200 98064 160000 98184 6 jtag_tms
port 298 nsew signal input
rlabel metal3 s 159200 50328 160000 50448 6 localMemory_wb_ack_o
port 299 nsew signal output
rlabel metal3 s 159200 53184 160000 53304 6 localMemory_wb_adr_i[0]
port 300 nsew signal input
rlabel metal3 s 159200 69640 160000 69760 6 localMemory_wb_adr_i[10]
port 301 nsew signal input
rlabel metal3 s 159200 71000 160000 71120 6 localMemory_wb_adr_i[11]
port 302 nsew signal input
rlabel metal3 s 159200 72496 160000 72616 6 localMemory_wb_adr_i[12]
port 303 nsew signal input
rlabel metal3 s 159200 73992 160000 74112 6 localMemory_wb_adr_i[13]
port 304 nsew signal input
rlabel metal3 s 159200 75352 160000 75472 6 localMemory_wb_adr_i[14]
port 305 nsew signal input
rlabel metal3 s 159200 76848 160000 76968 6 localMemory_wb_adr_i[15]
port 306 nsew signal input
rlabel metal3 s 159200 78344 160000 78464 6 localMemory_wb_adr_i[16]
port 307 nsew signal input
rlabel metal3 s 159200 79704 160000 79824 6 localMemory_wb_adr_i[17]
port 308 nsew signal input
rlabel metal3 s 159200 81200 160000 81320 6 localMemory_wb_adr_i[18]
port 309 nsew signal input
rlabel metal3 s 159200 82696 160000 82816 6 localMemory_wb_adr_i[19]
port 310 nsew signal input
rlabel metal3 s 159200 55088 160000 55208 6 localMemory_wb_adr_i[1]
port 311 nsew signal input
rlabel metal3 s 159200 84056 160000 84176 6 localMemory_wb_adr_i[20]
port 312 nsew signal input
rlabel metal3 s 159200 85552 160000 85672 6 localMemory_wb_adr_i[21]
port 313 nsew signal input
rlabel metal3 s 159200 87048 160000 87168 6 localMemory_wb_adr_i[22]
port 314 nsew signal input
rlabel metal3 s 159200 88408 160000 88528 6 localMemory_wb_adr_i[23]
port 315 nsew signal input
rlabel metal3 s 159200 56992 160000 57112 6 localMemory_wb_adr_i[2]
port 316 nsew signal input
rlabel metal3 s 159200 59032 160000 59152 6 localMemory_wb_adr_i[3]
port 317 nsew signal input
rlabel metal3 s 159200 60936 160000 61056 6 localMemory_wb_adr_i[4]
port 318 nsew signal input
rlabel metal3 s 159200 62432 160000 62552 6 localMemory_wb_adr_i[5]
port 319 nsew signal input
rlabel metal3 s 159200 63792 160000 63912 6 localMemory_wb_adr_i[6]
port 320 nsew signal input
rlabel metal3 s 159200 65288 160000 65408 6 localMemory_wb_adr_i[7]
port 321 nsew signal input
rlabel metal3 s 159200 66784 160000 66904 6 localMemory_wb_adr_i[8]
port 322 nsew signal input
rlabel metal3 s 159200 68144 160000 68264 6 localMemory_wb_adr_i[9]
port 323 nsew signal input
rlabel metal3 s 159200 50736 160000 50856 6 localMemory_wb_cyc_i
port 324 nsew signal input
rlabel metal3 s 159200 53728 160000 53848 6 localMemory_wb_data_i[0]
port 325 nsew signal input
rlabel metal3 s 159200 70048 160000 70168 6 localMemory_wb_data_i[10]
port 326 nsew signal input
rlabel metal3 s 159200 71544 160000 71664 6 localMemory_wb_data_i[11]
port 327 nsew signal input
rlabel metal3 s 159200 73040 160000 73160 6 localMemory_wb_data_i[12]
port 328 nsew signal input
rlabel metal3 s 159200 74400 160000 74520 6 localMemory_wb_data_i[13]
port 329 nsew signal input
rlabel metal3 s 159200 75896 160000 76016 6 localMemory_wb_data_i[14]
port 330 nsew signal input
rlabel metal3 s 159200 77392 160000 77512 6 localMemory_wb_data_i[15]
port 331 nsew signal input
rlabel metal3 s 159200 78752 160000 78872 6 localMemory_wb_data_i[16]
port 332 nsew signal input
rlabel metal3 s 159200 80248 160000 80368 6 localMemory_wb_data_i[17]
port 333 nsew signal input
rlabel metal3 s 159200 81744 160000 81864 6 localMemory_wb_data_i[18]
port 334 nsew signal input
rlabel metal3 s 159200 83104 160000 83224 6 localMemory_wb_data_i[19]
port 335 nsew signal input
rlabel metal3 s 159200 55632 160000 55752 6 localMemory_wb_data_i[1]
port 336 nsew signal input
rlabel metal3 s 159200 84600 160000 84720 6 localMemory_wb_data_i[20]
port 337 nsew signal input
rlabel metal3 s 159200 86096 160000 86216 6 localMemory_wb_data_i[21]
port 338 nsew signal input
rlabel metal3 s 159200 87456 160000 87576 6 localMemory_wb_data_i[22]
port 339 nsew signal input
rlabel metal3 s 159200 88952 160000 89072 6 localMemory_wb_data_i[23]
port 340 nsew signal input
rlabel metal3 s 159200 89904 160000 90024 6 localMemory_wb_data_i[24]
port 341 nsew signal input
rlabel metal3 s 159200 90856 160000 90976 6 localMemory_wb_data_i[25]
port 342 nsew signal input
rlabel metal3 s 159200 91808 160000 91928 6 localMemory_wb_data_i[26]
port 343 nsew signal input
rlabel metal3 s 159200 92760 160000 92880 6 localMemory_wb_data_i[27]
port 344 nsew signal input
rlabel metal3 s 159200 93712 160000 93832 6 localMemory_wb_data_i[28]
port 345 nsew signal input
rlabel metal3 s 159200 94664 160000 94784 6 localMemory_wb_data_i[29]
port 346 nsew signal input
rlabel metal3 s 159200 57536 160000 57656 6 localMemory_wb_data_i[2]
port 347 nsew signal input
rlabel metal3 s 159200 95752 160000 95872 6 localMemory_wb_data_i[30]
port 348 nsew signal input
rlabel metal3 s 159200 96704 160000 96824 6 localMemory_wb_data_i[31]
port 349 nsew signal input
rlabel metal3 s 159200 59440 160000 59560 6 localMemory_wb_data_i[3]
port 350 nsew signal input
rlabel metal3 s 159200 61344 160000 61464 6 localMemory_wb_data_i[4]
port 351 nsew signal input
rlabel metal3 s 159200 62840 160000 62960 6 localMemory_wb_data_i[5]
port 352 nsew signal input
rlabel metal3 s 159200 64336 160000 64456 6 localMemory_wb_data_i[6]
port 353 nsew signal input
rlabel metal3 s 159200 65696 160000 65816 6 localMemory_wb_data_i[7]
port 354 nsew signal input
rlabel metal3 s 159200 67192 160000 67312 6 localMemory_wb_data_i[8]
port 355 nsew signal input
rlabel metal3 s 159200 68688 160000 68808 6 localMemory_wb_data_i[9]
port 356 nsew signal input
rlabel metal3 s 159200 54136 160000 54256 6 localMemory_wb_data_o[0]
port 357 nsew signal output
rlabel metal3 s 159200 70592 160000 70712 6 localMemory_wb_data_o[10]
port 358 nsew signal output
rlabel metal3 s 159200 72088 160000 72208 6 localMemory_wb_data_o[11]
port 359 nsew signal output
rlabel metal3 s 159200 73448 160000 73568 6 localMemory_wb_data_o[12]
port 360 nsew signal output
rlabel metal3 s 159200 74944 160000 75064 6 localMemory_wb_data_o[13]
port 361 nsew signal output
rlabel metal3 s 159200 76440 160000 76560 6 localMemory_wb_data_o[14]
port 362 nsew signal output
rlabel metal3 s 159200 77800 160000 77920 6 localMemory_wb_data_o[15]
port 363 nsew signal output
rlabel metal3 s 159200 79296 160000 79416 6 localMemory_wb_data_o[16]
port 364 nsew signal output
rlabel metal3 s 159200 80656 160000 80776 6 localMemory_wb_data_o[17]
port 365 nsew signal output
rlabel metal3 s 159200 82152 160000 82272 6 localMemory_wb_data_o[18]
port 366 nsew signal output
rlabel metal3 s 159200 83648 160000 83768 6 localMemory_wb_data_o[19]
port 367 nsew signal output
rlabel metal3 s 159200 56040 160000 56160 6 localMemory_wb_data_o[1]
port 368 nsew signal output
rlabel metal3 s 159200 85008 160000 85128 6 localMemory_wb_data_o[20]
port 369 nsew signal output
rlabel metal3 s 159200 86504 160000 86624 6 localMemory_wb_data_o[21]
port 370 nsew signal output
rlabel metal3 s 159200 88000 160000 88120 6 localMemory_wb_data_o[22]
port 371 nsew signal output
rlabel metal3 s 159200 89360 160000 89480 6 localMemory_wb_data_o[23]
port 372 nsew signal output
rlabel metal3 s 159200 90312 160000 90432 6 localMemory_wb_data_o[24]
port 373 nsew signal output
rlabel metal3 s 159200 91400 160000 91520 6 localMemory_wb_data_o[25]
port 374 nsew signal output
rlabel metal3 s 159200 92352 160000 92472 6 localMemory_wb_data_o[26]
port 375 nsew signal output
rlabel metal3 s 159200 93304 160000 93424 6 localMemory_wb_data_o[27]
port 376 nsew signal output
rlabel metal3 s 159200 94256 160000 94376 6 localMemory_wb_data_o[28]
port 377 nsew signal output
rlabel metal3 s 159200 95208 160000 95328 6 localMemory_wb_data_o[29]
port 378 nsew signal output
rlabel metal3 s 159200 58080 160000 58200 6 localMemory_wb_data_o[2]
port 379 nsew signal output
rlabel metal3 s 159200 96160 160000 96280 6 localMemory_wb_data_o[30]
port 380 nsew signal output
rlabel metal3 s 159200 97112 160000 97232 6 localMemory_wb_data_o[31]
port 381 nsew signal output
rlabel metal3 s 159200 59984 160000 60104 6 localMemory_wb_data_o[3]
port 382 nsew signal output
rlabel metal3 s 159200 61888 160000 62008 6 localMemory_wb_data_o[4]
port 383 nsew signal output
rlabel metal3 s 159200 63384 160000 63504 6 localMemory_wb_data_o[5]
port 384 nsew signal output
rlabel metal3 s 159200 64744 160000 64864 6 localMemory_wb_data_o[6]
port 385 nsew signal output
rlabel metal3 s 159200 66240 160000 66360 6 localMemory_wb_data_o[7]
port 386 nsew signal output
rlabel metal3 s 159200 67736 160000 67856 6 localMemory_wb_data_o[8]
port 387 nsew signal output
rlabel metal3 s 159200 69096 160000 69216 6 localMemory_wb_data_o[9]
port 388 nsew signal output
rlabel metal3 s 159200 51280 160000 51400 6 localMemory_wb_error_o
port 389 nsew signal output
rlabel metal3 s 159200 54680 160000 54800 6 localMemory_wb_sel_i[0]
port 390 nsew signal input
rlabel metal3 s 159200 56584 160000 56704 6 localMemory_wb_sel_i[1]
port 391 nsew signal input
rlabel metal3 s 159200 58488 160000 58608 6 localMemory_wb_sel_i[2]
port 392 nsew signal input
rlabel metal3 s 159200 60392 160000 60512 6 localMemory_wb_sel_i[3]
port 393 nsew signal input
rlabel metal3 s 159200 51688 160000 51808 6 localMemory_wb_stall_o
port 394 nsew signal output
rlabel metal3 s 159200 52232 160000 52352 6 localMemory_wb_stb_i
port 395 nsew signal input
rlabel metal3 s 159200 52776 160000 52896 6 localMemory_wb_we_i
port 396 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 manufacturerID[0]
port 397 nsew signal input
rlabel metal2 s 73894 0 73950 800 6 manufacturerID[10]
port 398 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 manufacturerID[1]
port 399 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 manufacturerID[2]
port 400 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 manufacturerID[3]
port 401 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 manufacturerID[4]
port 402 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 manufacturerID[5]
port 403 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 manufacturerID[6]
port 404 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 manufacturerID[7]
port 405 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 manufacturerID[8]
port 406 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 manufacturerID[9]
port 407 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 partID[0]
port 408 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 partID[10]
port 409 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 partID[11]
port 410 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 partID[12]
port 411 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 partID[13]
port 412 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 partID[14]
port 413 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 partID[15]
port 414 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 partID[1]
port 415 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 partID[2]
port 416 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 partID[3]
port 417 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 partID[4]
port 418 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 partID[5]
port 419 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 partID[6]
port 420 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 partID[7]
port 421 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 partID[8]
port 422 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 partID[9]
port 423 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 probe_errorCode[0]
port 424 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 probe_errorCode[1]
port 425 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 probe_errorCode[2]
port 426 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 probe_errorCode[3]
port 427 nsew signal output
rlabel metal3 s 0 824 800 944 6 probe_isBranch
port 428 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 probe_isCompressed
port 429 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 probe_isLoad
port 430 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 probe_isStore
port 431 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 probe_jtagInstruction[0]
port 432 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 probe_jtagInstruction[1]
port 433 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 probe_jtagInstruction[2]
port 434 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 probe_jtagInstruction[3]
port 435 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 probe_jtagInstruction[4]
port 436 nsew signal output
rlabel metal3 s 0 13200 800 13320 6 probe_opcode[0]
port 437 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 probe_opcode[1]
port 438 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 probe_opcode[2]
port 439 nsew signal output
rlabel metal3 s 0 38224 800 38344 6 probe_opcode[3]
port 440 nsew signal output
rlabel metal3 s 0 43664 800 43784 6 probe_opcode[4]
port 441 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 probe_opcode[5]
port 442 nsew signal output
rlabel metal3 s 0 50736 800 50856 6 probe_opcode[6]
port 443 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 probe_programCounter[0]
port 444 nsew signal output
rlabel metal3 s 0 59712 800 59832 6 probe_programCounter[10]
port 445 nsew signal output
rlabel metal3 s 0 61480 800 61600 6 probe_programCounter[11]
port 446 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 probe_programCounter[12]
port 447 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 probe_programCounter[13]
port 448 nsew signal output
rlabel metal3 s 0 66784 800 66904 6 probe_programCounter[14]
port 449 nsew signal output
rlabel metal3 s 0 68552 800 68672 6 probe_programCounter[15]
port 450 nsew signal output
rlabel metal3 s 0 70320 800 70440 6 probe_programCounter[16]
port 451 nsew signal output
rlabel metal3 s 0 72224 800 72344 6 probe_programCounter[17]
port 452 nsew signal output
rlabel metal3 s 0 73992 800 74112 6 probe_programCounter[18]
port 453 nsew signal output
rlabel metal3 s 0 75760 800 75880 6 probe_programCounter[19]
port 454 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 probe_programCounter[1]
port 455 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 probe_programCounter[20]
port 456 nsew signal output
rlabel metal3 s 0 79296 800 79416 6 probe_programCounter[21]
port 457 nsew signal output
rlabel metal3 s 0 81064 800 81184 6 probe_programCounter[22]
port 458 nsew signal output
rlabel metal3 s 0 82832 800 82952 6 probe_programCounter[23]
port 459 nsew signal output
rlabel metal3 s 0 84600 800 84720 6 probe_programCounter[24]
port 460 nsew signal output
rlabel metal3 s 0 86504 800 86624 6 probe_programCounter[25]
port 461 nsew signal output
rlabel metal3 s 0 88272 800 88392 6 probe_programCounter[26]
port 462 nsew signal output
rlabel metal3 s 0 90040 800 90160 6 probe_programCounter[27]
port 463 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 probe_programCounter[28]
port 464 nsew signal output
rlabel metal3 s 0 93576 800 93696 6 probe_programCounter[29]
port 465 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 probe_programCounter[2]
port 466 nsew signal output
rlabel metal3 s 0 95344 800 95464 6 probe_programCounter[30]
port 467 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 probe_programCounter[31]
port 468 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 probe_programCounter[3]
port 469 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 probe_programCounter[4]
port 470 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 probe_programCounter[5]
port 471 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 probe_programCounter[6]
port 472 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 probe_programCounter[7]
port 473 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 probe_programCounter[8]
port 474 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 probe_programCounter[9]
port 475 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 probe_state[0]
port 476 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 probe_state[1]
port 477 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 probe_takeBranch
port 478 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 97424 6 vccd1
port 479 nsew power bidirectional
rlabel metal2 s 141882 0 141938 800 6 versionID[0]
port 480 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 versionID[1]
port 481 nsew signal input
rlabel metal2 s 149886 0 149942 800 6 versionID[2]
port 482 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 versionID[3]
port 483 nsew signal input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 97424 6 vssd1
port 484 nsew ground bidirectional
rlabel metal3 s 159200 144 160000 264 6 wb_clk_i
port 485 nsew signal input
rlabel metal3 s 159200 552 160000 672 6 wb_rst_i
port 486 nsew signal input
rlabel metal2 s 1214 99200 1270 100000 6 web0
port 487 nsew signal output
rlabel metal2 s 2042 99200 2098 100000 6 wmask0[0]
port 488 nsew signal output
rlabel metal2 s 2962 99200 3018 100000 6 wmask0[1]
port 489 nsew signal output
rlabel metal2 s 3790 99200 3846 100000 6 wmask0[2]
port 490 nsew signal output
rlabel metal2 s 4618 99200 4674 100000 6 wmask0[3]
port 491 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 160000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 30748496
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/ExperiarCore/runs/ExperiarCore/results/signoff/ExperiarCore.magic.gds
string GDS_START 1371514
<< end >>

