VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO UART
  CLASS BLOCK ;
  FOREIGN UART ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END clk
  PIN peripheralBus_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END peripheralBus_address[0]
  PIN peripheralBus_address[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END peripheralBus_address[10]
  PIN peripheralBus_address[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END peripheralBus_address[11]
  PIN peripheralBus_address[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END peripheralBus_address[12]
  PIN peripheralBus_address[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END peripheralBus_address[13]
  PIN peripheralBus_address[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END peripheralBus_address[14]
  PIN peripheralBus_address[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END peripheralBus_address[15]
  PIN peripheralBus_address[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END peripheralBus_address[16]
  PIN peripheralBus_address[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END peripheralBus_address[17]
  PIN peripheralBus_address[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END peripheralBus_address[18]
  PIN peripheralBus_address[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END peripheralBus_address[19]
  PIN peripheralBus_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END peripheralBus_address[1]
  PIN peripheralBus_address[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END peripheralBus_address[20]
  PIN peripheralBus_address[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END peripheralBus_address[21]
  PIN peripheralBus_address[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END peripheralBus_address[22]
  PIN peripheralBus_address[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END peripheralBus_address[23]
  PIN peripheralBus_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END peripheralBus_address[2]
  PIN peripheralBus_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END peripheralBus_address[3]
  PIN peripheralBus_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END peripheralBus_address[4]
  PIN peripheralBus_address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END peripheralBus_address[5]
  PIN peripheralBus_address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END peripheralBus_address[6]
  PIN peripheralBus_address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END peripheralBus_address[7]
  PIN peripheralBus_address[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END peripheralBus_address[8]
  PIN peripheralBus_address[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END peripheralBus_address[9]
  PIN peripheralBus_busy
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END peripheralBus_busy
  PIN peripheralBus_data[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END peripheralBus_data[0]
  PIN peripheralBus_data[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END peripheralBus_data[10]
  PIN peripheralBus_data[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END peripheralBus_data[11]
  PIN peripheralBus_data[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END peripheralBus_data[12]
  PIN peripheralBus_data[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END peripheralBus_data[13]
  PIN peripheralBus_data[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END peripheralBus_data[14]
  PIN peripheralBus_data[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END peripheralBus_data[15]
  PIN peripheralBus_data[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END peripheralBus_data[16]
  PIN peripheralBus_data[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END peripheralBus_data[17]
  PIN peripheralBus_data[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END peripheralBus_data[18]
  PIN peripheralBus_data[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END peripheralBus_data[19]
  PIN peripheralBus_data[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END peripheralBus_data[1]
  PIN peripheralBus_data[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END peripheralBus_data[20]
  PIN peripheralBus_data[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END peripheralBus_data[21]
  PIN peripheralBus_data[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END peripheralBus_data[22]
  PIN peripheralBus_data[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END peripheralBus_data[23]
  PIN peripheralBus_data[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END peripheralBus_data[24]
  PIN peripheralBus_data[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END peripheralBus_data[25]
  PIN peripheralBus_data[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END peripheralBus_data[26]
  PIN peripheralBus_data[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END peripheralBus_data[27]
  PIN peripheralBus_data[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END peripheralBus_data[28]
  PIN peripheralBus_data[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END peripheralBus_data[29]
  PIN peripheralBus_data[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END peripheralBus_data[2]
  PIN peripheralBus_data[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END peripheralBus_data[30]
  PIN peripheralBus_data[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END peripheralBus_data[31]
  PIN peripheralBus_data[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END peripheralBus_data[3]
  PIN peripheralBus_data[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END peripheralBus_data[4]
  PIN peripheralBus_data[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END peripheralBus_data[5]
  PIN peripheralBus_data[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END peripheralBus_data[6]
  PIN peripheralBus_data[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END peripheralBus_data[7]
  PIN peripheralBus_data[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END peripheralBus_data[8]
  PIN peripheralBus_data[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END peripheralBus_data[9]
  PIN peripheralBus_oe
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END peripheralBus_oe
  PIN peripheralBus_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END peripheralBus_we
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END rst
  PIN uart_en[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 14.320 350.000 14.920 ;
    END
  END uart_en[0]
  PIN uart_en[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 101.360 350.000 101.960 ;
    END
  END uart_en[1]
  PIN uart_en[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 189.080 350.000 189.680 ;
    END
  END uart_en[2]
  PIN uart_en[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 276.800 350.000 277.400 ;
    END
  END uart_en[3]
  PIN uart_rx[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 42.880 350.000 43.480 ;
    END
  END uart_rx[0]
  PIN uart_rx[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 130.600 350.000 131.200 ;
    END
  END uart_rx[1]
  PIN uart_rx[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 218.320 350.000 218.920 ;
    END
  END uart_rx[2]
  PIN uart_rx[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 306.040 350.000 306.640 ;
    END
  END uart_rx[3]
  PIN uart_tx[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 72.120 350.000 72.720 ;
    END
  END uart_tx[0]
  PIN uart_tx[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 159.840 350.000 160.440 ;
    END
  END uart_tx[1]
  PIN uart_tx[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 247.560 350.000 248.160 ;
    END
  END uart_tx[2]
  PIN uart_tx[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 335.280 350.000 335.880 ;
    END
  END uart_tx[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 5.520 10.640 344.080 337.520 ;
      LAYER met2 ;
        RECT 6.990 4.280 340.770 337.520 ;
        RECT 6.990 2.875 87.210 4.280 ;
        RECT 88.050 2.875 262.010 4.280 ;
        RECT 262.850 2.875 340.770 4.280 ;
      LAYER met3 ;
        RECT 4.000 336.280 346.000 337.445 ;
        RECT 4.000 335.600 345.600 336.280 ;
        RECT 4.400 334.880 345.600 335.600 ;
        RECT 4.400 334.200 346.000 334.880 ;
        RECT 4.000 330.160 346.000 334.200 ;
        RECT 4.400 328.760 346.000 330.160 ;
        RECT 4.000 324.040 346.000 328.760 ;
        RECT 4.400 322.640 346.000 324.040 ;
        RECT 4.000 317.920 346.000 322.640 ;
        RECT 4.400 316.520 346.000 317.920 ;
        RECT 4.000 311.800 346.000 316.520 ;
        RECT 4.400 310.400 346.000 311.800 ;
        RECT 4.000 307.040 346.000 310.400 ;
        RECT 4.000 306.360 345.600 307.040 ;
        RECT 4.400 305.640 345.600 306.360 ;
        RECT 4.400 304.960 346.000 305.640 ;
        RECT 4.000 300.240 346.000 304.960 ;
        RECT 4.400 298.840 346.000 300.240 ;
        RECT 4.000 294.120 346.000 298.840 ;
        RECT 4.400 292.720 346.000 294.120 ;
        RECT 4.000 288.000 346.000 292.720 ;
        RECT 4.400 286.600 346.000 288.000 ;
        RECT 4.000 282.560 346.000 286.600 ;
        RECT 4.400 281.160 346.000 282.560 ;
        RECT 4.000 277.800 346.000 281.160 ;
        RECT 4.000 276.440 345.600 277.800 ;
        RECT 4.400 276.400 345.600 276.440 ;
        RECT 4.400 275.040 346.000 276.400 ;
        RECT 4.000 270.320 346.000 275.040 ;
        RECT 4.400 268.920 346.000 270.320 ;
        RECT 4.000 264.880 346.000 268.920 ;
        RECT 4.400 263.480 346.000 264.880 ;
        RECT 4.000 258.760 346.000 263.480 ;
        RECT 4.400 257.360 346.000 258.760 ;
        RECT 4.000 252.640 346.000 257.360 ;
        RECT 4.400 251.240 346.000 252.640 ;
        RECT 4.000 248.560 346.000 251.240 ;
        RECT 4.000 247.160 345.600 248.560 ;
        RECT 4.000 246.520 346.000 247.160 ;
        RECT 4.400 245.120 346.000 246.520 ;
        RECT 4.000 241.080 346.000 245.120 ;
        RECT 4.400 239.680 346.000 241.080 ;
        RECT 4.000 234.960 346.000 239.680 ;
        RECT 4.400 233.560 346.000 234.960 ;
        RECT 4.000 228.840 346.000 233.560 ;
        RECT 4.400 227.440 346.000 228.840 ;
        RECT 4.000 222.720 346.000 227.440 ;
        RECT 4.400 221.320 346.000 222.720 ;
        RECT 4.000 219.320 346.000 221.320 ;
        RECT 4.000 217.920 345.600 219.320 ;
        RECT 4.000 217.280 346.000 217.920 ;
        RECT 4.400 215.880 346.000 217.280 ;
        RECT 4.000 211.160 346.000 215.880 ;
        RECT 4.400 209.760 346.000 211.160 ;
        RECT 4.000 205.040 346.000 209.760 ;
        RECT 4.400 203.640 346.000 205.040 ;
        RECT 4.000 199.600 346.000 203.640 ;
        RECT 4.400 198.200 346.000 199.600 ;
        RECT 4.000 193.480 346.000 198.200 ;
        RECT 4.400 192.080 346.000 193.480 ;
        RECT 4.000 190.080 346.000 192.080 ;
        RECT 4.000 188.680 345.600 190.080 ;
        RECT 4.000 187.360 346.000 188.680 ;
        RECT 4.400 185.960 346.000 187.360 ;
        RECT 4.000 181.240 346.000 185.960 ;
        RECT 4.400 179.840 346.000 181.240 ;
        RECT 4.000 175.800 346.000 179.840 ;
        RECT 4.400 174.400 346.000 175.800 ;
        RECT 4.000 169.680 346.000 174.400 ;
        RECT 4.400 168.280 346.000 169.680 ;
        RECT 4.000 163.560 346.000 168.280 ;
        RECT 4.400 162.160 346.000 163.560 ;
        RECT 4.000 160.840 346.000 162.160 ;
        RECT 4.000 159.440 345.600 160.840 ;
        RECT 4.000 157.440 346.000 159.440 ;
        RECT 4.400 156.040 346.000 157.440 ;
        RECT 4.000 152.000 346.000 156.040 ;
        RECT 4.400 150.600 346.000 152.000 ;
        RECT 4.000 145.880 346.000 150.600 ;
        RECT 4.400 144.480 346.000 145.880 ;
        RECT 4.000 139.760 346.000 144.480 ;
        RECT 4.400 138.360 346.000 139.760 ;
        RECT 4.000 134.320 346.000 138.360 ;
        RECT 4.400 132.920 346.000 134.320 ;
        RECT 4.000 131.600 346.000 132.920 ;
        RECT 4.000 130.200 345.600 131.600 ;
        RECT 4.000 128.200 346.000 130.200 ;
        RECT 4.400 126.800 346.000 128.200 ;
        RECT 4.000 122.080 346.000 126.800 ;
        RECT 4.400 120.680 346.000 122.080 ;
        RECT 4.000 115.960 346.000 120.680 ;
        RECT 4.400 114.560 346.000 115.960 ;
        RECT 4.000 110.520 346.000 114.560 ;
        RECT 4.400 109.120 346.000 110.520 ;
        RECT 4.000 104.400 346.000 109.120 ;
        RECT 4.400 103.000 346.000 104.400 ;
        RECT 4.000 102.360 346.000 103.000 ;
        RECT 4.000 100.960 345.600 102.360 ;
        RECT 4.000 98.280 346.000 100.960 ;
        RECT 4.400 96.880 346.000 98.280 ;
        RECT 4.000 92.160 346.000 96.880 ;
        RECT 4.400 90.760 346.000 92.160 ;
        RECT 4.000 86.720 346.000 90.760 ;
        RECT 4.400 85.320 346.000 86.720 ;
        RECT 4.000 80.600 346.000 85.320 ;
        RECT 4.400 79.200 346.000 80.600 ;
        RECT 4.000 74.480 346.000 79.200 ;
        RECT 4.400 73.120 346.000 74.480 ;
        RECT 4.400 73.080 345.600 73.120 ;
        RECT 4.000 71.720 345.600 73.080 ;
        RECT 4.000 69.040 346.000 71.720 ;
        RECT 4.400 67.640 346.000 69.040 ;
        RECT 4.000 62.920 346.000 67.640 ;
        RECT 4.400 61.520 346.000 62.920 ;
        RECT 4.000 56.800 346.000 61.520 ;
        RECT 4.400 55.400 346.000 56.800 ;
        RECT 4.000 50.680 346.000 55.400 ;
        RECT 4.400 49.280 346.000 50.680 ;
        RECT 4.000 45.240 346.000 49.280 ;
        RECT 4.400 43.880 346.000 45.240 ;
        RECT 4.400 43.840 345.600 43.880 ;
        RECT 4.000 42.480 345.600 43.840 ;
        RECT 4.000 39.120 346.000 42.480 ;
        RECT 4.400 37.720 346.000 39.120 ;
        RECT 4.000 33.000 346.000 37.720 ;
        RECT 4.400 31.600 346.000 33.000 ;
        RECT 4.000 26.880 346.000 31.600 ;
        RECT 4.400 25.480 346.000 26.880 ;
        RECT 4.000 21.440 346.000 25.480 ;
        RECT 4.400 20.040 346.000 21.440 ;
        RECT 4.000 15.320 346.000 20.040 ;
        RECT 4.400 13.920 345.600 15.320 ;
        RECT 4.000 9.200 346.000 13.920 ;
        RECT 4.400 7.800 346.000 9.200 ;
        RECT 4.000 3.760 346.000 7.800 ;
        RECT 4.400 2.895 346.000 3.760 ;
  END
END UART
END LIBRARY

