* NGSPICE file created from ExperiarCore.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

.subckt ExperiarCore addr0[0] addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6]
+ addr0[7] addr0[8] addr1[0] addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6]
+ addr1[7] addr1[8] clk0 clk1 coreIndex[0] coreIndex[1] coreIndex[2] coreIndex[3]
+ coreIndex[4] coreIndex[5] coreIndex[6] coreIndex[7] core_wb_ack_i core_wb_adr_o[0]
+ core_wb_adr_o[10] core_wb_adr_o[11] core_wb_adr_o[12] core_wb_adr_o[13] core_wb_adr_o[14]
+ core_wb_adr_o[15] core_wb_adr_o[16] core_wb_adr_o[17] core_wb_adr_o[18] core_wb_adr_o[19]
+ core_wb_adr_o[1] core_wb_adr_o[20] core_wb_adr_o[21] core_wb_adr_o[22] core_wb_adr_o[23]
+ core_wb_adr_o[24] core_wb_adr_o[25] core_wb_adr_o[26] core_wb_adr_o[27] core_wb_adr_o[2]
+ core_wb_adr_o[3] core_wb_adr_o[4] core_wb_adr_o[5] core_wb_adr_o[6] core_wb_adr_o[7]
+ core_wb_adr_o[8] core_wb_adr_o[9] core_wb_cyc_o core_wb_data_i[0] core_wb_data_i[10]
+ core_wb_data_i[11] core_wb_data_i[12] core_wb_data_i[13] core_wb_data_i[14] core_wb_data_i[15]
+ core_wb_data_i[16] core_wb_data_i[17] core_wb_data_i[18] core_wb_data_i[19] core_wb_data_i[1]
+ core_wb_data_i[20] core_wb_data_i[21] core_wb_data_i[22] core_wb_data_i[23] core_wb_data_i[24]
+ core_wb_data_i[25] core_wb_data_i[26] core_wb_data_i[27] core_wb_data_i[28] core_wb_data_i[29]
+ core_wb_data_i[2] core_wb_data_i[30] core_wb_data_i[31] core_wb_data_i[3] core_wb_data_i[4]
+ core_wb_data_i[5] core_wb_data_i[6] core_wb_data_i[7] core_wb_data_i[8] core_wb_data_i[9]
+ core_wb_data_o[0] core_wb_data_o[10] core_wb_data_o[11] core_wb_data_o[12] core_wb_data_o[13]
+ core_wb_data_o[14] core_wb_data_o[15] core_wb_data_o[16] core_wb_data_o[17] core_wb_data_o[18]
+ core_wb_data_o[19] core_wb_data_o[1] core_wb_data_o[20] core_wb_data_o[21] core_wb_data_o[22]
+ core_wb_data_o[23] core_wb_data_o[24] core_wb_data_o[25] core_wb_data_o[26] core_wb_data_o[27]
+ core_wb_data_o[28] core_wb_data_o[29] core_wb_data_o[2] core_wb_data_o[30] core_wb_data_o[31]
+ core_wb_data_o[3] core_wb_data_o[4] core_wb_data_o[5] core_wb_data_o[6] core_wb_data_o[7]
+ core_wb_data_o[8] core_wb_data_o[9] core_wb_error_i core_wb_sel_o[0] core_wb_sel_o[1]
+ core_wb_sel_o[2] core_wb_sel_o[3] core_wb_stall_i core_wb_stb_o core_wb_we_o csb0[0]
+ csb0[1] csb1[0] csb1[1] din0[0] din0[10] din0[11] din0[12] din0[13] din0[14] din0[15]
+ din0[16] din0[17] din0[18] din0[19] din0[1] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[2] din0[30] din0[31]
+ din0[3] din0[4] din0[5] din0[6] din0[7] din0[8] din0[9] dout0[0] dout0[10] dout0[11]
+ dout0[12] dout0[13] dout0[14] dout0[15] dout0[16] dout0[17] dout0[18] dout0[19]
+ dout0[1] dout0[20] dout0[21] dout0[22] dout0[23] dout0[24] dout0[25] dout0[26] dout0[27]
+ dout0[28] dout0[29] dout0[2] dout0[30] dout0[31] dout0[32] dout0[33] dout0[34] dout0[35]
+ dout0[36] dout0[37] dout0[38] dout0[39] dout0[3] dout0[40] dout0[41] dout0[42] dout0[43]
+ dout0[44] dout0[45] dout0[46] dout0[47] dout0[48] dout0[49] dout0[4] dout0[50] dout0[51]
+ dout0[52] dout0[53] dout0[54] dout0[55] dout0[56] dout0[57] dout0[58] dout0[59]
+ dout0[5] dout0[60] dout0[61] dout0[62] dout0[63] dout0[6] dout0[7] dout0[8] dout0[9]
+ dout1[0] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16] dout1[17]
+ dout1[18] dout1[19] dout1[1] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24] dout1[25]
+ dout1[26] dout1[27] dout1[28] dout1[29] dout1[2] dout1[30] dout1[31] dout1[32] dout1[33]
+ dout1[34] dout1[35] dout1[36] dout1[37] dout1[38] dout1[39] dout1[3] dout1[40] dout1[41]
+ dout1[42] dout1[43] dout1[44] dout1[45] dout1[46] dout1[47] dout1[48] dout1[49]
+ dout1[4] dout1[50] dout1[51] dout1[52] dout1[53] dout1[54] dout1[55] dout1[56] dout1[57]
+ dout1[58] dout1[59] dout1[5] dout1[60] dout1[61] dout1[62] dout1[63] dout1[6] dout1[7]
+ dout1[8] dout1[9] irq[0] irq[10] irq[11] irq[12] irq[13] irq[14] irq[15] irq[1]
+ irq[2] irq[3] irq[4] irq[5] irq[6] irq[7] irq[8] irq[9] jtag_tck jtag_tdi jtag_tdo
+ jtag_tms localMemory_wb_ack_o localMemory_wb_adr_i[0] localMemory_wb_adr_i[10] localMemory_wb_adr_i[11]
+ localMemory_wb_adr_i[12] localMemory_wb_adr_i[13] localMemory_wb_adr_i[14] localMemory_wb_adr_i[15]
+ localMemory_wb_adr_i[16] localMemory_wb_adr_i[17] localMemory_wb_adr_i[18] localMemory_wb_adr_i[19]
+ localMemory_wb_adr_i[1] localMemory_wb_adr_i[20] localMemory_wb_adr_i[21] localMemory_wb_adr_i[22]
+ localMemory_wb_adr_i[23] localMemory_wb_adr_i[2] localMemory_wb_adr_i[3] localMemory_wb_adr_i[4]
+ localMemory_wb_adr_i[5] localMemory_wb_adr_i[6] localMemory_wb_adr_i[7] localMemory_wb_adr_i[8]
+ localMemory_wb_adr_i[9] localMemory_wb_cyc_i localMemory_wb_data_i[0] localMemory_wb_data_i[10]
+ localMemory_wb_data_i[11] localMemory_wb_data_i[12] localMemory_wb_data_i[13] localMemory_wb_data_i[14]
+ localMemory_wb_data_i[15] localMemory_wb_data_i[16] localMemory_wb_data_i[17] localMemory_wb_data_i[18]
+ localMemory_wb_data_i[19] localMemory_wb_data_i[1] localMemory_wb_data_i[20] localMemory_wb_data_i[21]
+ localMemory_wb_data_i[22] localMemory_wb_data_i[23] localMemory_wb_data_i[24] localMemory_wb_data_i[25]
+ localMemory_wb_data_i[26] localMemory_wb_data_i[27] localMemory_wb_data_i[28] localMemory_wb_data_i[29]
+ localMemory_wb_data_i[2] localMemory_wb_data_i[30] localMemory_wb_data_i[31] localMemory_wb_data_i[3]
+ localMemory_wb_data_i[4] localMemory_wb_data_i[5] localMemory_wb_data_i[6] localMemory_wb_data_i[7]
+ localMemory_wb_data_i[8] localMemory_wb_data_i[9] localMemory_wb_data_o[0] localMemory_wb_data_o[10]
+ localMemory_wb_data_o[11] localMemory_wb_data_o[12] localMemory_wb_data_o[13] localMemory_wb_data_o[14]
+ localMemory_wb_data_o[15] localMemory_wb_data_o[16] localMemory_wb_data_o[17] localMemory_wb_data_o[18]
+ localMemory_wb_data_o[19] localMemory_wb_data_o[1] localMemory_wb_data_o[20] localMemory_wb_data_o[21]
+ localMemory_wb_data_o[22] localMemory_wb_data_o[23] localMemory_wb_data_o[24] localMemory_wb_data_o[25]
+ localMemory_wb_data_o[26] localMemory_wb_data_o[27] localMemory_wb_data_o[28] localMemory_wb_data_o[29]
+ localMemory_wb_data_o[2] localMemory_wb_data_o[30] localMemory_wb_data_o[31] localMemory_wb_data_o[3]
+ localMemory_wb_data_o[4] localMemory_wb_data_o[5] localMemory_wb_data_o[6] localMemory_wb_data_o[7]
+ localMemory_wb_data_o[8] localMemory_wb_data_o[9] localMemory_wb_error_o localMemory_wb_sel_i[0]
+ localMemory_wb_sel_i[1] localMemory_wb_sel_i[2] localMemory_wb_sel_i[3] localMemory_wb_stall_o
+ localMemory_wb_stb_i localMemory_wb_we_i manufacturerID[0] manufacturerID[10] manufacturerID[1]
+ manufacturerID[2] manufacturerID[3] manufacturerID[4] manufacturerID[5] manufacturerID[6]
+ manufacturerID[7] manufacturerID[8] manufacturerID[9] partID[0] partID[10] partID[11]
+ partID[12] partID[13] partID[14] partID[15] partID[1] partID[2] partID[3] partID[4]
+ partID[5] partID[6] partID[7] partID[8] partID[9] probe_env[0] probe_env[1] probe_jtagInstruction[0]
+ probe_jtagInstruction[1] probe_jtagInstruction[2] probe_jtagInstruction[3] probe_jtagInstruction[4]
+ probe_programCounter[0] probe_programCounter[10] probe_programCounter[11] probe_programCounter[12]
+ probe_programCounter[13] probe_programCounter[14] probe_programCounter[15] probe_programCounter[16]
+ probe_programCounter[17] probe_programCounter[18] probe_programCounter[19] probe_programCounter[1]
+ probe_programCounter[20] probe_programCounter[21] probe_programCounter[22] probe_programCounter[23]
+ probe_programCounter[24] probe_programCounter[25] probe_programCounter[26] probe_programCounter[27]
+ probe_programCounter[28] probe_programCounter[29] probe_programCounter[2] probe_programCounter[30]
+ probe_programCounter[31] probe_programCounter[3] probe_programCounter[4] probe_programCounter[5]
+ probe_programCounter[6] probe_programCounter[7] probe_programCounter[8] probe_programCounter[9]
+ probe_state vccd1 versionID[0] versionID[1] versionID[2] versionID[3] vssd1 wb_clk_i
+ wb_rst_i web0 wmask0[0] wmask0[1] wmask0[2] wmask0[3]
XFILLER_274_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09671_ input122/X input157/X _11241_/S vssd1 vssd1 vccd1 vccd1 _09672_/C sky130_fd_sc_hd__mux2_8
XFILLER_255_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18869_ _18511_/X _18937_/B _18867_/X _18868_/Y vssd1 vssd1 vccd1 vccd1 _18870_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20900_ _20998_/CLK _20900_/D vssd1 vssd1 vccd1 vccd1 _20900_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_270_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20831_ _21025_/CLK _20831_/D vssd1 vssd1 vccd1 vccd1 _20831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20762_ _20763_/CLK _20762_/D vssd1 vssd1 vccd1 vccd1 _20762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20693_ _20720_/CLK _20693_/D vssd1 vssd1 vccd1 vccd1 _20693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1807 _10284_/A vssd1 vssd1 vccd1 vccd1 _10373_/A sky130_fd_sc_hd__buf_8
Xfanout820 _15994_/B1 vssd1 vssd1 vccd1 vccd1 _16043_/B1 sky130_fd_sc_hd__buf_6
Xfanout1818 _19180_/Q vssd1 vssd1 vccd1 vccd1 _12512_/B sky130_fd_sc_hd__buf_6
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1829 _11670_/S vssd1 vssd1 vccd1 vccd1 _12513_/C sky130_fd_sc_hd__buf_12
X_20127_ _20438_/CLK _20127_/D vssd1 vssd1 vccd1 vccd1 _20127_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout831 _11785_/Y vssd1 vssd1 vccd1 vccd1 _13637_/A sky130_fd_sc_hd__buf_4
Xfanout842 _18375_/B vssd1 vssd1 vccd1 vccd1 _18385_/B sky130_fd_sc_hd__buf_4
X_09938_ _09939_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__or2_1
Xfanout853 _18157_/Y vssd1 vssd1 vccd1 vccd1 _18311_/S sky130_fd_sc_hd__buf_6
XFILLER_58_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout864 _15323_/A vssd1 vssd1 vccd1 vccd1 _15478_/C1 sky130_fd_sc_hd__buf_6
Xfanout875 _14948_/Y vssd1 vssd1 vccd1 vccd1 _15942_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_219_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20058_ _20690_/CLK _20058_/D vssd1 vssd1 vccd1 vccd1 _20058_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout886 _11018_/Y vssd1 vssd1 vccd1 vccd1 _14841_/S sky130_fd_sc_hd__buf_4
X_09869_ _12039_/A1 _10119_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _09869_/X sky130_fd_sc_hd__a21o_4
Xfanout897 _16718_/X vssd1 vssd1 vccd1 vccd1 _16974_/A1 sky130_fd_sc_hd__buf_6
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ _11898_/X _11899_/X _11902_/S vssd1 vssd1 vccd1 vccd1 _11900_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _12901_/B _12880_/B vssd1 vssd1 vccd1 vccd1 _12880_/X sky130_fd_sc_hd__or2_2
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_202 _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _19390_/Q _20681_/Q _12139_/S vssd1 vssd1 vccd1 vccd1 _11831_/X sky130_fd_sc_hd__mux2_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_224 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _19320_/Q _17938_/A1 _14558_/S vssd1 vssd1 vccd1 vccd1 _19320_/D sky130_fd_sc_hd__mux2_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11772_/A _11772_/B _13596_/A vssd1 vssd1 vccd1 vccd1 _11773_/A sky130_fd_sc_hd__o21bai_2
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_279 _20622_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13501_/A _13501_/B _13501_/C vssd1 vssd1 vccd1 vccd1 _13501_/X sky130_fd_sc_hd__or3_1
X_10713_ _12275_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10713_/Y sky130_fd_sc_hd__nor2_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14481_ _20236_/Q _19265_/Q _14483_/S vssd1 vssd1 vccd1 vccd1 _14482_/B sky130_fd_sc_hd__mux2_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _20168_/Q _11693_/B vssd1 vssd1 vccd1 vccd1 _11693_/X sky130_fd_sc_hd__or2_1
X_16220_ _19643_/Q _17872_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19643_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13432_ _13432_/A _13432_/B vssd1 vssd1 vccd1 vccd1 _15898_/A sky130_fd_sc_hd__xor2_4
X_10644_ _10456_/Y _10643_/Y _10640_/X vssd1 vssd1 vccd1 vccd1 _11405_/A sky130_fd_sc_hd__a21o_1
XFILLER_201_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16151_ _19599_/Q _16178_/S _16150_/Y _16165_/C1 vssd1 vssd1 vccd1 vccd1 _19599_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13363_ _20934_/Q _13363_/B vssd1 vssd1 vccd1 vccd1 _13363_/Y sky130_fd_sc_hd__nand2_1
X_10575_ _20566_/Q _12043_/B vssd1 vssd1 vccd1 vccd1 _10575_/X sky130_fd_sc_hd__or2_1
XFILLER_177_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15102_ _11189_/Y _15101_/X _15492_/A vssd1 vssd1 vccd1 vccd1 _15102_/Y sky130_fd_sc_hd__o21ai_1
X_12314_ _12241_/S _12313_/X _12312_/X _12314_/C1 vssd1 vssd1 vccd1 vccd1 _12314_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16082_ _19565_/Q _16081_/B _16081_/Y _16097_/B1 vssd1 vssd1 vccd1 vccd1 _19565_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13294_ _13289_/Y _13293_/X _14275_/A1 vssd1 vssd1 vccd1 vccd1 _13294_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_142_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19910_ _20694_/CLK _19910_/D vssd1 vssd1 vccd1 vccd1 _19910_/Q sky130_fd_sc_hd__dfxtp_1
X_15033_ _13637_/A _15032_/Y _14810_/X vssd1 vssd1 vccd1 vccd1 _15033_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_138_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12245_ _12245_/A1 _17949_/A1 _12244_/X _13675_/A vssd1 vssd1 vccd1 vccd1 _12245_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_181_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19841_ _19978_/CLK _19841_/D vssd1 vssd1 vccd1 vccd1 _19841_/Q sky130_fd_sc_hd__dfxtp_4
X_12176_ _11851_/C _12175_/X _12172_/X _12191_/C1 vssd1 vssd1 vccd1 vccd1 _12176_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11127_ _20152_/Q _11379_/B _12347_/C1 vssd1 vssd1 vccd1 vccd1 _11127_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19772_ _20084_/CLK _19772_/D vssd1 vssd1 vccd1 vccd1 _19772_/Q sky130_fd_sc_hd__dfxtp_1
X_16984_ _16950_/Y _16983_/X _16875_/B2 vssd1 vssd1 vccd1 vccd1 _16984_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11058_ _10553_/B _10470_/Y _11057_/X _10461_/X vssd1 vssd1 vccd1 vccd1 _11058_/Y
+ sky130_fd_sc_hd__o211ai_1
X_15935_ _20877_/Q _16042_/A2 fanout819/X vssd1 vssd1 vccd1 vccd1 _15935_/X sky130_fd_sc_hd__o21ba_1
X_18723_ _20962_/Q _18240_/Y _18749_/S vssd1 vssd1 vccd1 vccd1 _18724_/B sky130_fd_sc_hd__mux2_1
XFILLER_283_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20155_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10009_ _11948_/A1 _10008_/X _10007_/X vssd1 vssd1 vccd1 vccd1 _10009_/X sky130_fd_sc_hd__o21a_1
XFILLER_225_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18654_ _20937_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18654_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _15948_/A1 _12873_/X _15865_/X _15921_/B2 vssd1 vssd1 vccd1 vccd1 _15866_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_76_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17605_ _20363_/Q _17916_/A1 _17606_/S vssd1 vssd1 vccd1 vccd1 _20363_/D sky130_fd_sc_hd__mux2_1
X_14817_ _14813_/X _14816_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _14817_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18585_ _19499_/Q _18589_/B vssd1 vssd1 vccd1 vccd1 _18585_/Y sky130_fd_sc_hd__nand2_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15797_ _19724_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15797_/X sky130_fd_sc_hd__or2_1
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17536_ _20300_/Q _20299_/Q _20298_/Q _17536_/D vssd1 vssd1 vccd1 vccd1 _17537_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_178_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XExperiarCore_2007 vssd1 vssd1 vccd1 vccd1 ExperiarCore_2007/HI localMemory_wb_error_o
+ sky130_fd_sc_hd__conb_1
X_14748_ _19121_/Q _14764_/A2 _14747_/X _14758_/C1 vssd1 vssd1 vccd1 vccd1 _19498_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17467_ _17487_/A1 _17466_/Y _16451_/A vssd1 vssd1 vccd1 vccd1 _20268_/D sky130_fd_sc_hd__a21oi_1
X_14679_ _19438_/Q _17928_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19438_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19206_ _20426_/CLK _19206_/D vssd1 vssd1 vccd1 vccd1 _19206_/Q sky130_fd_sc_hd__dfxtp_1
X_16418_ _19751_/Q _19752_/Q _16418_/C vssd1 vssd1 vccd1 vccd1 _16420_/B sky130_fd_sc_hd__and3_4
XFILLER_149_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17398_ _20247_/Q _17337_/B _17530_/A2 _20296_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17398_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19137_ _19520_/CLK _19137_/D vssd1 vssd1 vccd1 vccd1 _19137_/Q sky130_fd_sc_hd__dfxtp_1
X_16349_ _19726_/Q _16348_/B _18720_/A vssd1 vssd1 vccd1 vccd1 _16350_/B sky130_fd_sc_hd__o21ai_1
XFILLER_145_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19068_ _20413_/Q vssd1 vssd1 vccd1 vccd1 _20413_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput401 _13794_/X vssd1 vssd1 vccd1 vccd1 din0[3] sky130_fd_sc_hd__buf_6
XFILLER_218_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput412 _19972_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[11] sky130_fd_sc_hd__buf_4
X_18019_ _20745_/Q _20744_/Q _18019_/C vssd1 vssd1 vccd1 vccd1 _18024_/C sky130_fd_sc_hd__and3_2
Xoutput423 _19982_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[21] sky130_fd_sc_hd__buf_4
XFILLER_161_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput434 _19992_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[31] sky130_fd_sc_hd__buf_4
XFILLER_114_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput445 _20257_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[0] sky130_fd_sc_hd__buf_4
Xoutput456 _19509_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[15] sky130_fd_sc_hd__buf_4
X_21030_ _21030_/CLK _21030_/D vssd1 vssd1 vccd1 vccd1 _21030_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput467 _19519_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[25] sky130_fd_sc_hd__buf_4
XFILLER_271_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput478 _19500_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[6] sky130_fd_sc_hd__buf_4
XFILLER_102_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09723_ _12144_/C1 _09712_/X _09715_/X _09722_/X _12152_/A1 vssd1 vssd1 vccd1 vccd1
+ _09723_/X sky130_fd_sc_hd__a311o_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09654_ _09681_/B _09681_/C _10553_/B vssd1 vssd1 vccd1 vccd1 _09678_/A sky130_fd_sc_hd__a21oi_1
XFILLER_243_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _09585_/A _19088_/Q _09585_/C _09606_/A vssd1 vssd1 vccd1 vccd1 _09596_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_83_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20814_ _21026_/CLK _20814_/D vssd1 vssd1 vccd1 vccd1 _20814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20745_ _21029_/CLK _20745_/D vssd1 vssd1 vccd1 vccd1 _20745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20676_ _20676_/CLK _20676_/D vssd1 vssd1 vccd1 vccd1 _20676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10360_ _12258_/S _10359_/X _11396_/S vssd1 vssd1 vccd1 vccd1 _10360_/X sky130_fd_sc_hd__o21a_1
XFILLER_136_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10291_ _10037_/Y _10290_/Y _09669_/X vssd1 vssd1 vccd1 vccd1 _10291_/X sky130_fd_sc_hd__a21o_1
XFILLER_275_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12030_ _12194_/A1 _17913_/A1 _12029_/X _09750_/Y vssd1 vssd1 vccd1 vccd1 _15931_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1604 _09618_/Y vssd1 vssd1 vccd1 vccd1 _12063_/C1 sky130_fd_sc_hd__buf_4
Xfanout1615 _11988_/S vssd1 vssd1 vccd1 vccd1 _12143_/S sky130_fd_sc_hd__buf_4
Xfanout1626 fanout1630/X vssd1 vssd1 vccd1 vccd1 _12376_/S sky130_fd_sc_hd__buf_8
XFILLER_132_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1637 _12400_/A1 vssd1 vssd1 vccd1 vccd1 _09689_/A sky130_fd_sc_hd__buf_8
XFILLER_104_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout650 _16067_/X vssd1 vssd1 vccd1 vccd1 _16077_/B sky130_fd_sc_hd__buf_2
XFILLER_219_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1648 _12531_/Y vssd1 vssd1 vccd1 vccd1 _18955_/A sky130_fd_sc_hd__buf_4
Xfanout1659 _09648_/Y vssd1 vssd1 vccd1 vccd1 _11239_/B1 sky130_fd_sc_hd__buf_8
XFILLER_219_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout661 _14737_/X vssd1 vssd1 vccd1 vccd1 _14773_/B sky130_fd_sc_hd__clkbuf_4
Xfanout672 _13906_/B vssd1 vssd1 vccd1 vccd1 _13921_/B sky130_fd_sc_hd__buf_4
XFILLER_120_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13981_ _14035_/A1 _09664_/B _10370_/X _14035_/B1 _19842_/Q vssd1 vssd1 vccd1 vccd1
+ _14067_/C sky130_fd_sc_hd__o32a_1
Xfanout683 _13863_/B vssd1 vssd1 vccd1 vccd1 _14527_/A2 sky130_fd_sc_hd__buf_4
XFILLER_19_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout694 _14099_/B vssd1 vssd1 vccd1 vccd1 _14107_/B sky130_fd_sc_hd__buf_4
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15720_ _20933_/Q _15995_/A2 _15719_/X vssd1 vssd1 vccd1 vccd1 _15720_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12932_ _19253_/Q _12964_/A2 _16945_/B _20001_/Q vssd1 vssd1 vccd1 vccd1 _16711_/A
+ sky130_fd_sc_hd__a22o_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _19543_/Q _16007_/A _15650_/X _16171_/A vssd1 vssd1 vccd1 vccd1 _19543_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_234_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12863_ _12851_/Y _13332_/B _12853_/B vssd1 vssd1 vccd1 vccd1 _13321_/B sky130_fd_sc_hd__o21a_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14602_ _19366_/Q _17852_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19366_/D sky130_fd_sc_hd__mux2_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11814_ _11903_/A1 _20713_/Q _11891_/B _11813_/X vssd1 vssd1 vccd1 vccd1 _11814_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_27_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18370_ _20840_/Q _18385_/B _18369_/Y _18740_/A vssd1 vssd1 vccd1 vccd1 _20840_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15582_/A _16028_/C vssd1 vssd1 vccd1 vccd1 _15582_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12794_ _12714_/X _12726_/C _12726_/A vssd1 vssd1 vccd1 vccd1 _12794_/X sky130_fd_sc_hd__a21o_1
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _20212_/Q _17321_/A2 _17305_/C _17320_/X _17330_/C1 vssd1 vssd1 vccd1 vccd1
+ _17321_/X sky130_fd_sc_hd__a221o_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _19303_/Q _17051_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19303_/D sky130_fd_sc_hd__mux2_1
XFILLER_199_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11795_/A _11795_/B _13416_/A _13415_/A vssd1 vssd1 vccd1 vccd1 _11745_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _20189_/Q _17235_/Y _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17252_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14464_ _18694_/A _14464_/B vssd1 vssd1 vccd1 vccd1 _19256_/D sky130_fd_sc_hd__and2_1
XFILLER_202_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11676_ _19384_/Q _20675_/Q _11676_/S vssd1 vssd1 vccd1 vccd1 _11676_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _19626_/Q _17855_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19626_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13415_ _13415_/A _13415_/B vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__xnor2_4
X_17183_ _20149_/Q _17708_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20149_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10627_ _10629_/A _10625_/X _10626_/X _12850_/A1 vssd1 vssd1 vccd1 vccd1 _10627_/X
+ sky130_fd_sc_hd__o211a_1
X_14395_ _14392_/B _14394_/Y _14417_/S vssd1 vssd1 vccd1 vccd1 _14395_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16134_ _16708_/B _16196_/S vssd1 vssd1 vccd1 vccd1 _16134_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13346_ _13346_/A _13346_/B _13346_/C vssd1 vssd1 vccd1 vccd1 _13347_/B sky130_fd_sc_hd__nand3_1
X_10558_ _11236_/B _10558_/B vssd1 vssd1 vccd1 vccd1 _10558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16065_ _19558_/Q _15814_/A _16064_/X _16187_/A vssd1 vssd1 vccd1 vccd1 _19558_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ _13586_/B _13586_/C _12795_/X vssd1 vssd1 vccd1 vccd1 _13600_/B sky130_fd_sc_hd__a21oi_2
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10489_ _11281_/A _20599_/Q _11268_/C vssd1 vssd1 vccd1 vccd1 _10489_/X sky130_fd_sc_hd__and3_1
X_15016_ _15016_/A vssd1 vssd1 vccd1 vccd1 _15016_/Y sky130_fd_sc_hd__inv_2
X_12228_ _12226_/X _12227_/X _12383_/A vssd1 vssd1 vccd1 vccd1 _12228_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19824_ _20669_/CLK _19824_/D vssd1 vssd1 vccd1 vccd1 _19824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12159_ _11367_/A _11726_/S _12158_/Y vssd1 vssd1 vccd1 vccd1 _12284_/A sky130_fd_sc_hd__o21a_2
XFILLER_284_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19755_ _20742_/CLK _19755_/D vssd1 vssd1 vccd1 vccd1 _19755_/Q sky130_fd_sc_hd__dfxtp_1
X_16967_ input61/X input96/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16967_/X sky130_fd_sc_hd__mux2_8
XFILLER_256_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18706_ _18985_/A _18706_/B vssd1 vssd1 vccd1 vccd1 _20953_/D sky130_fd_sc_hd__and2_1
X_15918_ _16002_/A1 _15904_/Y _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15918_/X sky130_fd_sc_hd__a21o_1
XFILLER_265_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19686_ _20481_/CLK _19686_/D vssd1 vssd1 vccd1 vccd1 _19686_/Q sky130_fd_sc_hd__dfxtp_1
X_16898_ _19233_/Q _16980_/A2 _16980_/B1 _19102_/Q _16897_/X vssd1 vssd1 vccd1 vccd1
+ _16898_/X sky130_fd_sc_hd__o221a_1
XFILLER_253_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15849_ _15849_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15849_/Y sky130_fd_sc_hd__nand2_1
X_18637_ _18520_/X _18688_/A2 _18635_/Y _18636_/Y vssd1 vssd1 vccd1 vccd1 _18638_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18568_ _18783_/A _18568_/B vssd1 vssd1 vccd1 vccd1 _20914_/D sky130_fd_sc_hd__nor2_1
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17519_ _17525_/A1 _17518_/Y _17430_/A vssd1 vssd1 vccd1 vccd1 _20294_/D sky130_fd_sc_hd__a21oi_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18499_ _18612_/B _18499_/B vssd1 vssd1 vccd1 vccd1 _18499_/X sky130_fd_sc_hd__or2_1
XFILLER_177_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20530_ _20662_/CLK _20530_/D vssd1 vssd1 vccd1 vccd1 _20530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20461_ _21047_/A _20461_/D vssd1 vssd1 vccd1 vccd1 _20461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20392_ _20580_/CLK _20392_/D vssd1 vssd1 vccd1 vccd1 _20392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21013_ _21013_/CLK _21013_/D vssd1 vssd1 vccd1 vccd1 _21013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput286 _13828_/X vssd1 vssd1 vccd1 vccd1 addr0[1] sky130_fd_sc_hd__buf_4
XFILLER_59_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput297 _13784_/X vssd1 vssd1 vccd1 vccd1 addr1[3] sky130_fd_sc_hd__buf_4
XFILLER_88_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09706_ _09698_/X _09699_/X _11980_/S vssd1 vssd1 vccd1 vccd1 _09706_/X sky130_fd_sc_hd__mux2_1
XFILLER_244_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09637_ _09612_/X _09636_/B _09610_/C vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__a21oi_4
XFILLER_71_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09568_ _12577_/A _15442_/A vssd1 vssd1 vccd1 vccd1 _11281_/B sky130_fd_sc_hd__or2_4
XFILLER_70_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09499_ _19214_/Q vssd1 vssd1 vccd1 vccd1 _13967_/S sky130_fd_sc_hd__inv_2
XFILLER_169_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11530_ _12144_/C1 _11519_/X _11522_/X _11529_/X _12152_/A1 vssd1 vssd1 vccd1 vccd1
+ _11530_/X sky130_fd_sc_hd__a311o_1
XFILLER_11_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20728_ _20760_/CLK _20728_/D vssd1 vssd1 vccd1 vccd1 _20728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11461_ _11459_/X _11460_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _11461_/X sky130_fd_sc_hd__mux2_1
X_20659_ _20659_/CLK _20659_/D vssd1 vssd1 vccd1 vccd1 _20659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ _20938_/Q _13363_/B _18683_/B vssd1 vssd1 vccd1 vccd1 _13200_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10412_ _19809_/Q _10603_/B _10410_/X _12085_/B2 _10411_/X vssd1 vssd1 vccd1 vccd1
+ _10412_/X sky130_fd_sc_hd__o221a_1
X_11392_ _19374_/Q _11392_/A2 _11390_/X _09738_/A _11391_/X vssd1 vssd1 vccd1 vccd1
+ _11392_/X sky130_fd_sc_hd__o221a_1
X_14180_ _19499_/Q _14171_/B _14179_/X vssd1 vssd1 vccd1 vccd1 _14181_/B sky130_fd_sc_hd__a21oi_4
XFILLER_164_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _13363_/B _13129_/Y _13130_/X _14110_/B vssd1 vssd1 vccd1 vccd1 _13131_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_164_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10343_ _09507_/A _10342_/X _10341_/X vssd1 vssd1 vccd1 vccd1 _10343_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13062_ _13056_/Y _13518_/A _13517_/B vssd1 vssd1 vccd1 vccd1 _13062_/Y sky130_fd_sc_hd__o21ai_2
X_10274_ _19509_/Q _15593_/A _11726_/S vssd1 vssd1 vccd1 vccd1 _11416_/B sky130_fd_sc_hd__mux2_4
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12013_ _19892_/Q _19793_/Q _12013_/S vssd1 vssd1 vccd1 vccd1 _12013_/X sky130_fd_sc_hd__mux2_1
Xfanout1401 _12081_/S0 vssd1 vssd1 vccd1 vccd1 _10092_/S sky130_fd_sc_hd__buf_8
X_17870_ _20643_/Q _17870_/A1 _17878_/S vssd1 vssd1 vccd1 vccd1 _20643_/D sky130_fd_sc_hd__mux2_1
XFILLER_239_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1412 fanout1430/X vssd1 vssd1 vccd1 vccd1 _10174_/S sky130_fd_sc_hd__buf_4
Xfanout1423 _11393_/S0 vssd1 vssd1 vccd1 vccd1 _12346_/S sky130_fd_sc_hd__buf_6
XFILLER_239_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1434 _11852_/B2 vssd1 vssd1 vccd1 vccd1 _12183_/C1 sky130_fd_sc_hd__buf_6
XFILLER_79_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1445 _11846_/C vssd1 vssd1 vccd1 vccd1 _11851_/C sky130_fd_sc_hd__buf_6
XFILLER_94_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16821_ _16932_/B1 _16818_/X _16820_/X _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16822_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1456 _09734_/Y vssd1 vssd1 vccd1 vccd1 _12411_/C sky130_fd_sc_hd__clkbuf_4
Xfanout1467 _12011_/S vssd1 vssd1 vccd1 vccd1 _11849_/S sky130_fd_sc_hd__buf_6
XFILLER_94_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1478 _12186_/S vssd1 vssd1 vccd1 vccd1 _12189_/A sky130_fd_sc_hd__buf_6
XFILLER_281_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout491 _17919_/X vssd1 vssd1 vccd1 vccd1 _17934_/S sky130_fd_sc_hd__buf_12
Xfanout1489 _09839_/A vssd1 vssd1 vccd1 vccd1 _12192_/A1 sky130_fd_sc_hd__buf_6
XFILLER_281_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16752_ _16822_/A _16752_/B vssd1 vssd1 vccd1 vccd1 _16752_/Y sky130_fd_sc_hd__nor2_1
X_19540_ _19541_/CLK _19540_/D vssd1 vssd1 vccd1 vccd1 _19540_/Q sky130_fd_sc_hd__dfxtp_4
X_13964_ _19187_/Q _14055_/C _14042_/S vssd1 vssd1 vccd1 vccd1 _13964_/X sky130_fd_sc_hd__mux2_1
XFILLER_247_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _15977_/A1 _12835_/Y _15702_/X _15703_/B2 vssd1 vssd1 vccd1 vccd1 _15705_/A
+ sky130_fd_sc_hd__o22a_1
X_12915_ _16037_/A _12486_/B _12484_/X _12914_/Y vssd1 vssd1 vccd1 vccd1 _12915_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16683_ _19938_/Q _17861_/A1 _16701_/S vssd1 vssd1 vccd1 vccd1 _19938_/D sky130_fd_sc_hd__mux2_1
X_19471_ _20698_/CLK _19471_/D vssd1 vssd1 vccd1 vccd1 _19471_/Q sky130_fd_sc_hd__dfxtp_1
X_13895_ _19113_/Q _19050_/S _13896_/B1 _19179_/Q _14458_/A vssd1 vssd1 vccd1 vccd1
+ _19113_/D sky130_fd_sc_hd__o221a_1
XFILLER_62_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18422_ _18422_/A _18422_/B vssd1 vssd1 vccd1 vccd1 _20865_/D sky130_fd_sc_hd__and2_1
XFILLER_222_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15634_ _20866_/Q _16042_/A2 fanout819/X vssd1 vssd1 vccd1 vccd1 _15634_/X sky130_fd_sc_hd__o21ba_1
XFILLER_62_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _12846_/A vssd1 vssd1 vccd1 vccd1 _12846_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _18508_/B _18363_/B vssd1 vssd1 vccd1 vccd1 _18353_/Y sky130_fd_sc_hd__nand2_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _21026_/Q _20994_/Q _15993_/S vssd1 vssd1 vccd1 vccd1 _15565_/X sky130_fd_sc_hd__mux2_1
XFILLER_261_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ _19502_/Q _12786_/B vssd1 vssd1 vccd1 vccd1 _12777_/X sky130_fd_sc_hd__and2_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _20207_/Q _17328_/A2 _17303_/X _17974_/B1 vssd1 vssd1 vccd1 vccd1 _20207_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _19294_/Q _17111_/A1 _14516_/S vssd1 vssd1 vccd1 vccd1 _19294_/D sky130_fd_sc_hd__mux2_1
X_18284_ _18299_/A1 _14373_/B _18283_/Y vssd1 vssd1 vccd1 vccd1 _18541_/B sky130_fd_sc_hd__o21ai_4
X_11728_ _13166_/B vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__clkinv_2
XFILLER_222_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15496_ _15611_/S _15214_/B _15610_/A1 vssd1 vssd1 vccd1 vccd1 _15496_/X sky130_fd_sc_hd__a21o_1
XFILLER_187_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ _17235_/A _17235_/B vssd1 vssd1 vccd1 vccd1 _17235_/Y sky130_fd_sc_hd__nand2_4
XFILLER_30_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14447_ _20219_/Q _19248_/Q _14477_/S vssd1 vssd1 vccd1 vccd1 _14448_/B sky130_fd_sc_hd__mux2_1
XFILLER_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11659_ _10430_/S _20707_/Q _12053_/S _11658_/X vssd1 vssd1 vccd1 vccd1 _11659_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17166_ _20132_/Q _17657_/A1 _17166_/S vssd1 vssd1 vccd1 vccd1 _20132_/D sky130_fd_sc_hd__mux2_1
X_14378_ _13139_/A _14377_/X _13239_/X vssd1 vssd1 vccd1 vccd1 _14379_/C sky130_fd_sc_hd__a21o_1
XFILLER_183_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16117_ _19583_/Q _16127_/A2 _16127_/B1 vssd1 vssd1 vccd1 vccd1 _16117_/X sky130_fd_sc_hd__o21a_1
X_13329_ _20964_/Q _13355_/B _13328_/Y _18593_/A2 vssd1 vssd1 vccd1 vccd1 _13329_/X
+ sky130_fd_sc_hd__a211o_1
X_17097_ _20067_/Q _17097_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20067_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16048_ _19765_/Q _14948_/Y _16047_/X _16048_/C1 vssd1 vssd1 vccd1 vccd1 _16048_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19807_ _20438_/CLK _19807_/D vssd1 vssd1 vccd1 vccd1 _19807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17999_ _20737_/Q _17995_/B _17998_/Y vssd1 vssd1 vccd1 vccd1 _20737_/D sky130_fd_sc_hd__o21a_1
XFILLER_229_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19738_ _20759_/CLK _19738_/D vssd1 vssd1 vccd1 vccd1 _19738_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1990 _19051_/A vssd1 vssd1 vccd1 vccd1 _18048_/A sky130_fd_sc_hd__buf_4
XFILLER_49_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19669_ _20179_/CLK _19669_/D vssd1 vssd1 vccd1 vccd1 _19669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_252_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20513_ _20585_/CLK _20513_/D vssd1 vssd1 vccd1 vccd1 _20513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20444_ _20702_/CLK _20444_/D vssd1 vssd1 vccd1 vccd1 _20444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20375_ _21047_/A _20375_/D vssd1 vssd1 vccd1 vccd1 _20375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_188_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19617_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_117_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21013_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10961_ _10958_/X _10959_/X _10960_/X _12429_/A1 _12430_/S vssd1 vssd1 vccd1 vccd1
+ _10961_/X sky130_fd_sc_hd__a221o_1
XFILLER_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ _12693_/A _12693_/B _12699_/C _12645_/Y _12636_/Y vssd1 vssd1 vccd1 vccd1
+ _12701_/B sky130_fd_sc_hd__o311a_2
XFILLER_232_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ _13680_/A _13684_/B vssd1 vssd1 vccd1 vccd1 _13680_/Y sky130_fd_sc_hd__nand2_4
XFILLER_252_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10892_ _11061_/A _16077_/A vssd1 vssd1 vccd1 vccd1 _10892_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12631_ _12479_/A _12657_/A2 _12682_/B _12630_/Y vssd1 vssd1 vccd1 vccd1 _12631_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15350_ _13568_/A _15185_/B _12579_/D vssd1 vssd1 vccd1 vccd1 _15350_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12562_ _12562_/A vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__inv_6
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ _14301_/A _14301_/B vssd1 vssd1 vccd1 vccd1 _14304_/A sky130_fd_sc_hd__nand2_1
XFILLER_211_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11513_ _11505_/X _11506_/X _11513_/S vssd1 vssd1 vccd1 vccd1 _11513_/X sky130_fd_sc_hd__mux2_1
X_15281_ _15021_/A _15268_/X _15280_/X vssd1 vssd1 vccd1 vccd1 _16774_/B sky130_fd_sc_hd__a21oi_4
XFILLER_200_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12493_ _12493_/A _12493_/B vssd1 vssd1 vccd1 vccd1 _12493_/X sky130_fd_sc_hd__or2_2
XFILLER_12_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17020_ _19998_/Q input207/X _17849_/S vssd1 vssd1 vccd1 vccd1 _19998_/D sky130_fd_sc_hd__mux2_1
XFILLER_138_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14232_ _14232_/A _14232_/B vssd1 vssd1 vccd1 vccd1 _14232_/X sky130_fd_sc_hd__xor2_1
X_11444_ _19815_/Q _19319_/Q _12146_/S vssd1 vssd1 vccd1 vccd1 _11444_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _14158_/B _14162_/Y _14202_/S vssd1 vssd1 vccd1 vccd1 _14163_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11375_ _11371_/X _11374_/X _11375_/S vssd1 vssd1 vccd1 vccd1 _11375_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13114_ _19243_/Q _13114_/B vssd1 vssd1 vccd1 vccd1 _13114_/X sky130_fd_sc_hd__or2_1
X_10326_ _11270_/A2 _10322_/X _10325_/X _09689_/C vssd1 vssd1 vccd1 vccd1 _10326_/X
+ sky130_fd_sc_hd__o211a_1
X_14094_ _19206_/Q _14106_/A2 _14093_/X _14104_/C1 vssd1 vssd1 vccd1 vccd1 _19206_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18971_ _21010_/Q _18971_/B vssd1 vssd1 vccd1 vccd1 _18971_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17922_ _20691_/Q _17922_/A1 _17934_/S vssd1 vssd1 vccd1 vccd1 _20691_/D sky130_fd_sc_hd__mux2_1
X_13045_ _20955_/Q _20889_/Q vssd1 vssd1 vccd1 vccd1 _13590_/A sky130_fd_sc_hd__nor2_1
X_10257_ _10262_/A _20380_/Q _20444_/Q _11042_/B vssd1 vssd1 vccd1 vccd1 _10257_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout1220 _13370_/B vssd1 vssd1 vccd1 vccd1 _13272_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_67_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1231 _12784_/B vssd1 vssd1 vccd1 vccd1 _12682_/B sky130_fd_sc_hd__buf_4
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17853_ _20626_/Q _17887_/A1 _17883_/S vssd1 vssd1 vccd1 vccd1 _20626_/D sky130_fd_sc_hd__mux2_1
XFILLER_239_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10188_ _10937_/A _20670_/Q _11191_/C vssd1 vssd1 vccd1 vccd1 _10188_/X sky130_fd_sc_hd__or3_1
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1242 _17382_/B1 vssd1 vssd1 vccd1 vccd1 _17530_/A2 sky130_fd_sc_hd__buf_4
XFILLER_67_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1253 _17335_/X vssd1 vssd1 vccd1 vccd1 _17371_/A2 sky130_fd_sc_hd__buf_6
Xfanout1264 _09689_/X vssd1 vssd1 vccd1 vccd1 _12075_/C1 sky130_fd_sc_hd__buf_6
XFILLER_266_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16804_ _16869_/A _16804_/B vssd1 vssd1 vccd1 vccd1 _16804_/Y sky130_fd_sc_hd__nand2_1
XFILLER_254_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1286 _09546_/Y vssd1 vssd1 vccd1 vccd1 _15922_/B2 sky130_fd_sc_hd__clkbuf_16
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14996_ _15314_/D _15022_/D vssd1 vssd1 vccd1 vccd1 _14996_/X sky130_fd_sc_hd__or2_4
X_17784_ _20561_/Q _17924_/A1 _17794_/S vssd1 vssd1 vccd1 vccd1 _20561_/D sky130_fd_sc_hd__mux2_1
Xfanout1297 _09540_/X vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__buf_6
XFILLER_219_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19523_ _19523_/CLK _19523_/D vssd1 vssd1 vccd1 vccd1 _19523_/Q sky130_fd_sc_hd__dfxtp_4
X_16735_ _20183_/Q _17219_/B _16717_/X vssd1 vssd1 vccd1 vccd1 _16735_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13947_ _19149_/Q _14522_/A _13906_/X vssd1 vssd1 vccd1 vccd1 _19149_/D sky130_fd_sc_hd__o21ba_1
XFILLER_207_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19454_ _20713_/CLK _19454_/D vssd1 vssd1 vccd1 vccd1 _19454_/Q sky130_fd_sc_hd__dfxtp_1
X_16666_ _19923_/Q _17178_/A1 _16666_/S vssd1 vssd1 vccd1 vccd1 _19923_/D sky130_fd_sc_hd__mux2_1
X_13878_ _19096_/Q _14527_/A2 _13900_/A2 _12510_/C _16195_/A vssd1 vssd1 vccd1 vccd1
+ _19096_/D sky130_fd_sc_hd__o221a_1
X_18405_ _20857_/Q _18195_/Y _18419_/S vssd1 vssd1 vccd1 vccd1 _18406_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15617_ _13426_/A _15982_/C _16056_/B1 vssd1 vssd1 vccd1 vccd1 _15617_/X sky130_fd_sc_hd__a21o_1
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12829_ _12839_/A _12829_/B _12829_/C _12829_/D vssd1 vssd1 vccd1 vccd1 _12866_/A
+ sky130_fd_sc_hd__nor4_2
X_16597_ _16598_/A _16594_/B _16595_/Y input9/X vssd1 vssd1 vccd1 vccd1 _16597_/X
+ sky130_fd_sc_hd__o22a_1
X_19385_ _19956_/CLK _19385_/D vssd1 vssd1 vccd1 vccd1 _19385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18336_ _20823_/Q _18349_/B _18335_/Y _18702_/A vssd1 vssd1 vccd1 vccd1 _20823_/D
+ sky130_fd_sc_hd__o211a_1
X_15548_ _15066_/S _15109_/X _15548_/B1 vssd1 vssd1 vccd1 vccd1 _15548_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_148_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18267_ _18728_/A _18267_/B vssd1 vssd1 vccd1 vccd1 _20807_/D sky130_fd_sc_hd__and2_1
X_15479_ _20925_/Q _15567_/A2 _15478_/X vssd1 vssd1 vccd1 vccd1 _15479_/X sky130_fd_sc_hd__o21a_1
X_17218_ _17219_/A _17219_/B _17219_/C vssd1 vssd1 vccd1 vccd1 _17224_/B sky130_fd_sc_hd__and3_1
XFILLER_129_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18198_ _19535_/Q _18198_/B vssd1 vssd1 vccd1 vccd1 _18198_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17149_ _20117_/Q _17708_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20117_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20160_ _20703_/CLK _20160_/D vssd1 vssd1 vccd1 vccd1 _20160_/Q sky130_fd_sc_hd__dfxtp_1
X_09971_ _19386_/Q _20677_/Q _12149_/S vssd1 vssd1 vccd1 vccd1 _09971_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20091_ _20155_/CLK _20091_/D vssd1 vssd1 vccd1 vccd1 _20091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_210_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20676_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_609 input228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20993_ _21025_/CLK _20993_/D vssd1 vssd1 vccd1 vccd1 _20993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20427_ _20428_/CLK _20427_/D vssd1 vssd1 vccd1 vccd1 _20427_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11160_ _12230_/A1 _20494_/Q _11161_/S _20526_/Q _12318_/A1 vssd1 vssd1 vccd1 vccd1
+ _11160_/X sky130_fd_sc_hd__o221a_1
X_20358_ _20717_/CLK _20358_/D vssd1 vssd1 vccd1 vccd1 _20358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10111_ _10112_/A _11412_/B vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__or2_4
XFILLER_134_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11091_ _12395_/S _11090_/X _11089_/X _12399_/A1 vssd1 vssd1 vccd1 vccd1 _11091_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20289_ _21004_/CLK _20289_/D vssd1 vssd1 vccd1 vccd1 _20289_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _10037_/Y _10041_/Y _09669_/X vssd1 vssd1 vccd1 vccd1 _10042_/X sky130_fd_sc_hd__a21o_1
XFILLER_276_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xsplit8 split8/A vssd1 vssd1 vccd1 vccd1 split8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14850_ _11416_/B _11735_/B _15983_/A vssd1 vssd1 vccd1 vccd1 _14850_/X sky130_fd_sc_hd__mux2_1
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _13802_/A1 _13678_/Y _13805_/B1 input216/X vssd1 vssd1 vccd1 vccd1 _13801_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14781_ _19515_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14781_/X sky130_fd_sc_hd__or2_1
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11993_ _20049_/Q _19924_/Q _11994_/S vssd1 vssd1 vccd1 vccd1 _11993_/X sky130_fd_sc_hd__mux2_1
X_16520_ _19827_/Q _17915_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19827_/D sky130_fd_sc_hd__mux2_1
XFILLER_217_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13732_ _13776_/B1 _13772_/B _13731_/X vssd1 vssd1 vccd1 vccd1 _13733_/B sky130_fd_sc_hd__a21oi_4
X_10944_ _20401_/Q _20337_/Q _20629_/Q _20593_/Q _11203_/S _11026_/C vssd1 vssd1 vccd1
+ vccd1 _10944_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16451_ _16451_/A _16451_/B _16451_/C vssd1 vssd1 vccd1 vccd1 _19764_/D sky130_fd_sc_hd__nor3_1
XFILLER_188_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13663_ _13663_/A _13663_/B _13735_/B vssd1 vssd1 vccd1 vccd1 _13663_/X sky130_fd_sc_hd__and3_4
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10875_ _11391_/A _19339_/Q _20694_/Q _12344_/S _11212_/S vssd1 vssd1 vccd1 vccd1
+ _10875_/X sky130_fd_sc_hd__a221o_1
XFILLER_204_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15402_ _15402_/A _15402_/B vssd1 vssd1 vccd1 vccd1 _15402_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19170_ _20426_/CLK _19170_/D vssd1 vssd1 vccd1 vccd1 _19170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _19523_/Q _19522_/Q _12901_/B vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__and3_1
X_16382_ _16386_/C _16382_/B vssd1 vssd1 vccd1 vccd1 _19738_/D sky130_fd_sc_hd__nor2_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13594_ _14524_/A1 _19224_/Q _13593_/X vssd1 vssd1 vccd1 vccd1 _13921_/A sky130_fd_sc_hd__a21oi_2
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18121_ _20782_/Q _18122_/C _18120_/Y vssd1 vssd1 vccd1 vccd1 _20782_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_85_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _20721_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15333_ _20729_/Q _15445_/A2 _15445_/B1 _20761_/Q vssd1 vssd1 vccd1 vccd1 _15333_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12545_ _20872_/Q _12549_/B _12545_/C vssd1 vssd1 vccd1 vccd1 _12551_/D sky130_fd_sc_hd__and3_1
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20568_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18052_ _20756_/Q _18053_/C _20757_/Q vssd1 vssd1 vccd1 vccd1 _18054_/B sky130_fd_sc_hd__a21oi_1
X_15264_ _15264_/A _15264_/B vssd1 vssd1 vccd1 vccd1 _15264_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12476_ _12454_/Y _16030_/D1 _12472_/X _12475_/X vssd1 vssd1 vccd1 vccd1 _12476_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17003_ _19246_/Q _17003_/B vssd1 vssd1 vccd1 vccd1 _17003_/X sky130_fd_sc_hd__or2_4
XFILLER_8_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14215_ _19224_/Q _14256_/A2 _14214_/X _14758_/C1 vssd1 vssd1 vccd1 vccd1 _19224_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_5 _15274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _20542_/Q _12139_/S vssd1 vssd1 vccd1 vccd1 _11427_/X sky130_fd_sc_hd__or2_1
X_15195_ _20949_/Q _15568_/A2 _15568_/B1 _20821_/Q _15194_/X vssd1 vssd1 vccd1 vccd1
+ _15195_/X sky130_fd_sc_hd__a221o_4
XFILLER_153_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _20269_/Q _14117_/A _14216_/B1 input240/X vssd1 vssd1 vccd1 vccd1 _14148_/B
+ sky130_fd_sc_hd__a22o_2
X_11358_ _19806_/Q _19310_/Q _11358_/S vssd1 vssd1 vccd1 vccd1 _11358_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10309_ _12513_/C _10297_/X _10301_/X _09621_/A vssd1 vssd1 vccd1 vccd1 _10309_/X
+ sky130_fd_sc_hd__o211a_1
X_14077_ _14099_/A _14099_/B _14077_/C vssd1 vssd1 vccd1 vccd1 _14077_/X sky130_fd_sc_hd__or3_1
XFILLER_140_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18954_ _19112_/Q _18954_/A2 _18967_/B1 _13183_/Y vssd1 vssd1 vccd1 vccd1 _18955_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11289_ _11026_/A _20493_/Q _11292_/S0 _20525_/Q vssd1 vssd1 vccd1 vccd1 _11289_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_141_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17905_ _20676_/Q _17905_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20676_/D sky130_fd_sc_hd__mux2_1
X_13028_ _20965_/Q _20899_/Q vssd1 vssd1 vccd1 vccd1 _13303_/B sky130_fd_sc_hd__nand2_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18885_ _19102_/Q _18954_/A2 _18967_/B1 _13427_/A vssd1 vssd1 vccd1 vccd1 _18886_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1050 _17189_/A1 vssd1 vssd1 vccd1 vccd1 _17923_/A1 sky130_fd_sc_hd__buf_4
XFILLER_267_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1061 _17892_/A1 vssd1 vssd1 vccd1 vccd1 _17683_/A1 sky130_fd_sc_hd__buf_4
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1072 _17919_/B vssd1 vssd1 vccd1 vccd1 _17676_/B sky130_fd_sc_hd__clkbuf_4
X_17836_ _20611_/Q _17874_/A1 _17840_/S vssd1 vssd1 vccd1 vccd1 _20611_/D sky130_fd_sc_hd__mux2_1
XFILLER_282_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1083 _12576_/Y vssd1 vssd1 vccd1 vccd1 _15326_/A sky130_fd_sc_hd__buf_6
Xfanout1094 _12210_/X vssd1 vssd1 vccd1 vccd1 _17706_/A1 sky130_fd_sc_hd__buf_6
XFILLER_266_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17767_ _20546_/Q _17835_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20546_/D sky130_fd_sc_hd__mux2_1
X_14979_ _14983_/A _14979_/B vssd1 vssd1 vccd1 vccd1 _14979_/Y sky130_fd_sc_hd__nor2_1
XFILLER_207_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19506_ _19506_/CLK _19506_/D vssd1 vssd1 vccd1 vccd1 _19506_/Q sky130_fd_sc_hd__dfxtp_4
X_16718_ _12952_/X _16717_/X _12930_/B vssd1 vssd1 vccd1 vccd1 _16718_/X sky130_fd_sc_hd__a21bo_4
XFILLER_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17698_ _20482_/Q _17801_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20482_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19437_ _20468_/CLK _19437_/D vssd1 vssd1 vccd1 vccd1 _19437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16649_ _19906_/Q _17686_/A1 _16666_/S vssd1 vssd1 vccd1 vccd1 _19906_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19368_ _20659_/CLK _19368_/D vssd1 vssd1 vccd1 vccd1 _19368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18319_ _18319_/A _18389_/B _18389_/C vssd1 vssd1 vccd1 vccd1 _18981_/B sky130_fd_sc_hd__or3_4
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19299_ _19697_/CLK _19299_/D vssd1 vssd1 vccd1 vccd1 _19299_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_148_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20212_ _20766_/CLK _20212_/D vssd1 vssd1 vccd1 vccd1 _20212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20143_ _20482_/CLK _20143_/D vssd1 vssd1 vccd1 vccd1 _20143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _11903_/A1 _20709_/Q _11891_/B _09953_/X vssd1 vssd1 vccd1 vccd1 _09954_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_104_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20074_ _20717_/CLK _20074_/D vssd1 vssd1 vccd1 vccd1 _20074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09885_ _09875_/X _09877_/X _09884_/X _11904_/S _12137_/A1 vssd1 vssd1 vccd1 vccd1
+ _09885_/X sky130_fd_sc_hd__o221a_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_406 _16985_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_261_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_417 _18589_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_428 _16037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20976_ _21000_/CLK _20976_/D vssd1 vssd1 vccd1 vccd1 _20976_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_439 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10660_ _20372_/Q _20436_/Q _12381_/S vssd1 vssd1 vccd1 vccd1 _10660_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10591_ _12051_/A1 _19906_/Q _11994_/S _20031_/Q _12056_/S vssd1 vssd1 vccd1 vccd1
+ _10591_/X sky130_fd_sc_hd__o221a_1
XFILLER_167_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ _11726_/S _11367_/B _12328_/Y _12329_/Y vssd1 vssd1 vccd1 vccd1 _12440_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12261_ _12259_/X _12260_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _12261_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14000_ _19199_/Q _14079_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _14000_/X sky130_fd_sc_hd__mux2_1
X_11212_ _11210_/X _11211_/X _11212_/S vssd1 vssd1 vccd1 vccd1 _11212_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12192_ _12192_/A1 _12179_/X _12183_/X _12191_/X _10409_/A vssd1 vssd1 vccd1 vccd1
+ _12192_/X sky130_fd_sc_hd__o311a_1
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11143_ _19560_/Q _14524_/B1 _19527_/Q vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_268_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_132_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20982_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11074_ _20120_/Q _20088_/Q _11074_/S vssd1 vssd1 vccd1 vccd1 _11074_/X sky130_fd_sc_hd__mux2_1
X_15951_ _12519_/A _15978_/A2 _15950_/Y vssd1 vssd1 vccd1 vccd1 _15952_/B sky130_fd_sc_hd__a21oi_1
XFILLER_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput120 dout1[21] vssd1 vssd1 vccd1 vccd1 input120/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput131 dout1[31] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput142 dout1[41] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__buf_2
X_10025_ input110/X input145/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10025_/X sky130_fd_sc_hd__mux2_8
X_14902_ _18136_/B _16720_/D vssd1 vssd1 vccd1 vccd1 _14902_/X sky130_fd_sc_hd__or2_1
Xinput153 dout1[51] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__clkbuf_2
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18670_ _20941_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18670_/Y sky130_fd_sc_hd__nand2_1
X_15882_ _15882_/A1 _15871_/X _15872_/X _15881_/X vssd1 vssd1 vccd1 vccd1 _15882_/X
+ sky130_fd_sc_hd__a22o_4
Xinput164 dout1[61] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_hd__clkbuf_2
XFILLER_264_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 irq[13] vssd1 vssd1 vccd1 vccd1 _12541_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_263_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 irq[9] vssd1 vssd1 vccd1 vccd1 _12544_/C sky130_fd_sc_hd__clkbuf_2
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _20377_/Q _17689_/A1 _17635_/S vssd1 vssd1 vccd1 vccd1 _20377_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput197 localMemory_wb_adr_i[16] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__clkbuf_2
X_14833_ _11051_/Y _12198_/B _14837_/S vssd1 vssd1 vccd1 vccd1 _14833_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _19129_/Q _14764_/A2 _14763_/X _18352_/C1 vssd1 vssd1 vccd1 vccd1 _19506_/D
+ sky130_fd_sc_hd__o211a_1
X_17552_ _20312_/Q _17931_/A1 _17567_/S vssd1 vssd1 vccd1 vccd1 _20312_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _11977_/A1 _11983_/A1 _19489_/Q _12129_/S vssd1 vssd1 vccd1 vccd1 _11976_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_251_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13715_ _13716_/B vssd1 vssd1 vccd1 vccd1 _13715_/Y sky130_fd_sc_hd__inv_2
X_16503_ _19810_/Q _17096_/A1 _16517_/S vssd1 vssd1 vccd1 vccd1 _19810_/D sky130_fd_sc_hd__mux2_1
X_17483_ _17487_/A1 _17482_/Y _18704_/A vssd1 vssd1 vccd1 vccd1 _20276_/D sky130_fd_sc_hd__a21oi_1
X_10927_ _12311_/A1 _10923_/X _10926_/X _09689_/A _10919_/X vssd1 vssd1 vccd1 vccd1
+ _10928_/C sky130_fd_sc_hd__o311a_1
XFILLER_147_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14695_ _19454_/Q _17944_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19454_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19222_ _19223_/CLK _19222_/D vssd1 vssd1 vccd1 vccd1 _19222_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13646_ _13657_/A _13646_/B vssd1 vssd1 vccd1 vccd1 _13676_/B sky130_fd_sc_hd__nor2_8
X_16434_ _19757_/Q _19758_/Q _16434_/C vssd1 vssd1 vccd1 vccd1 _16437_/B sky130_fd_sc_hd__and3_1
X_10858_ _12332_/A _20662_/Q _12337_/C vssd1 vssd1 vccd1 vccd1 _10858_/X sky130_fd_sc_hd__or3_1
XFILLER_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ _19574_/CLK _19153_/D vssd1 vssd1 vccd1 vccd1 _19153_/Q sky130_fd_sc_hd__dfxtp_4
X_16365_ _19732_/Q _16364_/B _18396_/A vssd1 vssd1 vccd1 vccd1 _16366_/B sky130_fd_sc_hd__o21ai_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _13047_/X _13048_/Y _13066_/X vssd1 vssd1 vccd1 vccd1 _13577_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _10786_/X _10787_/X _10788_/X _12420_/B1 _12265_/A vssd1 vssd1 vccd1 vccd1
+ _10789_/X sky130_fd_sc_hd__a221o_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15316_ _20792_/Q _14975_/Y _14978_/B _15021_/B _15315_/X vssd1 vssd1 vccd1 vccd1
+ _15316_/X sky130_fd_sc_hd__a221o_1
X_18104_ _18104_/A _18109_/C vssd1 vssd1 vccd1 vccd1 _18104_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12528_ _20914_/Q _18462_/A _13107_/B _18763_/A1 vssd1 vssd1 vccd1 vccd1 _12528_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_158_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16296_ _16300_/C _16296_/B vssd1 vssd1 vccd1 vccd1 _19706_/D sky130_fd_sc_hd__nor2_1
XFILLER_258_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19084_ _20410_/CLK _19084_/D vssd1 vssd1 vccd1 vccd1 _19084_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18035_ _20750_/Q _18036_/C _18034_/Y vssd1 vssd1 vccd1 vccd1 _20750_/D sky130_fd_sc_hd__o21a_1
X_15247_ _15348_/B2 _12680_/Y _13524_/A _12578_/A _10935_/B vssd1 vssd1 vccd1 vccd1
+ _15248_/C sky130_fd_sc_hd__o221a_1
XFILLER_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _12565_/B _12471_/B vssd1 vssd1 vccd1 vccd1 _12459_/Y sky130_fd_sc_hd__nand2_1
XFILLER_274_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15178_ _11053_/Y _12471_/X _12468_/X vssd1 vssd1 vccd1 vccd1 _15178_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14129_ _19495_/Q _14130_/B vssd1 vssd1 vccd1 vccd1 _14129_/X sky130_fd_sc_hd__and2_1
X_19986_ _19992_/CLK _19986_/D vssd1 vssd1 vccd1 vccd1 _19986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18937_ _21005_/Q _18937_/B vssd1 vssd1 vccd1 vccd1 _18937_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09670_ _19695_/Q _19657_/Q vssd1 vssd1 vccd1 vccd1 _09670_/Y sky130_fd_sc_hd__nand2_4
X_18868_ _20995_/Q _18937_/B vssd1 vssd1 vccd1 vccd1 _18868_/Y sky130_fd_sc_hd__nand2_1
XFILLER_267_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17819_ _20594_/Q _17857_/A1 _17844_/S vssd1 vssd1 vccd1 vccd1 _20594_/D sky130_fd_sc_hd__mux2_1
XFILLER_227_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18799_ _20985_/Q _18819_/B vssd1 vssd1 vccd1 vccd1 _18799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20830_ _20959_/CLK _20830_/D vssd1 vssd1 vccd1 vccd1 _20830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20761_ _20763_/CLK _20761_/D vssd1 vssd1 vccd1 vccd1 _20761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20692_ _20692_/CLK _20692_/D vssd1 vssd1 vccd1 vccd1 _20692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1808 _15103_/A1 vssd1 vssd1 vccd1 vccd1 _10284_/A sky130_fd_sc_hd__buf_4
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout810 _12592_/C vssd1 vssd1 vccd1 vccd1 _18864_/B1 sky130_fd_sc_hd__buf_2
Xfanout1819 _19178_/Q vssd1 vssd1 vccd1 vccd1 _11367_/A sky130_fd_sc_hd__buf_12
Xfanout821 _15323_/B vssd1 vssd1 vccd1 vccd1 _15994_/B1 sky130_fd_sc_hd__clkbuf_8
X_20126_ _20559_/CLK _20126_/D vssd1 vssd1 vccd1 vccd1 _20126_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout832 _18981_/X vssd1 vssd1 vccd1 vccd1 _18982_/B sky130_fd_sc_hd__buf_8
X_09937_ _19515_/Q _15768_/A _11649_/S vssd1 vssd1 vccd1 vccd1 _10016_/B sky130_fd_sc_hd__mux2_8
XFILLER_131_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout843 _18387_/B vssd1 vssd1 vccd1 vccd1 _18375_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout854 _15998_/A2 vssd1 vssd1 vccd1 vccd1 _15941_/A2 sky130_fd_sc_hd__buf_6
Xfanout865 _14963_/Y vssd1 vssd1 vccd1 vccd1 _15323_/A sky130_fd_sc_hd__buf_8
Xfanout876 _15604_/A2 vssd1 vssd1 vccd1 vccd1 _15453_/A2 sky130_fd_sc_hd__clkbuf_8
X_20057_ _20379_/CLK _20057_/D vssd1 vssd1 vccd1 vccd1 _20057_/Q sky130_fd_sc_hd__dfxtp_1
X_09868_ _19580_/Q _09867_/X _11229_/S vssd1 vssd1 vccd1 vccd1 _10119_/A sky130_fd_sc_hd__mux2_2
Xfanout887 _11018_/Y vssd1 vssd1 vccd1 vccd1 _15407_/S sky130_fd_sc_hd__buf_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout898 _16718_/X vssd1 vssd1 vccd1 vccd1 _17008_/A1 sky130_fd_sc_hd__buf_6
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _20355_/Q _12043_/B vssd1 vssd1 vccd1 vccd1 _09799_/X sky130_fd_sc_hd__or2_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 _19838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ _20421_/Q _12148_/S _11808_/X _12150_/S vssd1 vssd1 vccd1 vccd1 _11830_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_225 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_236 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11761_ _11761_/A _11761_/B _11745_/X vssd1 vssd1 vccd1 vccd1 _15789_/B sky130_fd_sc_hd__or3b_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20959_ _20959_/CLK _20959_/D vssd1 vssd1 vccd1 vccd1 _20959_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13500_ _20917_/Q _13602_/A1 _12525_/Y _13499_/Y _14110_/A vssd1 vssd1 vccd1 vccd1
+ _13500_/X sky130_fd_sc_hd__a221o_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _11375_/S _10711_/X _10708_/X _12431_/A1 vssd1 vssd1 vccd1 vccd1 _10713_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14480_ _18746_/A _14480_/B vssd1 vssd1 vccd1 vccd1 _19264_/D sky130_fd_sc_hd__and2_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _19168_/Q _11649_/S _11691_/Y vssd1 vssd1 vccd1 vccd1 _11729_/A sky130_fd_sc_hd__o21a_1
XFILLER_241_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _13431_/A _13431_/B vssd1 vssd1 vccd1 vccd1 _15949_/B sky130_fd_sc_hd__xnor2_4
XFILLER_186_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10643_ _13611_/A _11766_/B _11764_/B vssd1 vssd1 vccd1 vccd1 _10643_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16150_ _16804_/B _16178_/S vssd1 vssd1 vccd1 vccd1 _16150_/Y sky130_fd_sc_hd__nand2_1
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13362_ _13362_/A _13362_/B _13362_/C vssd1 vssd1 vccd1 vccd1 _13362_/X sky130_fd_sc_hd__and3_1
XFILLER_167_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10574_ _10057_/S _19439_/Q _11676_/S _10572_/X _10573_/X vssd1 vssd1 vccd1 vccd1
+ _10574_/X sky130_fd_sc_hd__a311o_1
XFILLER_167_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15101_ _12578_/B _12493_/B _15100_/Y _10935_/B vssd1 vssd1 vccd1 vccd1 _15101_/X
+ sky130_fd_sc_hd__o211a_1
X_12313_ _20656_/Q _20620_/Q _12313_/S vssd1 vssd1 vccd1 vccd1 _12313_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16081_ _16081_/A _16081_/B vssd1 vssd1 vccd1 vccd1 _16081_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13293_ _13607_/B _13290_/X _13291_/Y _13292_/Y _18612_/B vssd1 vssd1 vccd1 vccd1
+ _13293_/X sky130_fd_sc_hd__o311a_1
X_15032_ _12455_/Y _15520_/B2 _15150_/C1 vssd1 vssd1 vccd1 vccd1 _15032_/Y sky130_fd_sc_hd__a21oi_1
X_12244_ _12229_/X _12243_/X _12401_/A1 vssd1 vssd1 vccd1 vccd1 _12244_/X sky130_fd_sc_hd__a21o_2
X_19840_ _20742_/CLK _19840_/D vssd1 vssd1 vccd1 vccd1 _19840_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_269_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12175_ _12173_/X _12174_/X _12189_/A vssd1 vssd1 vccd1 vccd1 _12175_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11126_ _19664_/Q _11126_/B vssd1 vssd1 vccd1 vccd1 _11126_/X sky130_fd_sc_hd__or2_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19771_ _20630_/CLK _19771_/D vssd1 vssd1 vccd1 vccd1 _19771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16983_ input63/X input99/X _17009_/S vssd1 vssd1 vccd1 vccd1 _16983_/X sky130_fd_sc_hd__mux2_8
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18722_ _18724_/A _18722_/B vssd1 vssd1 vccd1 vccd1 _20961_/D sky130_fd_sc_hd__and2_1
XFILLER_277_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11057_ _11234_/A _10465_/Y _11235_/A vssd1 vssd1 vccd1 vccd1 _11057_/X sky130_fd_sc_hd__a21o_1
X_15934_ _20749_/Q _15934_/A2 _15934_/B1 _20781_/Q vssd1 vssd1 vccd1 vccd1 _15934_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10008_ _19418_/Q _20577_/Q _11947_/S vssd1 vssd1 vccd1 vccd1 _10008_/X sky130_fd_sc_hd__mux2_1
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18653_ _18960_/A _18653_/B vssd1 vssd1 vccd1 vccd1 _20936_/D sky130_fd_sc_hd__nor2_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _15526_/B _15848_/X _15864_/X _15976_/B2 vssd1 vssd1 vccd1 vccd1 _15865_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_225_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _20362_/Q _17881_/A1 _17606_/S vssd1 vssd1 vccd1 vccd1 _20362_/D sky130_fd_sc_hd__mux2_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14816_ _14814_/X _14815_/X _15058_/S vssd1 vssd1 vccd1 vccd1 _14816_/X sky130_fd_sc_hd__mux2_1
X_18584_ _20919_/Q _18592_/B vssd1 vssd1 vccd1 vccd1 _18584_/Y sky130_fd_sc_hd__nand2_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _19724_/Q _15961_/A2 _15961_/B1 _19756_/Q vssd1 vssd1 vccd1 vccd1 _15796_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17535_ _20299_/Q _17529_/X _17534_/X vssd1 vssd1 vccd1 vccd1 _20299_/D sky130_fd_sc_hd__o21ba_1
X_14747_ _19498_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14747_/X sky130_fd_sc_hd__or2_1
X_11959_ _11880_/A _11880_/B _11958_/X vssd1 vssd1 vccd1 vccd1 _11960_/B sky130_fd_sc_hd__a21oi_2
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14678_ _19437_/Q _17684_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19437_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17466_ _20268_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17466_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19205_ _20426_/CLK _19205_/D vssd1 vssd1 vccd1 vccd1 _19205_/Q sky130_fd_sc_hd__dfxtp_1
X_16417_ _19751_/Q _16418_/C _19752_/Q vssd1 vssd1 vccd1 vccd1 _16419_/B sky130_fd_sc_hd__a21oi_1
X_13629_ _13478_/B _13230_/X _15898_/A _13765_/A vssd1 vssd1 vccd1 vccd1 _13629_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_177_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17397_ _20247_/Q _17401_/A2 _17396_/X _17434_/A vssd1 vssd1 vccd1 vccd1 _20247_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19136_ _19511_/CLK _19136_/D vssd1 vssd1 vccd1 vccd1 _19136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16348_ _19726_/Q _16348_/B vssd1 vssd1 vccd1 vccd1 _16354_/C sky130_fd_sc_hd__and2_2
XFILLER_121_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19067_ _20412_/Q vssd1 vssd1 vccd1 vccd1 _20412_/D sky130_fd_sc_hd__clkbuf_2
X_16279_ _17952_/A _16279_/B _16279_/C vssd1 vssd1 vccd1 vccd1 _19701_/D sky130_fd_sc_hd__nor3_4
XFILLER_173_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput402 _13795_/X vssd1 vssd1 vccd1 vccd1 din0[4] sky130_fd_sc_hd__buf_4
X_18018_ _20744_/Q _18019_/C _20745_/Q vssd1 vssd1 vccd1 vccd1 _18020_/B sky130_fd_sc_hd__a21oi_1
Xoutput413 _19973_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[12] sky130_fd_sc_hd__buf_4
XFILLER_161_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput424 _19983_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[22] sky130_fd_sc_hd__buf_4
Xoutput435 _19964_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[3] sky130_fd_sc_hd__buf_4
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput446 _20258_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[1] sky130_fd_sc_hd__buf_4
Xoutput457 _19510_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[16] sky130_fd_sc_hd__buf_4
XFILLER_141_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput468 _19520_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[26] sky130_fd_sc_hd__buf_4
Xoutput479 _19501_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[7] sky130_fd_sc_hd__buf_4
XFILLER_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19969_ _20004_/CLK _19969_/D vssd1 vssd1 vccd1 vccd1 _19969_/Q sky130_fd_sc_hd__dfxtp_1
X_09722_ _12151_/A1 _09721_/X _09718_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _09722_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09653_ _09681_/B _09681_/C vssd1 vssd1 vccd1 vccd1 _10203_/A sky130_fd_sc_hd__nand2_1
XFILLER_95_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09584_ _19087_/Q _19086_/Q _09588_/C vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__or3b_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20813_ _21043_/CLK _20813_/D vssd1 vssd1 vccd1 vccd1 _20813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20744_ _21029_/CLK _20744_/D vssd1 vssd1 vccd1 vccd1 _20744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20675_ _20675_/CLK _20675_/D vssd1 vssd1 vccd1 vccd1 _20675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10290_ _11236_/B _10290_/B vssd1 vssd1 vccd1 vccd1 _10290_/Y sky130_fd_sc_hd__nand2_1
XFILLER_191_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1605 _11170_/B1 vssd1 vssd1 vccd1 vccd1 _11250_/S sky130_fd_sc_hd__buf_8
XFILLER_132_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1616 fanout1630/X vssd1 vssd1 vccd1 vccd1 _11988_/S sky130_fd_sc_hd__buf_4
Xfanout1627 fanout1630/X vssd1 vssd1 vccd1 vccd1 _12309_/S sky130_fd_sc_hd__buf_6
XFILLER_144_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1638 _09614_/X vssd1 vssd1 vccd1 vccd1 _12400_/A1 sky130_fd_sc_hd__buf_12
Xfanout640 _16170_/S vssd1 vssd1 vccd1 vccd1 _16190_/S sky130_fd_sc_hd__buf_8
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout651 _16036_/A2 vssd1 vssd1 vccd1 vccd1 _15814_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1649 _12531_/Y vssd1 vssd1 vccd1 vccd1 _18968_/A sky130_fd_sc_hd__buf_8
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20109_ _20712_/CLK _20109_/D vssd1 vssd1 vccd1 vccd1 _20109_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout662 _14397_/B vssd1 vssd1 vccd1 vccd1 _14437_/B sky130_fd_sc_hd__buf_4
X_13980_ _19160_/Q _14004_/A2 _14004_/B1 _13979_/X _16159_/C1 vssd1 vssd1 vccd1 vccd1
+ _19160_/D sky130_fd_sc_hd__o221a_1
XFILLER_282_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout673 _13943_/S vssd1 vssd1 vccd1 vccd1 _13906_/B sky130_fd_sc_hd__buf_4
XFILLER_247_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout684 _13986_/A2 vssd1 vssd1 vccd1 vccd1 _13863_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_281_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout695 _14069_/B vssd1 vssd1 vccd1 vccd1 _14099_/B sky130_fd_sc_hd__buf_4
X_12931_ _19250_/Q _12964_/A2 _16716_/A _19998_/Q vssd1 vssd1 vccd1 vccd1 _14119_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12862_ _13346_/A _13346_/B _12822_/Y _12861_/X vssd1 vssd1 vccd1 vccd1 _12871_/A
+ sky130_fd_sc_hd__a211o_4
X_15650_ _15650_/A _15650_/B _16007_/A vssd1 vssd1 vccd1 vccd1 _15650_/X sky130_fd_sc_hd__or3b_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _17919_/A _17574_/B _14601_/C vssd1 vssd1 vccd1 vccd1 _14601_/X sky130_fd_sc_hd__and3_4
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _11903_/A1 _12120_/A1 _19358_/Q _12129_/S vssd1 vssd1 vccd1 vccd1 _11813_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _15984_/B1 _15580_/X _10366_/A vssd1 vssd1 vccd1 vccd1 _15581_/X sky130_fd_sc_hd__o21a_1
XFILLER_221_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _13281_/A _12748_/B _12749_/C _12791_/A vssd1 vssd1 vccd1 vccd1 _12793_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ input5/X input280/X _17320_/S vssd1 vssd1 vccd1 vccd1 _17320_/X sky130_fd_sc_hd__mux2_1
X_14532_ _19302_/Q _17886_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19302_/D sky130_fd_sc_hd__mux2_1
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11795_/A _11795_/B _13416_/A vssd1 vssd1 vccd1 vccd1 _15734_/A sky130_fd_sc_hd__a21o_1
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _17251_/A _17275_/B _17269_/C vssd1 vssd1 vccd1 vccd1 _17251_/X sky130_fd_sc_hd__and3_1
X_14463_ _20227_/Q _19256_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14464_/B sky130_fd_sc_hd__mux2_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11675_ _20415_/Q _11676_/S _11653_/X _12063_/C1 vssd1 vssd1 vccd1 vccd1 _11675_/X
+ sky130_fd_sc_hd__o211a_1
X_16202_ _19625_/Q _17679_/A1 _16230_/S vssd1 vssd1 vccd1 vccd1 _19625_/D sky130_fd_sc_hd__mux2_1
X_13414_ _13414_/A _13414_/B vssd1 vssd1 vccd1 vccd1 _13414_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17182_ _20148_/Q _17950_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20148_/D sky130_fd_sc_hd__mux2_1
X_10626_ _12711_/A _19343_/Q _20698_/Q _10628_/S _10630_/C1 vssd1 vssd1 vccd1 vccd1
+ _10626_/X sky130_fd_sc_hd__a221o_1
X_14394_ _14394_/A _14394_/B vssd1 vssd1 vccd1 vccd1 _14394_/Y sky130_fd_sc_hd__xnor2_1
X_16133_ _16133_/A _16133_/B _16133_/C vssd1 vssd1 vccd1 vccd1 _16133_/X sky130_fd_sc_hd__and3_2
XFILLER_155_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13345_ _14295_/C1 _19232_/Q _14296_/A vssd1 vssd1 vccd1 vccd1 _13345_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ _19584_/Q _10556_/X _11229_/S vssd1 vssd1 vccd1 vccd1 _10558_/B sky130_fd_sc_hd__mux2_4
XFILLER_183_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _16064_/A _16064_/B _15814_/A vssd1 vssd1 vccd1 vccd1 _16064_/X sky130_fd_sc_hd__or3b_1
X_13276_ _13571_/A _13571_/B vssd1 vssd1 vccd1 vccd1 _13586_/C sky130_fd_sc_hd__and2_2
XFILLER_170_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10488_ _10478_/X _10481_/X _10484_/X _10487_/X _12513_/C _09621_/A vssd1 vssd1 vccd1
+ vccd1 _10488_/X sky130_fd_sc_hd__mux4_2
XFILLER_136_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15015_ _15021_/C _15018_/B vssd1 vssd1 vccd1 vccd1 _15015_/X sky130_fd_sc_hd__and2_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12227_ _09503_/A _12220_/X _12221_/X vssd1 vssd1 vccd1 vccd1 _12227_/X sky130_fd_sc_hd__o21a_1
XFILLER_142_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19823_ _20047_/CLK _19823_/D vssd1 vssd1 vccd1 vccd1 _19823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12158_ _12403_/A1 _12157_/Y _12158_/B1 vssd1 vssd1 vccd1 vccd1 _12158_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_256_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11109_ _12337_/A _20495_/Q _12248_/B1 _20527_/Q vssd1 vssd1 vccd1 vccd1 _11109_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19754_ _20962_/CLK _19754_/D vssd1 vssd1 vccd1 vccd1 _19754_/Q sky130_fd_sc_hd__dfxtp_2
X_16966_ _16974_/A1 _16965_/X _16982_/B1 vssd1 vssd1 vccd1 vccd1 _16966_/Y sky130_fd_sc_hd__o21ai_2
X_12089_ _20144_/Q _20112_/Q _12097_/S vssd1 vssd1 vccd1 vccd1 _12089_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18705_ _20953_/Q _18195_/Y _18719_/S vssd1 vssd1 vccd1 vccd1 _18706_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15917_ _15973_/A1 _15916_/X _15904_/Y vssd1 vssd1 vccd1 vccd1 _15917_/X sky130_fd_sc_hd__a21bo_1
XFILLER_225_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19685_ _20708_/CLK _19685_/D vssd1 vssd1 vccd1 vccd1 _19685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16897_ _20415_/Q _16963_/A2 _16963_/B1 vssd1 vssd1 vccd1 vccd1 _16897_/X sky130_fd_sc_hd__a21o_1
XFILLER_225_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18636_ _19512_/Q _18671_/B vssd1 vssd1 vccd1 vccd1 _18636_/Y sky130_fd_sc_hd__nand2_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _15365_/A _15846_/X _15847_/X _15844_/X vssd1 vssd1 vccd1 vccd1 _15848_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_225_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18567_ _20914_/Q _18619_/B _18566_/X vssd1 vssd1 vccd1 vccd1 _18568_/B sky130_fd_sc_hd__a21oi_1
X_15779_ _19755_/Q _15999_/A2 _15778_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15779_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17518_ _20294_/Q _17522_/B vssd1 vssd1 vccd1 vccd1 _17518_/Y sky130_fd_sc_hd__nand2_1
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18498_ _18856_/A _18498_/B vssd1 vssd1 vccd1 vccd1 _20892_/D sky130_fd_sc_hd__nor2_1
XFILLER_232_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17449_ _17460_/A2 _17446_/A _17447_/X _17448_/X _17434_/A vssd1 vssd1 vccd1 vccd1
+ _20263_/D sky130_fd_sc_hd__o221a_1
XFILLER_221_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20460_ _20687_/CLK _20460_/D vssd1 vssd1 vccd1 vccd1 _20460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19119_ _19505_/CLK _19119_/D vssd1 vssd1 vccd1 vccd1 _19119_/Q sky130_fd_sc_hd__dfxtp_2
X_20391_ _20583_/CLK _20391_/D vssd1 vssd1 vccd1 vccd1 _20391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21012_ _21018_/CLK _21012_/D vssd1 vssd1 vccd1 vccd1 _21012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput287 _13829_/X vssd1 vssd1 vccd1 vccd1 addr0[2] sky130_fd_sc_hd__buf_4
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput298 _13785_/X vssd1 vssd1 vccd1 vccd1 addr1[4] sky130_fd_sc_hd__buf_4
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ _09694_/X _09697_/X _09704_/X _11904_/S _12137_/A1 vssd1 vssd1 vccd1 vccd1
+ _09705_/X sky130_fd_sc_hd__o221a_1
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09636_ _09643_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _10553_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09567_ _09567_/A _19154_/Q _12579_/C vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__or3b_4
XFILLER_243_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09498_ _19216_/Q vssd1 vssd1 vccd1 vccd1 _09498_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20727_ _20727_/CLK _20727_/D vssd1 vssd1 vccd1 vccd1 _20727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11460_ _19351_/Q _20706_/Q _12185_/S vssd1 vssd1 vccd1 vccd1 _11460_/X sky130_fd_sc_hd__mux2_1
X_20658_ _20658_/CLK _20658_/D vssd1 vssd1 vccd1 vccd1 _20658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ _11290_/A _19313_/Q _11290_/C vssd1 vssd1 vccd1 vccd1 _10411_/X sky130_fd_sc_hd__or3_1
XFILLER_137_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11391_ _11391_/A _20665_/Q _11391_/C vssd1 vssd1 vccd1 vccd1 _11391_/X sky130_fd_sc_hd__or3_1
XFILLER_136_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20589_ _20657_/CLK _20589_/D vssd1 vssd1 vccd1 vccd1 _20589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13130_ _12629_/Y _13106_/B _12909_/X _13107_/A vssd1 vssd1 vccd1 vccd1 _13130_/X
+ sky130_fd_sc_hd__a31o_1
X_10342_ _19412_/Q _20571_/Q _10518_/S vssd1 vssd1 vccd1 vccd1 _10342_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _20949_/Q _20883_/Q _13505_/A vssd1 vssd1 vccd1 vccd1 _13518_/A sky130_fd_sc_hd__a21oi_2
XFILLER_180_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10273_ _12277_/A1 _17901_/A1 _10272_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _15593_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12012_ _12006_/X _12011_/X _12012_/S vssd1 vssd1 vccd1 vccd1 _12012_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1402 _12081_/S0 vssd1 vssd1 vccd1 vccd1 _10628_/S sky130_fd_sc_hd__buf_6
Xfanout1413 _11203_/S vssd1 vssd1 vccd1 vccd1 _11211_/S sky130_fd_sc_hd__buf_6
XFILLER_160_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1424 _11393_/S0 vssd1 vssd1 vccd1 vccd1 _12344_/S sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_39_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21047_/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16820_ _16846_/A _09522_/Y _16809_/X _16819_/Y vssd1 vssd1 vccd1 vccd1 _16820_/X
+ sky130_fd_sc_hd__o211a_4
Xfanout1435 _12085_/B2 vssd1 vssd1 vccd1 vccd1 _11718_/S sky130_fd_sc_hd__buf_6
Xfanout1446 _10611_/B vssd1 vssd1 vccd1 vccd1 _11846_/C sky130_fd_sc_hd__buf_6
Xfanout1457 _11391_/C vssd1 vssd1 vccd1 vccd1 _12337_/C sky130_fd_sc_hd__buf_6
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1468 _11204_/S vssd1 vssd1 vccd1 vccd1 _12011_/S sky130_fd_sc_hd__buf_6
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1479 _11945_/S vssd1 vssd1 vccd1 vccd1 _12186_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16751_ _16982_/B1 _16748_/X _16750_/X _16866_/B2 vssd1 vssd1 vccd1 vccd1 _16752_/B
+ sky130_fd_sc_hd__o2bb2a_2
Xfanout492 _17885_/X vssd1 vssd1 vccd1 vccd1 _17914_/S sky130_fd_sc_hd__clkbuf_16
X_13963_ _14041_/A1 _13969_/A2 _10809_/X _14041_/B1 _19836_/Q vssd1 vssd1 vccd1 vccd1
+ _14055_/C sky130_fd_sc_hd__o32a_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15702_ _15890_/B _15685_/Y _15701_/X _15976_/B2 vssd1 vssd1 vccd1 vccd1 _15702_/X
+ sky130_fd_sc_hd__o22a_1
X_19470_ _20718_/CLK _19470_/D vssd1 vssd1 vccd1 vccd1 _19470_/Q sky130_fd_sc_hd__dfxtp_1
X_12914_ _14433_/A _12914_/B vssd1 vssd1 vccd1 vccd1 _12914_/Y sky130_fd_sc_hd__xnor2_2
X_16682_ _19937_/Q _17894_/A1 _16704_/S vssd1 vssd1 vccd1 vccd1 _19937_/D sky130_fd_sc_hd__mux2_1
X_13894_ _19112_/Q _19050_/S _13896_/B1 _11367_/A _14458_/A vssd1 vssd1 vccd1 vccd1
+ _19112_/D sky130_fd_sc_hd__o221a_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18421_ _20865_/Q _18235_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18422_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15633_ _15322_/X _15323_/X _15140_/S vssd1 vssd1 vccd1 vccd1 _15633_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12845_ _12845_/A _12845_/B vssd1 vssd1 vccd1 vccd1 _12846_/A sky130_fd_sc_hd__or2_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _20831_/Q _18363_/B _18351_/Y _18352_/C1 vssd1 vssd1 vccd1 vccd1 _20831_/D
+ sky130_fd_sc_hd__o211a_1
X_15564_ _20736_/Q _16041_/A2 _16041_/B1 _20768_/Q vssd1 vssd1 vccd1 vccd1 _15564_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12774_/X _12775_/Y _12752_/B vssd1 vssd1 vccd1 vccd1 _12776_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_42_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _20206_/Q _17321_/A2 _17324_/C1 _17302_/X vssd1 vssd1 vccd1 vccd1 _17303_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_187_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11727_ _11729_/A _11733_/B vssd1 vssd1 vccd1 vccd1 _13166_/B sky130_fd_sc_hd__or2_2
X_14515_ _19293_/Q _17178_/A1 _14516_/S vssd1 vssd1 vccd1 vccd1 _19293_/D sky130_fd_sc_hd__mux2_1
XFILLER_222_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18283_ _19552_/Q _18308_/B vssd1 vssd1 vccd1 vccd1 _18283_/Y sky130_fd_sc_hd__nand2b_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ _11768_/X _15127_/B _15494_/X _12579_/D vssd1 vssd1 vccd1 vccd1 _15495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17234_ _17235_/A _17235_/B vssd1 vssd1 vccd1 vccd1 _17234_/X sky130_fd_sc_hd__and2_1
XFILLER_159_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14446_ _18985_/A _14446_/B vssd1 vssd1 vccd1 vccd1 _19247_/D sky130_fd_sc_hd__and2_1
X_11658_ _10430_/S _12051_/A1 _19352_/Q _12046_/B1 vssd1 vssd1 vccd1 vccd1 _11658_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10609_ _20634_/Q _11693_/B _11852_/B2 vssd1 vssd1 vccd1 vccd1 _10609_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17165_ _20131_/Q _17199_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20131_/D sky130_fd_sc_hd__mux2_1
XFILLER_196_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14377_ _14373_/B _14376_/Y _14417_/S vssd1 vssd1 vccd1 vccd1 _14377_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11589_ _11587_/X _11588_/X _11980_/S vssd1 vssd1 vccd1 vccd1 _11589_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16116_ _19582_/Q _16127_/A2 _16115_/X _16129_/B1 vssd1 vssd1 vccd1 vccd1 _19582_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13328_ _13355_/B _13328_/B vssd1 vssd1 vccd1 vccd1 _13328_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17096_ _20066_/Q _17096_/A1 _17111_/S vssd1 vssd1 vccd1 vccd1 _20066_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16047_ _20817_/Q _16047_/A2 _16041_/X _16049_/A1 _16046_/X vssd1 vssd1 vccd1 vccd1
+ _16047_/X sky130_fd_sc_hd__a221o_1
X_13259_ _13258_/A _13258_/B _13258_/C vssd1 vssd1 vccd1 vccd1 _13259_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_282_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19806_ _20665_/CLK _19806_/D vssd1 vssd1 vccd1 vccd1 _19806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17998_ _17998_/A _18003_/C vssd1 vssd1 vccd1 vccd1 _17998_/Y sky130_fd_sc_hd__nor2_1
XFILLER_257_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19737_ _20725_/CLK _19737_/D vssd1 vssd1 vccd1 vccd1 _19737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16949_ _16974_/A1 _16948_/X _16982_/B1 vssd1 vssd1 vccd1 vccd1 _16949_/Y sky130_fd_sc_hd__o21ai_2
Xfanout1980 _18814_/A vssd1 vssd1 vccd1 vccd1 _18598_/A sky130_fd_sc_hd__buf_6
XFILLER_38_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1991 _19051_/A vssd1 vssd1 vccd1 vccd1 _18054_/A sky130_fd_sc_hd__buf_4
XFILLER_77_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19668_ _20563_/CLK _19668_/D vssd1 vssd1 vccd1 vccd1 _19668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18619_ _20928_/Q _18619_/B vssd1 vssd1 vccd1 vccd1 _18619_/Y sky130_fd_sc_hd__nand2_1
XFILLER_213_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19599_ _19606_/CLK _19599_/D vssd1 vssd1 vccd1 vccd1 _19599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20512_ _20676_/CLK _20512_/D vssd1 vssd1 vccd1 vccd1 _20512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20443_ _20557_/CLK _20443_/D vssd1 vssd1 vccd1 vccd1 _20443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20374_ _20438_/CLK _20374_/D vssd1 vssd1 vccd1 vccd1 _20374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10960_ _11021_/A _20122_/Q _20090_/Q _11035_/S vssd1 vssd1 vccd1 vccd1 _10960_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09619_ _16454_/B _10152_/S _09689_/A _17538_/C vssd1 vssd1 vccd1 vccd1 _09619_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10891_ _09672_/A _13960_/A2 _10890_/X _11228_/B1 _19835_/Q vssd1 vssd1 vccd1 vccd1
+ _16077_/A sky130_fd_sc_hd__o32ai_4
XFILLER_216_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12630_ _19501_/Q _12639_/A vssd1 vssd1 vccd1 vccd1 _12630_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_157_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20962_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XPHY_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12561_ _12561_/A _13143_/B vssd1 vssd1 vccd1 vccd1 _12562_/A sky130_fd_sc_hd__nor2_8
XFILLER_240_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11512_ _11502_/X _11504_/X _11511_/X _12135_/A _12137_/A1 vssd1 vssd1 vccd1 vccd1
+ _11512_/X sky130_fd_sc_hd__o221a_1
X_14300_ _19512_/Q _14300_/B vssd1 vssd1 vccd1 vccd1 _14301_/B sky130_fd_sc_hd__or2_1
X_15280_ _19707_/Q _15279_/X _15454_/S vssd1 vssd1 vccd1 vccd1 _15280_/X sky130_fd_sc_hd__mux2_2
X_12492_ _19495_/Q _13107_/A vssd1 vssd1 vccd1 vccd1 _12493_/B sky130_fd_sc_hd__xnor2_1
XFILLER_221_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _14232_/A _14232_/B vssd1 vssd1 vccd1 vccd1 _14240_/B sky130_fd_sc_hd__nand2_1
X_11443_ _19640_/Q _12146_/S _11428_/X _12150_/S vssd1 vssd1 vccd1 vccd1 _11443_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14162_ _14162_/A _14162_/B vssd1 vssd1 vccd1 vccd1 _14162_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11374_ _11372_/X _11373_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _11374_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ _13100_/A _13100_/B _13112_/X vssd1 vssd1 vccd1 vccd1 _13245_/A sky130_fd_sc_hd__a21oi_4
XFILLER_166_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10325_ _11250_/S _10324_/X _10323_/X _11274_/B2 vssd1 vssd1 vccd1 vccd1 _10325_/X
+ sky130_fd_sc_hd__a211o_1
X_14093_ _14099_/A _14099_/B _14093_/C vssd1 vssd1 vccd1 vccd1 _14093_/X sky130_fd_sc_hd__or3_1
X_18970_ _18683_/Y _18970_/A2 _18968_/Y _18969_/Y vssd1 vssd1 vccd1 vccd1 _18970_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17921_ _20690_/Q _17921_/A1 _17934_/S vssd1 vssd1 vccd1 vccd1 _20690_/D sky130_fd_sc_hd__mux2_1
X_13044_ _20956_/Q _20890_/Q vssd1 vssd1 vccd1 vccd1 _13604_/B sky130_fd_sc_hd__nand2_2
X_10256_ _20476_/Q _11042_/B _11378_/S vssd1 vssd1 vccd1 vccd1 _10256_/X sky130_fd_sc_hd__o21a_1
XFILLER_239_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1210 _15026_/Y vssd1 vssd1 vccd1 vccd1 _16051_/A1 sky130_fd_sc_hd__buf_4
Xfanout1221 _13355_/B vssd1 vssd1 vccd1 vccd1 _13370_/B sky130_fd_sc_hd__clkbuf_4
X_17852_ _20625_/Q _17852_/A1 _17883_/S vssd1 vssd1 vccd1 vccd1 _20625_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1232 _12493_/A vssd1 vssd1 vccd1 vccd1 _12784_/B sky130_fd_sc_hd__buf_6
XFILLER_266_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10187_ _10937_/A _20506_/Q _11211_/S _20538_/Q vssd1 vssd1 vccd1 vccd1 _10187_/X
+ sky130_fd_sc_hd__o22a_1
Xfanout1243 _17337_/Y vssd1 vssd1 vccd1 vccd1 _17382_/B1 sky130_fd_sc_hd__buf_6
XFILLER_121_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16803_ _19968_/Q _16887_/A _16802_/Y _16896_/C1 vssd1 vssd1 vccd1 vccd1 _19968_/D
+ sky130_fd_sc_hd__a211o_1
Xfanout1265 _13675_/A vssd1 vssd1 vccd1 vccd1 _12401_/B1 sky130_fd_sc_hd__buf_6
Xfanout1276 _16034_/S vssd1 vssd1 vccd1 vccd1 _15895_/S sky130_fd_sc_hd__buf_12
XFILLER_266_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17783_ _20560_/Q _17923_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20560_/D sky130_fd_sc_hd__mux2_1
Xfanout1287 _12581_/A vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__buf_8
X_14995_ _15314_/D _15022_/D vssd1 vssd1 vccd1 vccd1 _14995_/Y sky130_fd_sc_hd__nor2_1
Xfanout1298 _14330_/B1 vssd1 vssd1 vccd1 vccd1 _14431_/B1 sky130_fd_sc_hd__buf_6
XFILLER_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19522_ _20296_/CLK _19522_/D vssd1 vssd1 vccd1 vccd1 _19522_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_207_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16734_ _19216_/Q _16862_/A2 _17005_/A2 _19085_/Q _16733_/X vssd1 vssd1 vccd1 vccd1
+ _16734_/X sky130_fd_sc_hd__o221a_1
X_13946_ _19148_/Q _13941_/B _13946_/B1 _13100_/X vssd1 vssd1 vccd1 vccd1 _19148_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19453_ _20712_/CLK _19453_/D vssd1 vssd1 vccd1 vccd1 _19453_/Q sky130_fd_sc_hd__dfxtp_1
X_16665_ _19922_/Q _17945_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19922_/D sky130_fd_sc_hd__mux2_1
X_13877_ _19095_/Q _13953_/A2 _13881_/B1 _19161_/Q _15288_/C1 vssd1 vssd1 vccd1 vccd1
+ _19095_/D sky130_fd_sc_hd__o221a_1
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18404_ _18418_/A _18404_/B vssd1 vssd1 vccd1 vccd1 _20856_/D sky130_fd_sc_hd__and2_1
X_15616_ _15890_/A _15527_/B _15614_/X _15615_/X _15609_/X vssd1 vssd1 vccd1 vccd1
+ _15616_/X sky130_fd_sc_hd__o41a_1
X_12828_ _12828_/A _12832_/B vssd1 vssd1 vccd1 vccd1 _12829_/D sky130_fd_sc_hd__nor2_2
X_19384_ _20675_/CLK _19384_/D vssd1 vssd1 vccd1 vccd1 _19384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16596_ _16598_/A _16594_/B _16595_/Y vssd1 vssd1 vccd1 vccd1 _16596_/X sky130_fd_sc_hd__o21a_1
XFILLER_250_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18335_ _18480_/B _18349_/B vssd1 vssd1 vccd1 vccd1 _18335_/Y sky130_fd_sc_hd__nand2_1
X_15547_ _15066_/S _15122_/Y _15545_/Y _15546_/Y vssd1 vssd1 vccd1 vccd1 _15547_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12757_/Y _12758_/X _12751_/X _12752_/Y vssd1 vssd1 vccd1 vccd1 _12759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18266_ _20807_/Q _18265_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18267_/B sky130_fd_sc_hd__mux2_1
X_15478_ _20893_/Q _14971_/A _15566_/B1 _15477_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15478_/X sky130_fd_sc_hd__a221o_1
XFILLER_147_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17217_ _20181_/Q _17708_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20181_/D sky130_fd_sc_hd__mux2_1
X_14429_ _13111_/Y _14428_/X _14437_/B _14437_/A vssd1 vssd1 vccd1 vccd1 _14429_/X
+ sky130_fd_sc_hd__a211o_1
X_18197_ _18418_/A _18197_/B vssd1 vssd1 vccd1 vccd1 _20793_/D sky130_fd_sc_hd__and2_1
XFILLER_129_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17148_ _20116_/Q _17950_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20116_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09970_ _20417_/Q _12149_/S _09948_/X _09901_/S vssd1 vssd1 vccd1 vccd1 _09970_/X
+ sky130_fd_sc_hd__o211a_1
X_17079_ _20051_/Q _17915_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20051_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20090_ _20672_/CLK _20090_/D vssd1 vssd1 vccd1 vccd1 _20090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20992_ _21025_/CLK _20992_/D vssd1 vssd1 vccd1 vccd1 _20992_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20426_ _20426_/CLK _20426_/D vssd1 vssd1 vccd1 vccd1 _20426_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20357_ _20678_/CLK _20357_/D vssd1 vssd1 vccd1 vccd1 _20357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _19506_/Q _15504_/A _11398_/S vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11090_ _19800_/Q _19304_/Q _11090_/S vssd1 vssd1 vccd1 vccd1 _11090_/X sky130_fd_sc_hd__mux2_1
X_20288_ _21010_/CLK _20288_/D vssd1 vssd1 vccd1 vccd1 _20288_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ _11236_/B _10041_/B vssd1 vssd1 vccd1 vccd1 _10041_/Y sky130_fd_sc_hd__nand2_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xsplit9 split9/A vssd1 vssd1 vccd1 vccd1 split9/X sky130_fd_sc_hd__clkbuf_2
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13800_ _13816_/A1 _13673_/Y _13816_/B1 input246/X vssd1 vssd1 vccd1 vccd1 _13800_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14780_ _19137_/Q _14798_/A2 _14779_/X _14780_/C1 vssd1 vssd1 vccd1 vccd1 _19514_/D
+ sky130_fd_sc_hd__o211a_1
X_11992_ _12056_/S _11991_/X _11990_/X _12144_/A1 vssd1 vssd1 vccd1 vccd1 _11992_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10943_ _19370_/Q _11291_/A2 _10941_/X _11291_/B2 _10942_/X vssd1 vssd1 vccd1 vccd1
+ _10943_/X sky130_fd_sc_hd__o221a_1
X_13731_ _13740_/B _13693_/X _13659_/B _13714_/S vssd1 vssd1 vccd1 vccd1 _13731_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_272_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16450_ _19763_/Q _19764_/Q _16450_/C vssd1 vssd1 vccd1 vccd1 _16451_/C sky130_fd_sc_hd__and3_1
X_10874_ _10871_/X _10872_/X _10873_/X _09731_/A _10866_/A vssd1 vssd1 vccd1 vccd1
+ _10874_/X sky130_fd_sc_hd__a221o_1
XFILLER_189_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13662_ _13662_/A vssd1 vssd1 vccd1 vccd1 _13735_/B sky130_fd_sc_hd__inv_6
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _19502_/Q _10935_/B _15400_/X vssd1 vssd1 vccd1 vccd1 _15402_/B sky130_fd_sc_hd__o21ai_2
X_12613_ _19521_/Q _12889_/A vssd1 vssd1 vccd1 vccd1 _12901_/B sky130_fd_sc_hd__and2_1
X_16381_ _19738_/Q _16380_/B _16381_/B1 vssd1 vssd1 vccd1 vccd1 _16382_/B sky130_fd_sc_hd__o21ai_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _18462_/A _13592_/X _13589_/X _13609_/A vssd1 vssd1 vccd1 vccd1 _13593_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18120_ _18126_/A _18120_/B vssd1 vssd1 vccd1 vccd1 _18120_/Y sky130_fd_sc_hd__nor2_1
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15332_ _19709_/Q _15475_/A2 _15475_/B1 _19741_/Q vssd1 vssd1 vccd1 vccd1 _15332_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_212_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12544_ _20875_/Q _12548_/B _12544_/C vssd1 vssd1 vccd1 vccd1 _12550_/C sky130_fd_sc_hd__and3_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18051_ _20756_/Q _18053_/C _18050_/Y vssd1 vssd1 vccd1 vccd1 _20756_/D sky130_fd_sc_hd__o21a_1
XFILLER_185_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15263_ _10885_/A _15500_/A0 _14878_/B vssd1 vssd1 vccd1 vccd1 _15263_/Y sky130_fd_sc_hd__a21oi_1
X_12475_ _12454_/A _12454_/B _12454_/C _15983_/A vssd1 vssd1 vccd1 vccd1 _12475_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17002_ _19991_/Q _17012_/A2 _17001_/Y _17998_/A vssd1 vssd1 vccd1 vccd1 _19991_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11426_ _20350_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _11426_/X sky130_fd_sc_hd__or2_1
X_14214_ _14255_/A _16068_/B _14214_/C vssd1 vssd1 vccd1 vccd1 _14214_/X sky130_fd_sc_hd__or3_1
XANTENNA_6 _15340_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ _20917_/Q _15567_/A2 _15193_/X vssd1 vssd1 vccd1 vccd1 _15194_/X sky130_fd_sc_hd__o21a_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_54_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20061_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14145_ _19217_/Q _14256_/A2 _14144_/X _18698_/A vssd1 vssd1 vccd1 vccd1 _19217_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11357_ _19631_/Q _19937_/Q _12300_/S vssd1 vssd1 vccd1 vccd1 _11357_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10308_ _10306_/X _10307_/X _10308_/S vssd1 vssd1 vccd1 vccd1 _10308_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14076_ _19197_/Q _14108_/A2 _14075_/X _16129_/B1 vssd1 vssd1 vccd1 vccd1 _19197_/D
+ sky130_fd_sc_hd__o211a_1
X_18953_ _18980_/A _18953_/B vssd1 vssd1 vccd1 vccd1 _21007_/D sky130_fd_sc_hd__nor2_1
X_11288_ _11286_/X _11287_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11288_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13027_ _20965_/Q _20899_/Q vssd1 vssd1 vccd1 vccd1 _13303_/A sky130_fd_sc_hd__or2_2
XFILLER_79_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17904_ _20675_/Q _17904_/A1 _17912_/S vssd1 vssd1 vccd1 vccd1 _20675_/D sky130_fd_sc_hd__mux2_1
X_10239_ _09623_/B _10235_/X _10238_/X _09689_/C vssd1 vssd1 vccd1 vccd1 _10239_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18884_ _18891_/A _18884_/B vssd1 vssd1 vccd1 vccd1 _20997_/D sky130_fd_sc_hd__nor2_1
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1040 _17887_/A1 vssd1 vssd1 vccd1 vccd1 _17051_/A1 sky130_fd_sc_hd__buf_2
XFILLER_266_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1051 _11049_/B1 vssd1 vssd1 vccd1 vccd1 _17189_/A1 sky130_fd_sc_hd__buf_2
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1062 _17892_/A1 vssd1 vssd1 vccd1 vccd1 _17649_/A1 sky130_fd_sc_hd__buf_2
X_17835_ _20610_/Q _17835_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20610_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1073 _17919_/B vssd1 vssd1 vccd1 vccd1 _17851_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1084 _17950_/A1 vssd1 vssd1 vccd1 vccd1 _17707_/A1 sky130_fd_sc_hd__buf_4
XFILLER_281_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1095 _12210_/X vssd1 vssd1 vccd1 vccd1 _17949_/A1 sky130_fd_sc_hd__buf_6
XFILLER_282_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17766_ _20545_/Q _17906_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20545_/D sky130_fd_sc_hd__mux2_1
X_14978_ _15021_/B _14978_/B vssd1 vssd1 vccd1 vccd1 _14978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19505_ _19505_/CLK _19505_/D vssd1 vssd1 vccd1 vccd1 _19505_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_281_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16717_ _17461_/A _16716_/Y _16715_/A vssd1 vssd1 vccd1 vccd1 _16717_/X sky130_fd_sc_hd__a21o_2
XFILLER_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13929_ _19133_/Q _13906_/B _13932_/B1 _13359_/Y vssd1 vssd1 vccd1 vccd1 _19133_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17697_ _20481_/Q _17800_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20481_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19436_ _20084_/CLK _19436_/D vssd1 vssd1 vccd1 vccd1 _19436_/Q sky130_fd_sc_hd__dfxtp_1
X_16648_ _19905_/Q _17058_/A1 _16670_/S vssd1 vssd1 vccd1 vccd1 _19905_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19367_ _20658_/CLK _19367_/D vssd1 vssd1 vccd1 vccd1 _19367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16579_ _16591_/A _16579_/B vssd1 vssd1 vccd1 vccd1 _19855_/D sky130_fd_sc_hd__or2_1
XFILLER_222_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18318_ _18318_/A _18318_/B _18318_/C vssd1 vssd1 vccd1 vccd1 _18389_/C sky130_fd_sc_hd__or3_1
XFILLER_203_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19298_ _20664_/CLK _19298_/D vssd1 vssd1 vccd1 vccd1 _19298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18249_ _18248_/B _14300_/B _18248_/Y vssd1 vssd1 vccd1 vccd1 _18520_/B sky130_fd_sc_hd__o21ai_4
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20211_ _20766_/CLK _20211_/D vssd1 vssd1 vccd1 vccd1 _20211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20142_ _20481_/CLK _20142_/D vssd1 vssd1 vccd1 vccd1 _20142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09953_ _11903_/A1 _12120_/A1 _19354_/Q _12129_/S vssd1 vssd1 vccd1 vccd1 _09953_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_132_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20073_ _20480_/CLK _20073_/D vssd1 vssd1 vccd1 vccd1 _20073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _09882_/X _09883_/X _11513_/S vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__mux2_1
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_407 _17001_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_418 _18690_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_429 _13790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20975_ _21006_/CLK _20975_/D vssd1 vssd1 vccd1 vccd1 _20975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10590_ _19276_/Q _20063_/Q _11676_/S vssd1 vssd1 vccd1 vccd1 _10590_/X sky130_fd_sc_hd__mux2_1
XFILLER_278_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _19691_/Q _20179_/Q _12417_/S vssd1 vssd1 vccd1 vccd1 _12260_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11211_ _19866_/Q _19767_/Q _11211_/S vssd1 vssd1 vccd1 vccd1 _11211_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20409_ _20668_/CLK _20409_/D vssd1 vssd1 vccd1 vccd1 _20409_/Q sky130_fd_sc_hd__dfxtp_4
X_12191_ _09986_/C _12186_/X _12190_/X _12191_/C1 vssd1 vssd1 vccd1 vccd1 _12191_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11142_ _11239_/A1 _13960_/A2 _11141_/X _09648_/Y _19832_/Q vssd1 vssd1 vccd1 vccd1
+ _16071_/A sky130_fd_sc_hd__o32ai_4
XFILLER_134_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11073_ _19664_/Q _20152_/Q _11074_/S vssd1 vssd1 vccd1 vccd1 _11073_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15950_ _15949_/A _15948_/X _15949_/Y vssd1 vssd1 vccd1 vccd1 _15950_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_277_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput110 dout1[12] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_hd__clkbuf_2
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput121 dout1[22] vssd1 vssd1 vccd1 vccd1 input121/X sky130_fd_sc_hd__clkbuf_2
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput132 dout1[32] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__buf_2
X_10024_ _11326_/A _11326_/B vssd1 vssd1 vccd1 vccd1 _10024_/X sky130_fd_sc_hd__and2_4
X_14901_ _18136_/B _16720_/D vssd1 vssd1 vccd1 vccd1 _14901_/Y sky130_fd_sc_hd__nor2_1
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput143 dout1[42] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__buf_2
XFILLER_209_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput154 dout1[52] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__clkbuf_2
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15881_ _19759_/Q _15999_/A2 _15880_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15881_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput165 dout1[62] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_hd__clkbuf_2
XFILLER_264_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 irq[14] vssd1 vssd1 vccd1 vccd1 _12538_/C sky130_fd_sc_hd__clkbuf_2
X_17620_ _20376_/Q _17931_/A1 _17635_/S vssd1 vssd1 vccd1 vccd1 _20376_/D sky130_fd_sc_hd__mux2_1
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_172_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21000_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput187 jtag_tck vssd1 vssd1 vccd1 vccd1 _17420_/A sky130_fd_sc_hd__buf_4
XFILLER_48_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14832_ _14828_/X _14831_/X _15170_/A vssd1 vssd1 vccd1 vccd1 _14832_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput198 localMemory_wb_adr_i[17] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__clkbuf_2
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_101_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20725_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17551_ _20311_/Q _17687_/A1 _17570_/S vssd1 vssd1 vccd1 vccd1 _20311_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14763_ _19506_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14763_/X sky130_fd_sc_hd__or2_1
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _19793_/Q _11897_/B _11974_/X _12123_/C1 vssd1 vssd1 vccd1 vccd1 _11975_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _19809_/Q _17095_/A1 _16517_/S vssd1 vssd1 vccd1 vccd1 _19809_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13714_ _13752_/B _13713_/X _13714_/S vssd1 vssd1 vccd1 vccd1 _13716_/B sky130_fd_sc_hd__mux2_8
X_17482_ _20276_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17482_/Y sky130_fd_sc_hd__nand2_1
X_10926_ _09618_/A _10924_/X _10925_/X _11345_/S vssd1 vssd1 vccd1 vccd1 _10926_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14694_ _19453_/Q _17666_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19453_/D sky130_fd_sc_hd__mux2_1
X_19221_ _19223_/CLK _19221_/D vssd1 vssd1 vccd1 vccd1 _19221_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16433_ _19757_/Q _16434_/C _19758_/Q vssd1 vssd1 vccd1 vccd1 _16435_/B sky130_fd_sc_hd__a21oi_1
X_10857_ _12332_/A _20498_/Q _12334_/S0 _20530_/Q vssd1 vssd1 vccd1 vccd1 _10857_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_232_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13645_ _13663_/A _13663_/B _13708_/B vssd1 vssd1 vccd1 vccd1 _13645_/X sky130_fd_sc_hd__and3_4
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19152_ _19621_/CLK _19152_/D vssd1 vssd1 vccd1 vccd1 _19152_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _19732_/Q _16364_/B vssd1 vssd1 vccd1 vccd1 _16370_/C sky130_fd_sc_hd__and2_2
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _12427_/A1 _20124_/Q _20092_/Q _11126_/B vssd1 vssd1 vccd1 vccd1 _10788_/X
+ sky130_fd_sc_hd__a22o_1
X_13576_ _20922_/Q _13602_/A1 _13575_/X _18616_/B vssd1 vssd1 vccd1 vccd1 _13576_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _20776_/Q _18103_/B vssd1 vssd1 vccd1 vccd1 _18109_/C sky130_fd_sc_hd__and2_2
X_15315_ _15323_/A _14965_/X _14972_/X _15313_/X _15314_/X vssd1 vssd1 vccd1 vccd1
+ _15315_/X sky130_fd_sc_hd__o311a_1
XFILLER_185_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19083_ _20428_/Q vssd1 vssd1 vccd1 vccd1 _20428_/D sky130_fd_sc_hd__clkbuf_2
X_12527_ _19215_/Q _18462_/A _13575_/C vssd1 vssd1 vccd1 vccd1 _12527_/X sky130_fd_sc_hd__and3_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16295_ _19706_/Q _16293_/A _16381_/B1 vssd1 vssd1 vccd1 vccd1 _16296_/B sky130_fd_sc_hd__o21ai_1
XFILLER_158_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18034_ _18795_/A _18034_/B vssd1 vssd1 vccd1 vccd1 _18034_/Y sky130_fd_sc_hd__nor2_1
X_15246_ _15246_/A _15246_/B _15246_/C vssd1 vssd1 vccd1 vccd1 _15248_/B sky130_fd_sc_hd__or3_1
X_12458_ _12565_/B _12471_/B vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__and2_1
XFILLER_160_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11409_ _11409_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11409_/X sky130_fd_sc_hd__and2_1
X_12389_ _20427_/Q _20363_/Q _12389_/S vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15177_ _15612_/S _15164_/X _15176_/X vssd1 vssd1 vccd1 vccd1 _15177_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14128_ _20267_/Q _14117_/A _14216_/B1 input226/X vssd1 vssd1 vccd1 vccd1 _14130_/B
+ sky130_fd_sc_hd__a22o_4
X_19985_ _19992_/CLK _19985_/D vssd1 vssd1 vccd1 vccd1 _19985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14059_ _14107_/A _14069_/B _14059_/C vssd1 vssd1 vccd1 vccd1 _14059_/X sky130_fd_sc_hd__or3_1
X_18936_ _18663_/Y _18970_/A2 _18934_/Y _18935_/Y vssd1 vssd1 vccd1 vccd1 _18936_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_268_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18867_ _18624_/Y _18867_/A2 _18865_/Y _18866_/Y vssd1 vssd1 vccd1 vccd1 _18867_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_267_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17818_ _20593_/Q _17890_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20593_/D sky130_fd_sc_hd__mux2_1
XFILLER_283_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18798_ _18585_/Y _18818_/A2 _18797_/X _18901_/S vssd1 vssd1 vccd1 vccd1 _18798_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17749_ _20528_/Q _17889_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20528_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20760_ _20760_/CLK _20760_/D vssd1 vssd1 vccd1 vccd1 _20760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19419_ _20714_/CLK _19419_/D vssd1 vssd1 vccd1 vccd1 _19419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20691_ _20720_/CLK _20691_/D vssd1 vssd1 vccd1 vccd1 _20691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout800 _12479_/A vssd1 vssd1 vccd1 vccd1 _14803_/A1 sky130_fd_sc_hd__buf_6
XFILLER_277_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout811 _12590_/Y vssd1 vssd1 vccd1 vccd1 _12592_/C sky130_fd_sc_hd__buf_6
XFILLER_277_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20125_ _20468_/CLK _20125_/D vssd1 vssd1 vccd1 vccd1 _20125_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1809 _19528_/Q vssd1 vssd1 vccd1 vccd1 _15103_/A1 sky130_fd_sc_hd__buf_2
Xfanout822 _15323_/B vssd1 vssd1 vccd1 vccd1 _15566_/B1 sky130_fd_sc_hd__buf_8
X_09936_ _12194_/A1 _09936_/A2 _09935_/X _12194_/B2 vssd1 vssd1 vccd1 vccd1 _15768_/A
+ sky130_fd_sc_hd__a22o_2
Xfanout833 _18981_/X vssd1 vssd1 vccd1 vccd1 _18983_/B sky130_fd_sc_hd__clkbuf_8
Xfanout844 _18357_/B vssd1 vssd1 vccd1 vccd1 _18387_/B sky130_fd_sc_hd__clkbuf_4
Xfanout855 _16047_/A2 vssd1 vssd1 vccd1 vccd1 _15016_/A sky130_fd_sc_hd__buf_6
XFILLER_246_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout866 _15993_/S vssd1 vssd1 vccd1 vccd1 _16040_/S sky130_fd_sc_hd__buf_8
X_20056_ _20061_/CLK _20056_/D vssd1 vssd1 vccd1 vccd1 _20056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout877 _14948_/Y vssd1 vssd1 vccd1 vccd1 _15604_/A2 sky130_fd_sc_hd__buf_4
X_09867_ _11242_/A1 _14011_/A2 _09866_/X _11242_/B1 _19852_/Q vssd1 vssd1 vccd1 vccd1
+ _09867_/X sky130_fd_sc_hd__o32a_1
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout888 _18688_/A2 vssd1 vssd1 vccd1 vccd1 _18684_/A2 sky130_fd_sc_hd__buf_6
XFILLER_245_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout899 _15996_/B1 vssd1 vssd1 vccd1 vccd1 _16016_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_246_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09798_ _10430_/S _20711_/Q _10426_/S _09797_/X vssd1 vssd1 vccd1 vccd1 _09798_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_261_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 _19838_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_237 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_248 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11760_ _15763_/A _15763_/B _11752_/X _11757_/Y vssd1 vssd1 vccd1 vccd1 _11883_/C
+ sky130_fd_sc_hd__a211oi_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_259 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ _20990_/CLK _20958_/D vssd1 vssd1 vccd1 vccd1 _20958_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_199_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _12420_/B1 _10710_/X _10709_/X vssd1 vssd1 vccd1 vccd1 _10711_/X sky130_fd_sc_hd__o21a_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11922_/A1 _13712_/A _12158_/B1 vssd1 vssd1 vccd1 vccd1 _11691_/Y sky130_fd_sc_hd__o21ai_1
X_20889_ _21019_/CLK _20889_/D vssd1 vssd1 vccd1 vccd1 _20889_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13430_ _13430_/A vssd1 vssd1 vccd1 vccd1 _13430_/Y sky130_fd_sc_hd__inv_2
X_10642_ _10638_/B _10642_/B vssd1 vssd1 vccd1 vccd1 _11766_/B sky130_fd_sc_hd__nand2b_2
XFILLER_167_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _13361_/A _13361_/B _13361_/C _13361_/D vssd1 vssd1 vccd1 vccd1 _13388_/B
+ sky130_fd_sc_hd__or4_1
X_10573_ _10057_/S _10581_/A1 _19471_/Q _12136_/B1 vssd1 vssd1 vccd1 vccd1 _10573_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15100_ _15520_/B2 _15099_/X _15098_/X vssd1 vssd1 vccd1 vccd1 _15100_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12312_ _12312_/A1 _20524_/Q _12309_/S _12294_/X vssd1 vssd1 vccd1 vccd1 _12312_/X
+ sky130_fd_sc_hd__o211a_1
X_16080_ _19564_/Q _16079_/B _16079_/Y _16097_/B1 vssd1 vssd1 vccd1 vccd1 _19564_/D
+ sky130_fd_sc_hd__o211a_1
X_13292_ _20959_/Q _13607_/B vssd1 vssd1 vccd1 vccd1 _13292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12243_ _11275_/A _12232_/X _12235_/X _12242_/X _12400_/A1 vssd1 vssd1 vccd1 vccd1
+ _12243_/X sky130_fd_sc_hd__a311o_2
XFILLER_177_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15031_ _19494_/Q _12578_/B _15030_/X vssd1 vssd1 vccd1 vccd1 _15031_/X sky130_fd_sc_hd__o21a_1
XFILLER_142_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12174_ _20146_/Q _20114_/Q _12174_/S vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11125_ _12357_/A1 _11124_/X _11123_/X vssd1 vssd1 vccd1 vccd1 _11125_/X sky130_fd_sc_hd__o21a_1
XFILLER_174_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19770_ _20465_/CLK _19770_/D vssd1 vssd1 vccd1 vccd1 _19770_/Q sky130_fd_sc_hd__dfxtp_1
X_16982_ _17008_/A1 _16981_/X _16982_/B1 vssd1 vssd1 vccd1 vccd1 _16982_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_150_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18721_ _20961_/Q _18235_/Y _18749_/S vssd1 vssd1 vccd1 vccd1 _18722_/B sky130_fd_sc_hd__mux2_1
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ _19529_/Q _09613_/A _09613_/B _19593_/Q vssd1 vssd1 vccd1 vccd1 _11056_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15933_ _19729_/Q _15933_/B vssd1 vssd1 vccd1 vccd1 _15933_/X sky130_fd_sc_hd__or2_1
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ _11946_/A1 _19354_/Q _20709_/Q _11947_/S _11946_/C1 vssd1 vssd1 vccd1 vccd1
+ _10007_/X sky130_fd_sc_hd__a221o_1
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18652_ _18532_/X _18684_/A2 _18650_/Y _18651_/Y vssd1 vssd1 vccd1 vccd1 _18653_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15864_ _16024_/A1 _15862_/X _15863_/X _15843_/A _15975_/B2 vssd1 vssd1 vccd1 vccd1
+ _15864_/X sky130_fd_sc_hd__a32o_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _20361_/Q _17948_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20361_/D sky130_fd_sc_hd__mux2_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _11414_/B _11734_/B _14815_/S vssd1 vssd1 vccd1 vccd1 _14815_/X sky130_fd_sc_hd__mux2_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _18783_/A _18583_/B vssd1 vssd1 vccd1 vccd1 _20918_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _15795_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15795_/Y sky130_fd_sc_hd__nand2_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17534_ _17537_/A _17537_/B _17533_/X _17532_/A vssd1 vssd1 vccd1 vccd1 _17534_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_233_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _19120_/Q _14764_/A2 _14745_/X _18714_/A vssd1 vssd1 vccd1 vccd1 _19497_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11958_ _11877_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__and2b_1
XFILLER_251_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _11275_/A _10905_/X _10908_/X _12311_/C1 vssd1 vssd1 vccd1 vccd1 _10909_/X
+ sky130_fd_sc_hd__o31a_1
X_17465_ _17495_/A1 _17464_/Y _18801_/A vssd1 vssd1 vccd1 vccd1 _20267_/D sky130_fd_sc_hd__a21oi_1
X_14677_ _19436_/Q _17683_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19436_/D sky130_fd_sc_hd__mux2_1
XFILLER_225_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11889_ _19890_/Q _19791_/Q _11889_/S vssd1 vssd1 vccd1 vccd1 _11889_/X sky130_fd_sc_hd__mux2_1
X_19204_ _20428_/CLK _19204_/D vssd1 vssd1 vccd1 vccd1 _19204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16416_ _19751_/Q _16418_/C _16415_/Y vssd1 vssd1 vccd1 vccd1 _19751_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13628_ _13478_/B _13240_/X _13439_/C _13765_/A vssd1 vssd1 vccd1 vccd1 _13628_/X
+ sky130_fd_sc_hd__a22o_4
X_17396_ _20246_/Q _17337_/B _17530_/A2 _20295_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17396_/X sky130_fd_sc_hd__a221o_1
XFILLER_220_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19135_ _19511_/CLK _19135_/D vssd1 vssd1 vccd1 vccd1 _19135_/Q sky130_fd_sc_hd__dfxtp_1
X_16347_ _18863_/A _16347_/B _16348_/B vssd1 vssd1 vccd1 vccd1 _19725_/D sky130_fd_sc_hd__nor3_1
X_13559_ _19222_/Q _13559_/B vssd1 vssd1 vccd1 vccd1 _13559_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_285_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19066_ _20411_/Q vssd1 vssd1 vccd1 vccd1 _20411_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16278_ _16278_/A _16278_/B vssd1 vssd1 vccd1 vccd1 _19694_/D sky130_fd_sc_hd__nor2_1
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18017_ _20744_/Q _18019_/C _18016_/Y vssd1 vssd1 vccd1 vccd1 _20744_/D sky130_fd_sc_hd__o21a_1
X_15229_ _09744_/B _12682_/A _16009_/B vssd1 vssd1 vccd1 vccd1 _15229_/X sky130_fd_sc_hd__mux2_1
Xoutput403 _13796_/X vssd1 vssd1 vccd1 vccd1 din0[5] sky130_fd_sc_hd__buf_4
Xoutput414 _19974_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[13] sky130_fd_sc_hd__buf_4
XFILLER_160_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput425 _19984_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[23] sky130_fd_sc_hd__buf_4
Xoutput436 _19965_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[4] sky130_fd_sc_hd__buf_4
Xoutput447 _20259_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[2] sky130_fd_sc_hd__buf_4
XFILLER_5_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput458 _19511_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[17] sky130_fd_sc_hd__buf_4
XFILLER_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput469 _19521_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[27] sky130_fd_sc_hd__buf_4
XFILLER_259_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19968_ _19978_/CLK _19968_/D vssd1 vssd1 vccd1 vccd1 _19968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09721_ _09719_/X _09720_/X _11917_/S vssd1 vssd1 vccd1 vccd1 _09721_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18919_ _19107_/Q _18954_/A2 _18967_/B1 _15816_/A vssd1 vssd1 vccd1 vccd1 _18920_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19899_ _20061_/CLK _19899_/D vssd1 vssd1 vccd1 vccd1 _19899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09652_ _11242_/A1 _14041_/A2 _09647_/X _09649_/X _11229_/S vssd1 vssd1 vccd1 vccd1
+ _09681_/C sky130_fd_sc_hd__o311ai_4
XFILLER_228_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09583_ _09583_/A _09583_/B _09588_/C vssd1 vssd1 vccd1 vccd1 _09606_/A sky130_fd_sc_hd__and3_1
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20812_ _20812_/CLK _20812_/D vssd1 vssd1 vccd1 vccd1 _20812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20743_ _21029_/CLK _20743_/D vssd1 vssd1 vccd1 vccd1 _20743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20674_ _20678_/CLK _20674_/D vssd1 vssd1 vccd1 vccd1 _20674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1606 _09618_/Y vssd1 vssd1 vccd1 vccd1 _11170_/B1 sky130_fd_sc_hd__buf_8
Xfanout1617 _09806_/S vssd1 vssd1 vccd1 vccd1 _12056_/S sky130_fd_sc_hd__buf_6
Xfanout630 _13881_/B1 vssd1 vssd1 vccd1 vccd1 _13900_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_266_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1628 _11359_/S vssd1 vssd1 vccd1 vccd1 _12317_/S sky130_fd_sc_hd__buf_4
XFILLER_278_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout641 _16178_/S vssd1 vssd1 vccd1 vccd1 _16164_/B sky130_fd_sc_hd__buf_4
Xfanout1639 _17524_/B vssd1 vssd1 vccd1 vccd1 _17522_/B sky130_fd_sc_hd__buf_4
X_20108_ _20568_/CLK _20108_/D vssd1 vssd1 vccd1 vccd1 _20108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_265_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09919_ _09986_/A _19483_/Q _19451_/Q _09931_/S _12016_/C1 vssd1 vssd1 vccd1 vccd1
+ _09919_/X sky130_fd_sc_hd__a221o_1
Xfanout652 _16036_/A2 vssd1 vssd1 vccd1 vccd1 _15980_/A2 sky130_fd_sc_hd__buf_4
Xfanout663 _14115_/Y vssd1 vssd1 vccd1 vccd1 _14397_/B sky130_fd_sc_hd__buf_4
Xfanout674 _13901_/X vssd1 vssd1 vccd1 vccd1 _13943_/S sky130_fd_sc_hd__buf_6
XFILLER_219_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout685 _13862_/X vssd1 vssd1 vccd1 vccd1 _13986_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_274_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout696 _14073_/B vssd1 vssd1 vccd1 vccd1 _14069_/B sky130_fd_sc_hd__buf_6
X_12930_ _12950_/B2 _12930_/B vssd1 vssd1 vccd1 vccd1 _12930_/X sky130_fd_sc_hd__and2b_2
X_20039_ _20681_/CLK _20039_/D vssd1 vssd1 vccd1 vccd1 _20039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12861_ _13248_/A _13332_/A _13346_/C vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__or3_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _17884_/A _17744_/A vssd1 vssd1 vccd1 vccd1 _14601_/C sky130_fd_sc_hd__nor2_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _20581_/Q _11897_/B _11811_/X _11892_/C1 vssd1 vssd1 vccd1 vccd1 _11812_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _16058_/A2 _15264_/B _15580_/S vssd1 vssd1 vccd1 vccd1 _15580_/X sky130_fd_sc_hd__mux2_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12701_/A _12701_/B _12791_/X vssd1 vssd1 vccd1 vccd1 _13346_/A sky130_fd_sc_hd__a21o_4
XFILLER_233_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _17919_/A _17574_/B _14531_/C vssd1 vssd1 vccd1 vccd1 _14531_/X sky130_fd_sc_hd__and3_4
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11743_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _13416_/A sky130_fd_sc_hd__nor2_8
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17250_ _20189_/Q _17268_/A2 _17248_/X _17249_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1
+ _20189_/D sky130_fd_sc_hd__o221a_1
XFILLER_159_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _18692_/A _14462_/B vssd1 vssd1 vccd1 vccd1 _19255_/D sky130_fd_sc_hd__and2_1
XFILLER_169_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11674_ _11995_/S _11673_/X _11672_/X _11684_/A1 vssd1 vssd1 vccd1 vccd1 _11674_/X
+ sky130_fd_sc_hd__a211o_1
X_16201_ _19624_/Q _17051_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19624_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13413_ _13413_/A _13413_/B vssd1 vssd1 vccd1 vccd1 _15816_/A sky130_fd_sc_hd__xor2_4
X_17181_ _20147_/Q _17949_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20147_/D sky130_fd_sc_hd__mux2_1
X_10625_ _19407_/Q _20566_/Q _10628_/S vssd1 vssd1 vccd1 vccd1 _10625_/X sky130_fd_sc_hd__mux2_1
X_14393_ _14382_/Y _14386_/B _14384_/B vssd1 vssd1 vccd1 vccd1 _14394_/B sky130_fd_sc_hd__o21ai_2
XFILLER_195_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16132_ _09650_/X _16132_/A2 _16131_/X vssd1 vssd1 vccd1 vccd1 _19590_/D sky130_fd_sc_hd__o21a_1
XFILLER_154_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10556_ _11242_/A1 _14038_/A2 _10555_/X _11242_/B1 _19856_/Q vssd1 vssd1 vccd1 vccd1
+ _10556_/X sky130_fd_sc_hd__o32a_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13344_ _13334_/X _13338_/Y _13343_/Y vssd1 vssd1 vccd1 vccd1 _14296_/A sky130_fd_sc_hd__a21oi_1
XFILLER_128_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16063_ _12708_/A _16063_/A2 _13181_/B _16063_/B2 vssd1 vssd1 vccd1 vccd1 _16064_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10487_ _10485_/X _10486_/X _11259_/S vssd1 vssd1 vccd1 vccd1 _10487_/X sky130_fd_sc_hd__mux2_1
X_13275_ _13275_/A1 _19236_/Q _14794_/C1 _13274_/Y vssd1 vssd1 vccd1 vccd1 _13412_/B
+ sky130_fd_sc_hd__o211a_4
X_15014_ _15019_/A _15014_/B _15133_/B _15014_/D vssd1 vssd1 vccd1 vccd1 _15018_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_142_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12226_ _12218_/X _12219_/X _12391_/S vssd1 vssd1 vccd1 vccd1 _12226_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19822_ _20649_/CLK _19822_/D vssd1 vssd1 vccd1 vccd1 _19822_/Q sky130_fd_sc_hd__dfxtp_1
X_12157_ _12157_/A1 _17948_/A1 _12153_/X vssd1 vssd1 vccd1 vccd1 _12157_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _11106_/X _11107_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _11108_/X sky130_fd_sc_hd__mux2_1
XFILLER_257_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19753_ _20962_/CLK _19753_/D vssd1 vssd1 vccd1 vccd1 _19753_/Q sky130_fd_sc_hd__dfxtp_1
X_12088_ _12082_/X _12087_/X _12088_/S vssd1 vssd1 vccd1 vccd1 _12088_/X sky130_fd_sc_hd__mux2_1
X_16965_ _17006_/A1 _15916_/X _16945_/X _16964_/X vssd1 vssd1 vccd1 vccd1 _16965_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_238_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18704_ _18704_/A _18704_/B vssd1 vssd1 vccd1 vccd1 _20952_/D sky130_fd_sc_hd__nor2_1
X_11039_ _19401_/Q _20560_/Q _11039_/S vssd1 vssd1 vccd1 vccd1 _11039_/X sky130_fd_sc_hd__mux2_1
X_15916_ _16000_/A1 _15905_/X _15906_/X _15915_/X vssd1 vssd1 vccd1 vccd1 _15916_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_204_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19684_ _20568_/CLK _19684_/D vssd1 vssd1 vccd1 vccd1 _19684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_265_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16896_ _19978_/Q _16849_/A _16895_/Y _16896_/C1 vssd1 vssd1 vccd1 vccd1 _19978_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_264_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18635_ _20932_/Q _18686_/B vssd1 vssd1 vccd1 vccd1 _18635_/Y sky130_fd_sc_hd__nand2_1
XFILLER_252_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _14843_/S _15359_/X _15363_/X _15258_/A vssd1 vssd1 vccd1 vccd1 _15847_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18566_ _19494_/Q _18570_/B _18459_/Y _18565_/B vssd1 vssd1 vccd1 vccd1 _18566_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _20807_/Q _15941_/A2 _15771_/X _15941_/B2 _15777_/X vssd1 vssd1 vccd1 vccd1
+ _15778_/X sky130_fd_sc_hd__a221o_1
XFILLER_212_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17517_ _17525_/A1 _17516_/Y _17430_/A vssd1 vssd1 vccd1 vccd1 _20293_/D sky130_fd_sc_hd__a21oi_1
X_14729_ _19486_/Q _17944_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19486_/D sky130_fd_sc_hd__mux2_1
X_18497_ _20892_/Q _18474_/S _18496_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18498_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_590 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17448_ _20264_/Q _17446_/A _17451_/A _17443_/A vssd1 vssd1 vccd1 vccd1 _17448_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ _20238_/Q _17381_/A2 _17378_/X _18740_/A vssd1 vssd1 vccd1 vccd1 _20238_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20716_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19118_ _19511_/CLK _19118_/D vssd1 vssd1 vccd1 vccd1 _19118_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_145_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20390_ _20481_/CLK _20390_/D vssd1 vssd1 vccd1 vccd1 _20390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19049_ _21043_/Q _19049_/A2 _19048_/X _18730_/A vssd1 vssd1 vccd1 vccd1 _21043_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_204_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20645_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21011_ _21011_/CLK _21011_/D vssd1 vssd1 vccd1 vccd1 _21011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput288 _13830_/X vssd1 vssd1 vccd1 vccd1 addr0[3] sky130_fd_sc_hd__buf_4
XFILLER_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput299 _13786_/X vssd1 vssd1 vccd1 vccd1 addr1[5] sky130_fd_sc_hd__buf_4
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09704_ _09702_/X _09703_/X _11980_/S vssd1 vssd1 vccd1 vccd1 _09704_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09635_ _09589_/X _09610_/C _09634_/X _09686_/A vssd1 vssd1 vccd1 vccd1 _09636_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09566_ _09567_/A _19154_/Q _12579_/C vssd1 vssd1 vccd1 vccd1 _15303_/A sky130_fd_sc_hd__nor3b_4
XFILLER_270_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09497_ _19226_/Q vssd1 vssd1 vccd1 vccd1 _09497_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20726_ _20759_/CLK _20726_/D vssd1 vssd1 vccd1 vccd1 _20726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20657_ _20657_/CLK _20657_/D vssd1 vssd1 vccd1 vccd1 _20657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10410_ _11290_/A _19908_/Q _11292_/S0 _20033_/Q vssd1 vssd1 vccd1 vccd1 _10410_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _11391_/A _20501_/Q _12346_/S _20533_/Q vssd1 vssd1 vccd1 vccd1 _11390_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_176_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20588_ _20694_/CLK _20588_/D vssd1 vssd1 vccd1 vccd1 _20588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10341_ _10356_/A _19348_/Q _20703_/Q _10518_/S _11304_/S vssd1 vssd1 vccd1 vccd1
+ _10341_/X sky130_fd_sc_hd__a221o_1
XFILLER_152_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13060_ _20948_/Q _20882_/Q _13060_/C _13060_/D vssd1 vssd1 vccd1 vccd1 _13505_/A
+ sky130_fd_sc_hd__and4_1
X_10272_ _10260_/X _10271_/X _12275_/A vssd1 vssd1 vccd1 vccd1 _10272_/X sky130_fd_sc_hd__mux2_4
XFILLER_3_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12011_ _12009_/X _12010_/X _12011_/S vssd1 vssd1 vccd1 vccd1 _12011_/X sky130_fd_sc_hd__mux2_1
Xfanout1403 _09736_/Y vssd1 vssd1 vccd1 vccd1 _12081_/S0 sky130_fd_sc_hd__buf_6
XFILLER_239_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1414 fanout1430/X vssd1 vssd1 vccd1 vccd1 _11203_/S sky130_fd_sc_hd__buf_6
Xfanout1425 fanout1430/X vssd1 vssd1 vccd1 vccd1 _11393_/S0 sky130_fd_sc_hd__buf_4
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1436 _11852_/B2 vssd1 vssd1 vccd1 vccd1 _12085_/B2 sky130_fd_sc_hd__buf_8
XFILLER_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1447 _10405_/C vssd1 vssd1 vccd1 vccd1 _09834_/C sky130_fd_sc_hd__buf_6
Xfanout1458 _11391_/C vssd1 vssd1 vccd1 vccd1 _12254_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_47_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1469 _10630_/C1 vssd1 vssd1 vccd1 vccd1 _12091_/S sky130_fd_sc_hd__buf_8
X_16750_ _16799_/S _09520_/Y _16726_/X _16749_/Y vssd1 vssd1 vccd1 vccd1 _16750_/X
+ sky130_fd_sc_hd__o211a_4
X_13962_ _19154_/Q _19050_/S _14043_/B1 _13961_/X _14458_/A vssd1 vssd1 vccd1 vccd1
+ _19154_/D sky130_fd_sc_hd__o221a_1
Xfanout493 _17885_/X vssd1 vssd1 vccd1 vccd1 _17912_/S sky130_fd_sc_hd__buf_6
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _16024_/A1 _15699_/X _15700_/Y _13427_/A _15975_/B2 vssd1 vssd1 vccd1 vccd1
+ _15701_/X sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_79_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19560_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12913_ _13106_/A _13106_/B _13106_/C _13106_/D vssd1 vssd1 vccd1 vccd1 _12913_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16681_ _19936_/Q _17859_/A1 _16704_/S vssd1 vssd1 vccd1 vccd1 _19936_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13893_ _19111_/Q _14527_/A2 _13896_/B1 _12519_/A _14458_/A vssd1 vssd1 vccd1 vccd1
+ _19111_/D sky130_fd_sc_hd__o221a_1
XFILLER_74_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18420_ _18708_/A _18420_/B vssd1 vssd1 vccd1 vccd1 _20864_/D sky130_fd_sc_hd__and2_1
X_15632_ _20738_/Q _16041_/A2 _16041_/B1 _20770_/Q vssd1 vssd1 vccd1 vccd1 _15632_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_250_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _19510_/Q _12855_/B _19511_/Q vssd1 vssd1 vccd1 vccd1 _12845_/B sky130_fd_sc_hd__a21oi_1
XFILLER_15_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _18505_/B _18363_/B vssd1 vssd1 vccd1 vccd1 _18351_/Y sky130_fd_sc_hd__nand2_1
X_15563_ _19716_/Q _15595_/A2 _15595_/B1 _19748_/Q vssd1 vssd1 vccd1 vccd1 _15563_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _15380_/A _12784_/B vssd1 vssd1 vccd1 vccd1 _12775_/Y sky130_fd_sc_hd__nand2_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17302_/A _17329_/S _17302_/C vssd1 vssd1 vccd1 vccd1 _17302_/X sky130_fd_sc_hd__and3_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14514_ _19292_/Q _17945_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19292_/D sky130_fd_sc_hd__mux2_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _18730_/A _18282_/B vssd1 vssd1 vccd1 vccd1 _20810_/D sky130_fd_sc_hd__and2_1
X_11726_ _19512_/Q _11725_/Y _11726_/S vssd1 vssd1 vccd1 vccd1 _11733_/B sky130_fd_sc_hd__mux2_4
XFILLER_187_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _15494_/A _15494_/B vssd1 vssd1 vccd1 vccd1 _15494_/X sky130_fd_sc_hd__or2_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17233_ _17235_/A _17336_/B vssd1 vssd1 vccd1 vccd1 _17233_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14445_ _20218_/Q _19247_/Q _14477_/S vssd1 vssd1 vccd1 vccd1 _14446_/B sky130_fd_sc_hd__mux2_1
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11657_ _20575_/Q _12044_/B _11656_/X _12051_/C1 vssd1 vssd1 vccd1 vccd1 _11657_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10608_ _10602_/X _10603_/X _10604_/X _10607_/X _12088_/S vssd1 vssd1 vccd1 vccd1
+ _10608_/X sky130_fd_sc_hd__a311o_1
X_17164_ _20130_/Q _17689_/A1 _17166_/S vssd1 vssd1 vccd1 vccd1 _20130_/D sky130_fd_sc_hd__mux2_1
X_14376_ _14376_/A _14376_/B vssd1 vssd1 vccd1 vccd1 _14376_/Y sky130_fd_sc_hd__xnor2_1
X_11588_ _20137_/Q _20105_/Q _11979_/S vssd1 vssd1 vccd1 vccd1 _11588_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16115_ _09672_/X _09673_/X _16131_/A2 vssd1 vssd1 vccd1 vccd1 _16115_/X sky130_fd_sc_hd__a21bo_1
XFILLER_116_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _13327_/A _13327_/B vssd1 vssd1 vccd1 vccd1 _13328_/B sky130_fd_sc_hd__xnor2_1
XFILLER_127_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10539_ _12581_/A _15443_/A _10509_/Y vssd1 vssd1 vccd1 vccd1 _10641_/B sky130_fd_sc_hd__o21ba_4
X_17095_ _20065_/Q _17095_/A1 _17111_/S vssd1 vssd1 vccd1 vccd1 _20065_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16046_ _16046_/A1 _16045_/X _16042_/X vssd1 vssd1 vccd1 vccd1 _16046_/X sky130_fd_sc_hd__o21a_4
X_13258_ _13258_/A _13258_/B _13258_/C vssd1 vssd1 vccd1 vccd1 _13258_/X sky130_fd_sc_hd__and3_1
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12209_ _12366_/A1 _10124_/B _10037_/B vssd1 vssd1 vccd1 vccd1 _12209_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13189_ _15954_/A _13189_/B vssd1 vssd1 vccd1 vccd1 _17041_/B sky130_fd_sc_hd__nand2_8
XFILLER_285_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19805_ _20467_/CLK _19805_/D vssd1 vssd1 vccd1 vccd1 _19805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17997_ _20737_/Q _20736_/Q _17997_/C vssd1 vssd1 vccd1 vccd1 _18003_/C sky130_fd_sc_hd__and3_2
XFILLER_229_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19736_ _20725_/CLK _19736_/D vssd1 vssd1 vccd1 vccd1 _19736_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1970 _13595_/A vssd1 vssd1 vccd1 vccd1 _16241_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16948_ _16981_/A1 _15861_/X _16945_/X _16947_/X vssd1 vssd1 vccd1 vccd1 _16948_/X
+ sky130_fd_sc_hd__o211a_2
Xfanout1981 _18814_/A vssd1 vssd1 vccd1 vccd1 _18821_/A sky130_fd_sc_hd__buf_6
XFILLER_238_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1992 _18056_/A vssd1 vssd1 vccd1 vccd1 _18064_/A sky130_fd_sc_hd__buf_4
XFILLER_253_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19667_ _20155_/CLK _19667_/D vssd1 vssd1 vccd1 vccd1 _19667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16879_ _20623_/Q _16945_/B _16945_/C vssd1 vssd1 vccd1 vccd1 _16879_/X sky130_fd_sc_hd__and3_4
XFILLER_64_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18618_ _18856_/A _18618_/B vssd1 vssd1 vccd1 vccd1 _20927_/D sky130_fd_sc_hd__nor2_1
XFILLER_252_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19598_ _19606_/CLK _19598_/D vssd1 vssd1 vccd1 vccd1 _19598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18549_ _18980_/A _18549_/B vssd1 vssd1 vccd1 vccd1 _20909_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20511_ _20675_/CLK _20511_/D vssd1 vssd1 vccd1 vccd1 _20511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20442_ _20557_/CLK _20442_/D vssd1 vssd1 vccd1 vccd1 _20442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20373_ _20718_/CLK _20373_/D vssd1 vssd1 vccd1 vccd1 _20373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09618_ _09618_/A _10979_/C vssd1 vssd1 vccd1 vccd1 _09618_/Y sky130_fd_sc_hd__nand2_8
XFILLER_284_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ input151/X input136/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10890_/X sky130_fd_sc_hd__mux2_8
XFILLER_271_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09549_ _19153_/Q _19152_/Q _09734_/B _12490_/B vssd1 vssd1 vccd1 vccd1 _12574_/A
+ sky130_fd_sc_hd__or4_4
XPHY_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12560_ _13636_/A _13694_/A vssd1 vssd1 vccd1 vccd1 _13143_/B sky130_fd_sc_hd__nor2_4
XFILLER_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11511_ _11509_/X _11510_/X _11902_/S vssd1 vssd1 vccd1 vccd1 _11511_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20709_ _20713_/CLK _20709_/D vssd1 vssd1 vccd1 vccd1 _20709_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_197_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20353_/CLK sky130_fd_sc_hd__clkbuf_16
X_12491_ _19158_/Q _12479_/A _12657_/A2 _16005_/A1 _12584_/C vssd1 vssd1 vccd1 vccd1
+ _12496_/A sky130_fd_sc_hd__a32o_2
XFILLER_8_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14230_ _14240_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14232_/B sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_126_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20621_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_11442_ _12143_/S _11441_/X _11440_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _11442_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11373_ _19670_/Q _20158_/Q _11377_/S vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__mux2_1
X_14161_ _14161_/A _14161_/B vssd1 vssd1 vccd1 vccd1 _14162_/B sky130_fd_sc_hd__or2_2
XFILLER_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10324_ _19281_/Q _20068_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10324_/X sky130_fd_sc_hd__mux2_1
X_13112_ _09488_/A _19245_/Q _16191_/A _13111_/Y vssd1 vssd1 vccd1 vccd1 _13112_/X
+ sky130_fd_sc_hd__o211a_2
X_14092_ _19205_/Q _14104_/A2 _14091_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1 _19205_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10255_ _20316_/Q _11379_/B vssd1 vssd1 vccd1 vccd1 _10255_/X sky130_fd_sc_hd__or2_1
X_17920_ _20689_/Q _17920_/A1 _17934_/S vssd1 vssd1 vccd1 vccd1 _20689_/D sky130_fd_sc_hd__mux2_1
X_13043_ _20956_/Q _20890_/Q vssd1 vssd1 vccd1 vccd1 _13043_/Y sky130_fd_sc_hd__nor2_2
XFILLER_285_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1200 _17324_/C1 vssd1 vssd1 vccd1 vccd1 _17291_/B1 sky130_fd_sc_hd__buf_4
XFILLER_266_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1211 _16002_/A1 vssd1 vssd1 vccd1 vccd1 _15283_/A sky130_fd_sc_hd__buf_4
XFILLER_267_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17851_ _17851_/A _17851_/B _17851_/C vssd1 vssd1 vccd1 vccd1 _17851_/X sky130_fd_sc_hd__and3_4
X_10186_ _10184_/X _10185_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _10186_/X sky130_fd_sc_hd__mux2_1
Xfanout1222 _13305_/B vssd1 vssd1 vccd1 vccd1 _13355_/B sky130_fd_sc_hd__buf_4
Xfanout1233 _11230_/A vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__buf_4
XFILLER_278_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1244 _17370_/B1 vssd1 vssd1 vccd1 vccd1 _17362_/B1 sky130_fd_sc_hd__buf_6
XFILLER_266_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16802_ _16798_/Y _16801_/X _17011_/B1 vssd1 vssd1 vccd1 vccd1 _16802_/Y sky130_fd_sc_hd__a21oi_4
Xfanout1255 _16716_/A vssd1 vssd1 vccd1 vccd1 _16945_/B sky130_fd_sc_hd__buf_6
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17782_ _20559_/Q _17782_/A1 _17794_/S vssd1 vssd1 vccd1 vccd1 _20559_/D sky130_fd_sc_hd__mux2_1
Xfanout1266 _09689_/X vssd1 vssd1 vccd1 vccd1 _13675_/A sky130_fd_sc_hd__clkbuf_16
X_14994_ _15019_/A _15021_/B vssd1 vssd1 vccd1 vccd1 _15022_/D sky130_fd_sc_hd__nand2_4
Xfanout1277 _16034_/S vssd1 vssd1 vccd1 vccd1 _15949_/A sky130_fd_sc_hd__buf_4
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1288 _12581_/A vssd1 vssd1 vccd1 vccd1 _15150_/C1 sky130_fd_sc_hd__buf_4
XFILLER_266_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1299 _14117_/Y vssd1 vssd1 vccd1 vccd1 _14330_/B1 sky130_fd_sc_hd__buf_6
X_16733_ _20398_/Q _17004_/A2 _17004_/B1 vssd1 vssd1 vccd1 vccd1 _16733_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19521_ _19523_/CLK _19521_/D vssd1 vssd1 vccd1 vccd1 _19521_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_281_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13945_ _19147_/Q _13941_/B _13946_/B1 _13112_/X vssd1 vssd1 vccd1 vccd1 _19147_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19452_ _20451_/CLK _19452_/D vssd1 vssd1 vccd1 vccd1 _19452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16664_ _19921_/Q _17910_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19921_/D sky130_fd_sc_hd__mux2_1
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13876_ _19094_/Q _13953_/A2 _13881_/B1 _19160_/Q _15288_/C1 vssd1 vssd1 vccd1 vccd1
+ _19094_/D sky130_fd_sc_hd__o221a_1
XFILLER_250_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18403_ _20856_/Q _18190_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18404_/B sky130_fd_sc_hd__mux2_1
X_15615_ _14815_/S _15610_/Y _15626_/B _15468_/A vssd1 vssd1 vccd1 vccd1 _15615_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_216_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19383_ _20646_/CLK _19383_/D vssd1 vssd1 vccd1 vccd1 _19383_/Q sky130_fd_sc_hd__dfxtp_1
X_12827_ _19513_/Q _12857_/B vssd1 vssd1 vccd1 vccd1 _12829_/C sky130_fd_sc_hd__nor2_2
X_16595_ _16595_/A vssd1 vssd1 vccd1 vccd1 _16595_/Y sky130_fd_sc_hd__inv_2
XFILLER_250_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18334_ _20822_/Q _18341_/B _18333_/Y _18700_/A vssd1 vssd1 vccd1 vccd1 _20822_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15546_ _14841_/S _15254_/X _15066_/S vssd1 vssd1 vccd1 vccd1 _15546_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _19505_/Q _12758_/B vssd1 vssd1 vccd1 vccd1 _12758_/X sky130_fd_sc_hd__and2_1
XFILLER_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18265_ _18529_/B vssd1 vssd1 vccd1 vccd1 _18265_/Y sky130_fd_sc_hd__inv_2
X_11709_ _19416_/Q _12025_/S _11708_/X _09834_/C vssd1 vssd1 vccd1 vccd1 _11709_/X
+ sky130_fd_sc_hd__o211a_1
X_15477_ _21023_/Q _20991_/Q _15508_/S vssd1 vssd1 vccd1 vccd1 _15477_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12689_ _12653_/A _12653_/B _12653_/C vssd1 vssd1 vccd1 vccd1 _12692_/D sky130_fd_sc_hd__o21a_1
X_17216_ _20180_/Q _17950_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20180_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14428_ _14427_/A _14423_/B _14427_/Y _09488_/A vssd1 vssd1 vccd1 vccd1 _14428_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18196_ _20793_/Q _18195_/Y _18311_/S vssd1 vssd1 vccd1 vccd1 _18197_/B sky130_fd_sc_hd__mux2_1
XFILLER_163_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17147_ _20115_/Q _17949_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20115_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14359_ _14437_/A _14437_/B _14359_/C vssd1 vssd1 vccd1 vccd1 _14359_/X sky130_fd_sc_hd__or3_1
XFILLER_183_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17078_ _20050_/Q _17112_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20050_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16029_ _13181_/A _15982_/C _16056_/B1 _16028_/X vssd1 vssd1 vccd1 vccd1 _16029_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_276_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19719_ _20268_/CLK _19719_/D vssd1 vssd1 vccd1 vccd1 _19719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20991_ _21023_/CLK _20991_/D vssd1 vssd1 vccd1 vccd1 _20991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20425_ _20425_/CLK _20425_/D vssd1 vssd1 vccd1 vccd1 _20425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20356_ _20706_/CLK _20356_/D vssd1 vssd1 vccd1 vccd1 _20356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20287_ _21010_/CLK _20287_/D vssd1 vssd1 vccd1 vccd1 _20287_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10040_ _19587_/Q _10039_/X _11243_/S vssd1 vssd1 vccd1 vccd1 _10041_/B sky130_fd_sc_hd__mux2_2
XFILLER_276_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11991_ _19825_/Q _19329_/Q _11994_/S vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13730_ _13730_/A _13730_/B vssd1 vssd1 vccd1 vccd1 _13772_/B sky130_fd_sc_hd__or2_2
XFILLER_217_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10942_ _11290_/A _20661_/Q _11290_/C vssd1 vssd1 vccd1 vccd1 _10942_/X sky130_fd_sc_hd__or3_1
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ _13661_/A _13661_/B vssd1 vssd1 vccd1 vccd1 _13662_/A sky130_fd_sc_hd__nand2_2
XFILLER_32_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10873_ _11391_/A _20123_/Q _20091_/Q _12344_/S vssd1 vssd1 vccd1 vccd1 _10873_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15400_ _15520_/B2 _15378_/X _15379_/Y _15399_/X vssd1 vssd1 vccd1 vccd1 _15400_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_188_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _19520_/Q _19519_/Q _12884_/B vssd1 vssd1 vccd1 vccd1 _12889_/A sky130_fd_sc_hd__and3_1
X_16380_ _19738_/Q _16380_/B vssd1 vssd1 vccd1 vccd1 _16386_/C sky130_fd_sc_hd__and2_2
XFILLER_169_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13591_/Y _20955_/Q _13607_/B vssd1 vssd1 vccd1 vccd1 _13592_/X sky130_fd_sc_hd__mux2_2
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15331_ _15331_/A _16009_/B vssd1 vssd1 vccd1 vccd1 _15331_/Y sky130_fd_sc_hd__nand2_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12543_ _20866_/Q _12548_/B _12543_/C vssd1 vssd1 vccd1 vccd1 _12551_/C sky130_fd_sc_hd__and3_4
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18050_ _20756_/Q _18053_/C _18054_/A vssd1 vssd1 vccd1 vccd1 _18050_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15262_ _15066_/S _15261_/X _15548_/B1 vssd1 vssd1 vccd1 vccd1 _15262_/Y sky130_fd_sc_hd__o21ai_2
X_12474_ _14894_/A _14898_/A vssd1 vssd1 vccd1 vccd1 _12474_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17001_ _16998_/Y _17000_/Y _17011_/B1 vssd1 vssd1 vccd1 vccd1 _17001_/Y sky130_fd_sc_hd__a21oi_4
X_14213_ _14524_/A1 _14212_/X _13593_/X vssd1 vssd1 vccd1 vccd1 _14214_/C sky130_fd_sc_hd__a21o_1
X_11425_ _11514_/A1 _20706_/Q _12124_/S _11424_/X vssd1 vssd1 vccd1 vccd1 _11425_/X
+ sky130_fd_sc_hd__a31o_1
X_15193_ _20885_/Q _14971_/A _15566_/B1 _15192_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15193_/X sky130_fd_sc_hd__a221o_1
XFILLER_172_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _16804_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14144_ _14255_/A _14204_/B _14144_/C vssd1 vssd1 vccd1 vccd1 _14144_/X sky130_fd_sc_hd__or3_1
XFILLER_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11356_ _11359_/S _11355_/X _11354_/X _11363_/A1 vssd1 vssd1 vccd1 vccd1 _11356_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _10302_/X _10303_/X _11256_/S vssd1 vssd1 vccd1 vccd1 _10307_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14075_ _14107_/A _14107_/B _14075_/C vssd1 vssd1 vccd1 vccd1 _14075_/X sky130_fd_sc_hd__or3_1
XFILLER_180_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18952_ _18547_/X _18978_/B _18950_/X _18951_/Y vssd1 vssd1 vccd1 vccd1 _18953_/B
+ sky130_fd_sc_hd__o211a_1
X_11287_ _19623_/Q _19929_/Q _19267_/Q _20054_/Q _11292_/S0 _11290_/C vssd1 vssd1
+ vccd1 vccd1 _11287_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_94_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20688_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_140_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17903_ _20674_/Q _17903_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20674_/D sky130_fd_sc_hd__mux2_1
X_13026_ _20966_/Q _20900_/Q vssd1 vssd1 vccd1 vccd1 _13367_/B sky130_fd_sc_hd__nand2_2
X_10238_ _11170_/B1 _10237_/X _10236_/X _09688_/A vssd1 vssd1 vccd1 vccd1 _10238_/X
+ sky130_fd_sc_hd__a211o_1
X_18883_ _18517_/X _18978_/B _18881_/X _18882_/Y vssd1 vssd1 vccd1 vccd1 _18884_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_239_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1030 _15527_/Y vssd1 vssd1 vccd1 vccd1 _15544_/A sky130_fd_sc_hd__buf_2
XFILLER_239_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1041 _17887_/A1 vssd1 vssd1 vccd1 vccd1 _17921_/A1 sky130_fd_sc_hd__buf_8
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_23_wb_clk_i _20408_/CLK vssd1 vssd1 vccd1 vccd1 _20683_/CLK sky130_fd_sc_hd__clkbuf_16
X_10169_ _20131_/Q _20099_/Q _12428_/S vssd1 vssd1 vccd1 vccd1 _10169_/X sky130_fd_sc_hd__mux2_1
Xfanout1052 _10978_/X vssd1 vssd1 vccd1 vccd1 _11049_/B1 sky130_fd_sc_hd__buf_4
X_17834_ _20609_/Q _17906_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20609_/D sky130_fd_sc_hd__mux2_1
XFILLER_266_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1063 _10728_/X vssd1 vssd1 vccd1 vccd1 _17892_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_227_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1074 _17885_/B vssd1 vssd1 vccd1 vccd1 _17919_/B sky130_fd_sc_hd__buf_2
XFILLER_254_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1085 _17950_/A1 vssd1 vssd1 vccd1 vccd1 _17114_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_48_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1096 _17914_/A1 vssd1 vssd1 vccd1 vccd1 _17705_/A1 sky130_fd_sc_hd__buf_4
X_14977_ _14978_/B vssd1 vssd1 vccd1 vccd1 _14977_/Y sky130_fd_sc_hd__inv_2
X_17765_ _20544_/Q _17871_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20544_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19504_ _19506_/CLK _19504_/D vssd1 vssd1 vccd1 vccd1 _19504_/Q sky130_fd_sc_hd__dfxtp_4
X_16716_ _16716_/A _16716_/B vssd1 vssd1 vccd1 vccd1 _16716_/Y sky130_fd_sc_hd__nand2_1
X_13928_ _19132_/Q _13906_/B _13932_/B1 _13411_/B vssd1 vssd1 vccd1 vccd1 _19132_/D
+ sky130_fd_sc_hd__o22a_1
X_17696_ _20480_/Q _17696_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20480_/D sky130_fd_sc_hd__mux2_1
XFILLER_235_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16647_ _19904_/Q _17684_/A1 _16670_/S vssd1 vssd1 vccd1 vccd1 _19904_/D sky130_fd_sc_hd__mux2_1
X_19435_ _20687_/CLK _19435_/D vssd1 vssd1 vccd1 vccd1 _19435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_262_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13859_ _13860_/B _13860_/C vssd1 vssd1 vccd1 vccd1 _16068_/A sky130_fd_sc_hd__or2_4
XFILLER_211_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16578_ _19855_/Q _16578_/A2 _16578_/B1 input26/X vssd1 vssd1 vccd1 vccd1 _16579_/B
+ sky130_fd_sc_hd__o22a_1
X_19366_ _20657_/CLK _19366_/D vssd1 vssd1 vccd1 vccd1 _19366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18317_ _18985_/A _18317_/B vssd1 vssd1 vccd1 vccd1 _20817_/D sky130_fd_sc_hd__and2_1
X_15529_ _16002_/A1 _15528_/Y _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15529_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19297_ _20084_/CLK _19297_/D vssd1 vssd1 vccd1 vccd1 _19297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18248_ _19545_/Q _18248_/B vssd1 vssd1 vccd1 vccd1 _18248_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_136_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18179_ _18163_/A _14158_/B _18178_/Y vssd1 vssd1 vccd1 vccd1 _18477_/B sky130_fd_sc_hd__o21ai_4
XFILLER_144_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20210_ _20766_/CLK _20210_/D vssd1 vssd1 vccd1 vccd1 _20210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20141_ _20712_/CLK _20141_/D vssd1 vssd1 vccd1 vccd1 _20141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09952_ _20577_/Q _11897_/B _09951_/X _11892_/C1 vssd1 vssd1 vccd1 vccd1 _09952_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20072_ _20679_/CLK _20072_/D vssd1 vssd1 vccd1 vccd1 _20072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _20139_/Q _20107_/Q _11527_/S vssd1 vssd1 vccd1 vccd1 _09883_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_408 _17574_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_419 _09624_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20974_ _21040_/CLK _20974_/D vssd1 vssd1 vccd1 vccd1 _20974_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_272_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11210_ _11191_/A _19463_/Q _19431_/Q _11211_/S vssd1 vssd1 vccd1 vccd1 _11210_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12190_ _11849_/S _12187_/X _12189_/X _12190_/C1 vssd1 vssd1 vccd1 vccd1 _12190_/X
+ sky130_fd_sc_hd__o211a_1
X_20408_ _20408_/CLK _20408_/D vssd1 vssd1 vccd1 vccd1 _20408_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ input118/X input133/X _11241_/S vssd1 vssd1 vccd1 vccd1 _11141_/X sky130_fd_sc_hd__mux2_8
X_20339_ _20426_/CLK _20339_/D vssd1 vssd1 vccd1 vccd1 _20339_/Q sky130_fd_sc_hd__dfxtp_1
X_11072_ _19931_/Q _12213_/B vssd1 vssd1 vccd1 vccd1 _11072_/X sky130_fd_sc_hd__or2_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput100 dout0[61] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput111 dout1[13] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput122 dout1[23] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_hd__clkbuf_2
X_10023_ _10284_/A _11234_/B split7/A vssd1 vssd1 vccd1 vccd1 _11326_/B sky130_fd_sc_hd__o21ai_2
X_14900_ _16945_/C _17219_/A _18134_/A vssd1 vssd1 vccd1 vccd1 _16720_/D sky130_fd_sc_hd__a21o_2
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput133 dout1[33] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_hd__buf_2
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _20811_/Q _15941_/A2 _15873_/X _15941_/B2 _15879_/X vssd1 vssd1 vccd1 vccd1
+ _15880_/X sky130_fd_sc_hd__a221o_2
XFILLER_264_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput144 dout1[43] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput155 dout1[53] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__clkbuf_2
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 dout1[63] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_hd__buf_2
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput177 irq[15] vssd1 vssd1 vccd1 vccd1 _12547_/C sky130_fd_sc_hd__clkbuf_2
X_14831_ _14829_/X _14830_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _14831_/X sky130_fd_sc_hd__mux2_1
XFILLER_248_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 jtag_tdi vssd1 vssd1 vccd1 vccd1 _17236_/A sky130_fd_sc_hd__buf_12
Xinput199 localMemory_wb_adr_i[18] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__clkbuf_2
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _20310_/Q _17686_/A1 _17567_/S vssd1 vssd1 vccd1 vccd1 _20310_/D sky130_fd_sc_hd__mux2_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14762_ _19128_/Q _14764_/A2 _14761_/X _18352_/C1 vssd1 vssd1 vccd1 vccd1 _19505_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ _19892_/Q _11979_/S vssd1 vssd1 vccd1 vccd1 _11974_/X sky130_fd_sc_hd__or2_1
XFILLER_251_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16501_ _19808_/Q _17060_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19808_/D sky130_fd_sc_hd__mux2_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _13685_/A _13676_/B _13675_/Y _13655_/A vssd1 vssd1 vccd1 vccd1 _13713_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_17481_ _17487_/A1 _17480_/Y _18704_/A vssd1 vssd1 vccd1 vccd1 _20275_/D sky130_fd_sc_hd__a21oi_1
X_10925_ _11008_/A1 _19466_/Q _19434_/Q _10924_/S _11338_/A1 vssd1 vssd1 vccd1 vccd1
+ _10925_/X sky130_fd_sc_hd__a221o_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14693_ _19452_/Q _17802_/A1 _14699_/S vssd1 vssd1 vccd1 vccd1 _19452_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19220_ _19223_/CLK _19220_/D vssd1 vssd1 vccd1 vccd1 _19220_/Q sky130_fd_sc_hd__dfxtp_4
X_16432_ _19757_/Q _16434_/C _16431_/Y vssd1 vssd1 vccd1 vccd1 _19757_/D sky130_fd_sc_hd__o21a_1
XFILLER_204_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13644_ _13657_/A _13644_/B vssd1 vssd1 vccd1 vccd1 _13708_/B sky130_fd_sc_hd__nor2_8
Xclkbuf_leaf_141_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19696_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10856_ _10854_/X _10855_/X _12414_/S vssd1 vssd1 vccd1 vccd1 _10856_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19151_ _19620_/CLK _19151_/D vssd1 vssd1 vccd1 vccd1 _19151_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _18821_/A _16363_/B _16364_/B vssd1 vssd1 vccd1 vccd1 _19731_/D sky130_fd_sc_hd__nor3_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13587_/B _13575_/B _13575_/C vssd1 vssd1 vccd1 vccd1 _13575_/X sky130_fd_sc_hd__and3b_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _19668_/Q _11126_/B _12419_/C1 vssd1 vssd1 vccd1 vccd1 _10787_/X sky130_fd_sc_hd__o21a_1
X_18102_ _18104_/A _18102_/B _18103_/B vssd1 vssd1 vccd1 vccd1 _20775_/D sky130_fd_sc_hd__nor3_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _20979_/Q _15314_/B _15314_/C _15314_/D vssd1 vssd1 vccd1 vccd1 _15314_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_158_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19082_ _20427_/Q vssd1 vssd1 vccd1 vccd1 _20427_/D sky130_fd_sc_hd__clkbuf_2
X_12526_ _13350_/A _13107_/B vssd1 vssd1 vccd1 vccd1 _14110_/B sky130_fd_sc_hd__or2_4
X_16294_ _19705_/Q _19706_/Q _16294_/C vssd1 vssd1 vccd1 vccd1 _16300_/C sky130_fd_sc_hd__and3_2
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18033_ _20750_/Q _18036_/C vssd1 vssd1 vccd1 vccd1 _18034_/B sky130_fd_sc_hd__and2_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _15026_/Y _15229_/X _15673_/B1 vssd1 vssd1 vccd1 vccd1 _15246_/C sky130_fd_sc_hd__o21a_1
XFILLER_172_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12457_ _14895_/A _12464_/C vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__nand2_2
X_11408_ _10456_/Y _10641_/A _10641_/B _10640_/X _11407_/X vssd1 vssd1 vccd1 vccd1
+ _11408_/X sky130_fd_sc_hd__a311o_1
XFILLER_126_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15176_ _15611_/S _15172_/X _15174_/X _15175_/Y _15610_/A1 vssd1 vssd1 vccd1 vccd1
+ _15176_/X sky130_fd_sc_hd__a311o_1
X_12388_ _11094_/S _12387_/X _12386_/X _12398_/C1 vssd1 vssd1 vccd1 vccd1 _12388_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14127_ _19215_/Q _14205_/A2 _14126_/X _18698_/A vssd1 vssd1 vccd1 vccd1 _19215_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11339_ _19406_/Q _20565_/Q _11342_/S vssd1 vssd1 vccd1 vccd1 _11339_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19984_ _20862_/CLK _19984_/D vssd1 vssd1 vccd1 vccd1 _19984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14058_ _19188_/Q _14108_/A2 _14057_/X _14458_/A vssd1 vssd1 vccd1 vccd1 _19188_/D
+ sky130_fd_sc_hd__o211a_1
X_18935_ _19142_/Q _18976_/A2 _18767_/B vssd1 vssd1 vccd1 vccd1 _18935_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13009_ _20974_/Q _20908_/Q vssd1 vssd1 vccd1 vccd1 _13009_/Y sky130_fd_sc_hd__nor2_1
XFILLER_268_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18866_ _19132_/Q _12533_/B _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18866_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_283_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17817_ _20592_/Q _17889_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20592_/D sky130_fd_sc_hd__mux2_1
XFILLER_282_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18797_ _09493_/Y _18796_/X _18968_/A vssd1 vssd1 vccd1 vccd1 _18797_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17748_ _20527_/Q _17888_/A1 _17776_/S vssd1 vssd1 vccd1 vccd1 _20527_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17679_ _20463_/Q _17679_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20463_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19418_ _20714_/CLK _19418_/D vssd1 vssd1 vccd1 vccd1 _19418_/Q sky130_fd_sc_hd__dfxtp_1
X_20690_ _20690_/CLK _20690_/D vssd1 vssd1 vccd1 vccd1 _20690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19349_ _20704_/CLK _19349_/D vssd1 vssd1 vccd1 vccd1 _19349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20124_ _20563_/CLK _20124_/D vssd1 vssd1 vccd1 vccd1 _20124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout801 _12476_/X vssd1 vssd1 vccd1 vccd1 _12479_/A sky130_fd_sc_hd__buf_6
X_09935_ _09926_/X _09934_/Y _09839_/A _09918_/X vssd1 vssd1 vccd1 vccd1 _09935_/X
+ sky130_fd_sc_hd__o2bb2a_2
Xfanout812 _13776_/B1 vssd1 vssd1 vccd1 vccd1 _13663_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_132_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout823 _15017_/Y vssd1 vssd1 vccd1 vccd1 _15323_/B sky130_fd_sc_hd__buf_6
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout834 _18749_/S vssd1 vssd1 vccd1 vccd1 _18753_/S sky130_fd_sc_hd__buf_6
XFILLER_113_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout845 _18357_/B vssd1 vssd1 vccd1 vccd1 _18363_/B sky130_fd_sc_hd__clkbuf_8
Xfanout856 _15998_/A2 vssd1 vssd1 vccd1 vccd1 _16047_/A2 sky130_fd_sc_hd__buf_6
X_20055_ _20694_/CLK _20055_/D vssd1 vssd1 vccd1 vccd1 _20055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09866_ input120/X input155/X _11241_/S vssd1 vssd1 vccd1 vccd1 _09866_/X sky130_fd_sc_hd__mux2_8
XFILLER_219_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout867 _15309_/S vssd1 vssd1 vccd1 vccd1 _15993_/S sky130_fd_sc_hd__buf_8
XFILLER_131_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout878 _15933_/B vssd1 vssd1 vccd1 vccd1 _15990_/B sky130_fd_sc_hd__clkbuf_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout889 _18563_/X vssd1 vssd1 vccd1 vccd1 _18688_/A2 sky130_fd_sc_hd__buf_4
XFILLER_133_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09797_ _10430_/S _12060_/A1 _19356_/Q _12046_/B1 vssd1 vssd1 vccd1 vccd1 _09797_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_280_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 _19840_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_216 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_227 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_238 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20957_ _21023_/CLK _20957_/D vssd1 vssd1 vccd1 vccd1 _20957_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _19405_/Q _20564_/Q _12417_/S vssd1 vssd1 vccd1 vccd1 _10710_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _13670_/A1 _17904_/A1 _11686_/X _12075_/C1 vssd1 vssd1 vccd1 vccd1 _13712_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_202_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20888_ _20949_/CLK _20888_/D vssd1 vssd1 vccd1 vccd1 _20888_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ _10641_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__nand2_1
XFILLER_139_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13360_ _14776_/C1 _13345_/X _13359_/A vssd1 vssd1 vccd1 vccd1 _13361_/D sky130_fd_sc_hd__a21bo_1
XFILLER_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10572_ _19874_/Q _11676_/S _10571_/X _12051_/C1 vssd1 vssd1 vccd1 vccd1 _10572_/X
+ sky130_fd_sc_hd__o211a_1
X_12311_ _12311_/A1 _12302_/X _12310_/X _12311_/C1 vssd1 vssd1 vccd1 vccd1 _12311_/X
+ sky130_fd_sc_hd__a211o_2
X_13291_ _13290_/A _13290_/B _13290_/C vssd1 vssd1 vccd1 vccd1 _13291_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15030_ _15520_/B2 _14893_/X _15029_/X _16005_/A1 vssd1 vssd1 vccd1 vccd1 _15030_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12242_ _12314_/C1 _12241_/X _12238_/X _12399_/C1 vssd1 vssd1 vccd1 vccd1 _12242_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12173_ _19690_/Q _20178_/Q _12174_/S vssd1 vssd1 vccd1 vccd1 _12173_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ _19400_/Q _20559_/Q _11126_/B vssd1 vssd1 vccd1 vccd1 _11124_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16981_ _16981_/A1 _15972_/X _16945_/X _16980_/X vssd1 vssd1 vccd1 vccd1 _16981_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_77_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18720_ _18720_/A _18720_/B vssd1 vssd1 vccd1 vccd1 _20960_/D sky130_fd_sc_hd__and2_1
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ _11053_/Y _11055_/B vssd1 vssd1 vccd1 vccd1 _13495_/A sky130_fd_sc_hd__nand2b_4
XFILLER_110_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15932_ _19729_/Q _15989_/A2 _15989_/B1 _19761_/Q vssd1 vssd1 vccd1 vccd1 _15932_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_283_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10006_ _10004_/X _10005_/X _11945_/S vssd1 vssd1 vccd1 vccd1 _10006_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18651_ _19516_/Q _18651_/B vssd1 vssd1 vccd1 vccd1 _18651_/Y sky130_fd_sc_hd__nand2_1
X_15863_ _16002_/A1 _15849_/Y _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15863_/X sky130_fd_sc_hd__a21o_1
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _20360_/Q _17913_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20360_/D sky130_fd_sc_hd__mux2_1
XFILLER_92_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14814_ _11416_/B _11735_/B _14815_/S vssd1 vssd1 vccd1 vccd1 _14814_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18582_ _18477_/X _18564_/A _18580_/Y _18581_/Y vssd1 vssd1 vccd1 vccd1 _18583_/B
+ sky130_fd_sc_hd__o211a_1
X_15794_ _15789_/X _15790_/Y _15793_/X vssd1 vssd1 vccd1 vccd1 _15794_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _17526_/C _20249_/Q _17522_/B vssd1 vssd1 vccd1 vccd1 _17533_/X sky130_fd_sc_hd__a21o_1
X_14745_ _19497_/Q _14773_/B vssd1 vssd1 vccd1 vccd1 _14745_/X sky130_fd_sc_hd__or2_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _11961_/B vssd1 vssd1 vccd1 vccd1 _13433_/A sky130_fd_sc_hd__clkinv_4
XFILLER_205_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10908_ _19802_/Q _09689_/D _10906_/X _09688_/A _10907_/X vssd1 vssd1 vccd1 vccd1
+ _10908_/X sky130_fd_sc_hd__o221a_1
X_17464_ _20267_/Q _17494_/B vssd1 vssd1 vccd1 vccd1 _17464_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14676_ _19435_/Q _17857_/A1 _14685_/S vssd1 vssd1 vccd1 vccd1 _19435_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11888_ _20390_/Q _20454_/Q _11891_/B vssd1 vssd1 vccd1 vccd1 _11888_/X sky130_fd_sc_hd__mux2_1
X_19203_ _20663_/CLK _19203_/D vssd1 vssd1 vccd1 vccd1 _19203_/Q sky130_fd_sc_hd__dfxtp_1
X_16415_ _19751_/Q _16418_/C _18821_/A vssd1 vssd1 vccd1 vccd1 _16415_/Y sky130_fd_sc_hd__a21oi_1
X_13627_ _13478_/B _13242_/C _15843_/A _13765_/A vssd1 vssd1 vccd1 vccd1 _13627_/X
+ sky130_fd_sc_hd__a22o_4
X_10839_ _19628_/Q _12323_/S _10824_/X _12324_/S vssd1 vssd1 vccd1 vccd1 _10839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17395_ _20246_/Q _17401_/A2 _17394_/X _17434_/A vssd1 vssd1 vccd1 vccd1 _20246_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19134_ _19511_/CLK _19134_/D vssd1 vssd1 vccd1 vccd1 _19134_/Q sky130_fd_sc_hd__dfxtp_1
X_16346_ _19724_/Q _19725_/Q _16346_/C vssd1 vssd1 vccd1 vccd1 _16348_/B sky130_fd_sc_hd__and3_1
XFILLER_201_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13558_ _13558_/A _13558_/B vssd1 vssd1 vccd1 vccd1 _13558_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_201_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19065_ _20410_/Q vssd1 vssd1 vccd1 vccd1 _20410_/D sky130_fd_sc_hd__clkbuf_2
X_12509_ _18765_/C _12585_/C _12509_/C vssd1 vssd1 vccd1 vccd1 _13107_/B sky130_fd_sc_hd__nor3_4
X_16277_ _19693_/Q _17708_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19693_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13489_ _09481_/Y _13564_/B _20948_/Q vssd1 vssd1 vccd1 vccd1 _13489_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15228_ _15218_/X _15226_/Y _15227_/X _15326_/A vssd1 vssd1 vccd1 vccd1 _15248_/A
+ sky130_fd_sc_hd__a31o_1
X_18016_ _20744_/Q _18019_/C _18104_/A vssd1 vssd1 vccd1 vccd1 _18016_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput404 _13797_/X vssd1 vssd1 vccd1 vccd1 din0[6] sky130_fd_sc_hd__buf_4
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput415 _19975_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[14] sky130_fd_sc_hd__buf_4
Xoutput426 _19985_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[24] sky130_fd_sc_hd__buf_4
XFILLER_154_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput437 _19966_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[5] sky130_fd_sc_hd__buf_4
Xoutput448 _20260_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[3] sky130_fd_sc_hd__buf_4
XFILLER_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15159_ _15165_/S _15062_/X _15158_/X vssd1 vssd1 vccd1 vccd1 _15159_/Y sky130_fd_sc_hd__o21ai_1
Xoutput459 _19512_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[18] sky130_fd_sc_hd__buf_4
XFILLER_102_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19967_ _20004_/CLK _19967_/D vssd1 vssd1 vccd1 vccd1 _19967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09720_ _19290_/Q _20077_/Q _11979_/S vssd1 vssd1 vccd1 vccd1 _09720_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18918_ _18973_/A _18918_/B vssd1 vssd1 vccd1 vccd1 _21002_/D sky130_fd_sc_hd__nor2_1
XFILLER_274_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19898_ _20341_/CLK _19898_/D vssd1 vssd1 vccd1 vccd1 _19898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09651_ _19590_/Q _09666_/B vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18849_ _18856_/A _18849_/B vssd1 vssd1 vccd1 vccd1 _20992_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09582_ _14112_/A _19085_/Q _19084_/Q vssd1 vssd1 vccd1 vccd1 _09588_/C sky130_fd_sc_hd__and3b_2
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20811_ _20812_/CLK _20811_/D vssd1 vssd1 vccd1 vccd1 _20811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_wb_clk_i ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_169_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20742_ _20742_/CLK _20742_/D vssd1 vssd1 vccd1 vccd1 _20742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20673_ _20673_/CLK _20673_/D vssd1 vssd1 vccd1 vccd1 _20673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1607 _12301_/S vssd1 vssd1 vccd1 vccd1 _12324_/S sky130_fd_sc_hd__buf_6
Xfanout1618 _10585_/S vssd1 vssd1 vccd1 vccd1 _09806_/S sky130_fd_sc_hd__buf_8
Xfanout620 _14205_/A2 vssd1 vssd1 vccd1 vccd1 _14398_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1629 fanout1630/X vssd1 vssd1 vccd1 vccd1 _11359_/S sky130_fd_sc_hd__buf_6
Xfanout631 _13889_/B1 vssd1 vssd1 vccd1 vccd1 _13881_/B1 sky130_fd_sc_hd__buf_4
Xfanout642 _16170_/S vssd1 vssd1 vccd1 vccd1 _16178_/S sky130_fd_sc_hd__buf_4
X_09918_ _09912_/X _09917_/X _12012_/S vssd1 vssd1 vccd1 vccd1 _09918_/X sky130_fd_sc_hd__mux2_1
X_20107_ _20482_/CLK _20107_/D vssd1 vssd1 vccd1 vccd1 _20107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout653 _16036_/A2 vssd1 vssd1 vccd1 vccd1 _16007_/A sky130_fd_sc_hd__buf_4
XFILLER_247_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout664 _14115_/Y vssd1 vssd1 vccd1 vccd1 _16068_/B sky130_fd_sc_hd__buf_6
Xfanout675 _13902_/B vssd1 vssd1 vccd1 vccd1 _17745_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_246_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout686 _14040_/A2 vssd1 vssd1 vccd1 vccd1 _19050_/S sky130_fd_sc_hd__clkbuf_8
X_20038_ _20673_/CLK _20038_/D vssd1 vssd1 vccd1 vccd1 _20038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09849_ _19887_/Q _19788_/Q _10397_/S vssd1 vssd1 vccd1 vccd1 _09849_/X sky130_fd_sc_hd__mux2_1
Xfanout697 _14073_/B vssd1 vssd1 vccd1 vccd1 _16133_/B sky130_fd_sc_hd__buf_6
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12860_ _12860_/A _12860_/B vssd1 vssd1 vccd1 vccd1 _13346_/C sky130_fd_sc_hd__xnor2_2
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _19422_/Q _11891_/B vssd1 vssd1 vccd1 vccd1 _11811_/X sky130_fd_sc_hd__or2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12791_/A _12791_/B _12791_/C _12791_/D vssd1 vssd1 vccd1 vccd1 _12791_/X
+ sky130_fd_sc_hd__or4_4
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _17918_/A _16672_/A vssd1 vssd1 vccd1 vccd1 _14531_/C sky130_fd_sc_hd__nor2_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11742_/A _11742_/B vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__and2_4
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _20226_/Q _19255_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14462_/B sky130_fd_sc_hd__mux2_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _20643_/Q _20607_/Q _11682_/S vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16200_ _19623_/Q _17886_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19623_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13412_ _13412_/A _13412_/B _13412_/C _13412_/D vssd1 vssd1 vccd1 vccd1 _13412_/X
+ sky130_fd_sc_hd__or4_4
X_17180_ _20146_/Q _17705_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20146_/D sky130_fd_sc_hd__mux2_1
X_10624_ _12850_/A1 _10620_/X _10623_/X _12085_/B2 vssd1 vssd1 vccd1 vccd1 _10624_/X
+ sky130_fd_sc_hd__o22a_1
X_14392_ _19521_/Q _14392_/B vssd1 vssd1 vccd1 vccd1 _14394_/A sky130_fd_sc_hd__xnor2_1
XFILLER_139_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16131_ _19590_/Q _16131_/A2 _16131_/B1 vssd1 vssd1 vccd1 vccd1 _16131_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13343_ _18593_/A2 _13342_/X _14306_/A1 vssd1 vssd1 vccd1 vccd1 _13343_/Y sky130_fd_sc_hd__o21ai_1
X_10555_ input124/X input159/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10555_/X sky130_fd_sc_hd__mux2_8
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16062_ _15948_/A1 _12914_/Y _16061_/X _16062_/B2 vssd1 vssd1 vccd1 vccd1 _16064_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_13274_ _13269_/X _13273_/X _13275_/A1 vssd1 vssd1 vccd1 vccd1 _13274_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_170_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ _11273_/A1 _19472_/Q _19440_/Q _10485_/S vssd1 vssd1 vccd1 vccd1 _10486_/X
+ sky130_fd_sc_hd__a22o_1
X_15013_ _15133_/B _15142_/S vssd1 vssd1 vccd1 vccd1 _15013_/Y sky130_fd_sc_hd__nor2_4
XFILLER_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12225_ _12215_/X _12217_/X _12224_/X _12383_/A _09502_/A vssd1 vssd1 vccd1 vccd1
+ _12225_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19821_ _20047_/CLK _19821_/D vssd1 vssd1 vccd1 vccd1 _19821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12156_ _12156_/A1 _12154_/X _12155_/X vssd1 vssd1 vccd1 vccd1 _12156_/X sky130_fd_sc_hd__a21o_1
XFILLER_78_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11107_ _19625_/Q _19931_/Q _19269_/Q _20056_/Q _12272_/B2 _12406_/C vssd1 vssd1
+ vccd1 vccd1 _11107_/X sky130_fd_sc_hd__mux4_1
X_19752_ _20621_/CLK _19752_/D vssd1 vssd1 vccd1 vccd1 _19752_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16964_ _19241_/Q _17003_/B _16964_/B1 _19110_/Q _16963_/X vssd1 vssd1 vccd1 vccd1
+ _16964_/X sky130_fd_sc_hd__o221a_1
X_12087_ _12085_/X _12086_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _12087_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18703_ _09479_/Y _18483_/B _18719_/S vssd1 vssd1 vccd1 vccd1 _18704_/B sky130_fd_sc_hd__mux2_1
XFILLER_204_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11038_ _12430_/S _11037_/Y _11034_/Y _11384_/S vssd1 vssd1 vccd1 vccd1 _11038_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_204_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15915_ _19760_/Q _15942_/A2 _15914_/X _15999_/C1 vssd1 vssd1 vccd1 vccd1 _15915_/X
+ sky130_fd_sc_hd__a211o_1
X_19683_ _20482_/CLK _19683_/D vssd1 vssd1 vccd1 vccd1 _19683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16895_ _16892_/Y _16894_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16895_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_77_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18634_ _18891_/A _18634_/B vssd1 vssd1 vccd1 vccd1 _20931_/D sky130_fd_sc_hd__nor2_1
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _11880_/B _12471_/X _15845_/Y _11878_/A vssd1 vssd1 vccd1 vccd1 _15846_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18565_ _18570_/B _18565_/B vssd1 vssd1 vccd1 vccd1 _18565_/Y sky130_fd_sc_hd__nor2_8
XFILLER_92_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ _16017_/C1 _15776_/X _15772_/X vssd1 vssd1 vccd1 vccd1 _15777_/X sky130_fd_sc_hd__o21a_2
XFILLER_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12989_ _19232_/Q _19231_/Q _19230_/Q _19229_/Q vssd1 vssd1 vccd1 vccd1 _12990_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_240_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17516_ _20293_/Q _17522_/B vssd1 vssd1 vccd1 vccd1 _17516_/Y sky130_fd_sc_hd__nand2_1
X_14728_ _19485_/Q _17666_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19485_/D sky130_fd_sc_hd__mux2_1
X_18496_ _18604_/B _18496_/B vssd1 vssd1 vccd1 vccd1 _18496_/X sky130_fd_sc_hd__or2_2
XANTENNA_580 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_591 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17447_ _17457_/A _17437_/X _17446_/Y _17445_/X _17443_/C vssd1 vssd1 vccd1 vccd1
+ _17447_/X sky130_fd_sc_hd__o32a_1
X_14659_ _19421_/Q _17666_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19421_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17378_ _20237_/Q _17378_/A2 _17382_/B1 _20286_/Q _17380_/C1 vssd1 vssd1 vccd1 vccd1
+ _17378_/X sky130_fd_sc_hd__a221o_4
XFILLER_220_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19117_ _19520_/CLK _19117_/D vssd1 vssd1 vccd1 vccd1 _19117_/Q sky130_fd_sc_hd__dfxtp_4
X_16329_ _19718_/Q _16330_/C _19719_/Q vssd1 vssd1 vccd1 vccd1 _16331_/B sky130_fd_sc_hd__a21oi_1
XFILLER_146_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19048_ _18315_/Y _19048_/A2 _19048_/B1 _12553_/C _19048_/C1 vssd1 vssd1 vccd1 vccd1
+ _19048_/X sky130_fd_sc_hd__a221o_1
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21010_ _21010_/CLK _21010_/D vssd1 vssd1 vccd1 vccd1 _21010_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput289 _13831_/X vssd1 vssd1 vccd1 vccd1 addr0[4] sky130_fd_sc_hd__buf_4
XFILLER_101_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09703_ _20141_/Q _20109_/Q _11889_/S vssd1 vssd1 vccd1 vccd1 _09703_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09634_ _14112_/A _19090_/Q _19088_/Q _19089_/Q vssd1 vssd1 vccd1 vccd1 _09634_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09565_ _09562_/X _14898_/A _09556_/X vssd1 vssd1 vccd1 vccd1 _12577_/A sky130_fd_sc_hd__a21oi_4
XFILLER_243_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09496_ _19231_/Q vssd1 vssd1 vccd1 vccd1 _09496_/Y sky130_fd_sc_hd__inv_2
XFILLER_270_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20725_ _20725_/CLK _20725_/D vssd1 vssd1 vccd1 vccd1 _20725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20656_ _20663_/CLK _20656_/D vssd1 vssd1 vccd1 vccd1 _20656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20587_ _20719_/CLK _20587_/D vssd1 vssd1 vccd1 vccd1 _20587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10340_ _10335_/X _10339_/X _12504_/A vssd1 vssd1 vccd1 vccd1 _10340_/X sky130_fd_sc_hd__a21o_1
XFILLER_165_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10271_ _10265_/X _10270_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _10271_/X sky130_fd_sc_hd__mux2_1
X_12010_ _20424_/Q _20360_/Q _20652_/Q _20616_/Q _12185_/S _12008_/C vssd1 vssd1 vccd1
+ vccd1 _12010_/X sky130_fd_sc_hd__mux4_1
XFILLER_215_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1404 _10345_/S vssd1 vssd1 vccd1 vccd1 _11295_/S sky130_fd_sc_hd__buf_6
XFILLER_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1415 fanout1422/X vssd1 vssd1 vccd1 vccd1 _12428_/S sky130_fd_sc_hd__buf_6
XFILLER_132_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1426 _12248_/B1 vssd1 vssd1 vccd1 vccd1 _12352_/S sky130_fd_sc_hd__buf_6
Xfanout1437 _09735_/Y vssd1 vssd1 vccd1 vccd1 _11852_/B2 sky130_fd_sc_hd__buf_8
XFILLER_238_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1448 _10405_/C vssd1 vssd1 vccd1 vccd1 _12084_/C sky130_fd_sc_hd__buf_6
Xfanout1459 _09734_/Y vssd1 vssd1 vccd1 vccd1 _11391_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_247_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13961_ _19186_/Q _14053_/C _14042_/S vssd1 vssd1 vccd1 vccd1 _13961_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout494 _17885_/X vssd1 vssd1 vccd1 vccd1 _17917_/S sky130_fd_sc_hd__buf_12
XFILLER_171_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12912_ _12912_/A _12912_/B vssd1 vssd1 vccd1 vccd1 _13106_/D sky130_fd_sc_hd__nand2_1
XFILLER_58_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15700_ _16051_/A1 _15686_/Y _16051_/B1 vssd1 vssd1 vccd1 vccd1 _15700_/Y sky130_fd_sc_hd__o21ai_1
X_16680_ _19935_/Q _17649_/A1 _16704_/S vssd1 vssd1 vccd1 vccd1 _19935_/D sky130_fd_sc_hd__mux2_1
XFILLER_247_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13892_ _19110_/Q _14040_/A2 _13896_/B1 _12513_/A _14458_/A vssd1 vssd1 vccd1 vccd1
+ _19110_/D sky130_fd_sc_hd__o221a_1
XFILLER_207_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15631_ _19718_/Q _15989_/A2 _15989_/B1 _19750_/Q vssd1 vssd1 vccd1 vccd1 _15631_/X
+ sky130_fd_sc_hd__a22o_1
X_12843_ _15659_/A _15527_/A vssd1 vssd1 vccd1 vccd1 _12843_/X sky130_fd_sc_hd__or2_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ _16002_/A1 _15561_/Y _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15562_/X sky130_fd_sc_hd__a21o_1
X_18350_ _20830_/Q _18349_/B _18349_/Y _18718_/A vssd1 vssd1 vccd1 vccd1 _20830_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_261_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _14803_/A1 _12582_/C _12784_/B _12773_/X vssd1 vssd1 vccd1 vccd1 _12774_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_203_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _20206_/Q _17328_/A2 _17299_/X _17300_/X _17974_/B1 vssd1 vssd1 vccd1 vccd1
+ _20206_/D sky130_fd_sc_hd__o221a_1
X_14513_ _19291_/Q _17876_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19291_/D sky130_fd_sc_hd__mux2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_48_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20586_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _15686_/A vssd1 vssd1 vccd1 vccd1 _11725_/Y sky130_fd_sc_hd__inv_2
XFILLER_261_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15493_ _19538_/Q _15492_/A _15492_/Y _16159_/C1 vssd1 vssd1 vccd1 vccd1 _19538_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18281_ _20810_/Q _18280_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18282_/B sky130_fd_sc_hd__mux2_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17232_ _17235_/A _17336_/B vssd1 vssd1 vccd1 vccd1 _17232_/X sky130_fd_sc_hd__and2_2
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14444_ _20298_/Q _17522_/B _17528_/B vssd1 vssd1 vccd1 vccd1 _14444_/X sky130_fd_sc_hd__or3_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11656_ _19416_/Q _11978_/S vssd1 vssd1 vccd1 vccd1 _11656_/X sky130_fd_sc_hd__or2_1
XFILLER_168_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17163_ _20129_/Q _17163_/A1 _17166_/S vssd1 vssd1 vccd1 vccd1 _20129_/D sky130_fd_sc_hd__mux2_1
X_10607_ _19807_/Q _10603_/B _10605_/X _12085_/B2 _10606_/X vssd1 vssd1 vccd1 vccd1
+ _10607_/X sky130_fd_sc_hd__o221a_1
X_14375_ _14366_/A _14363_/Y _14365_/B vssd1 vssd1 vccd1 vccd1 _14376_/B sky130_fd_sc_hd__o21a_1
X_11587_ _19681_/Q _20169_/Q _11979_/S vssd1 vssd1 vccd1 vccd1 _11587_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16114_ _09787_/X _16126_/A2 _16113_/X vssd1 vssd1 vccd1 vccd1 _19581_/D sky130_fd_sc_hd__o21a_1
XFILLER_155_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13326_ _13029_/Y _13326_/B vssd1 vssd1 vccd1 vccd1 _13327_/B sky130_fd_sc_hd__nand2b_1
XFILLER_182_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17094_ _20064_/Q _17896_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20064_/D sky130_fd_sc_hd__mux2_1
X_10538_ _12433_/A1 _10474_/X _10537_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _15443_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_127_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16045_ _20977_/Q _16045_/A2 _16016_/S _20849_/Q _16044_/X vssd1 vssd1 vccd1 vccd1
+ _16045_/X sky130_fd_sc_hd__a221o_1
X_13257_ _13334_/A _13253_/X _13254_/Y _13256_/Y vssd1 vssd1 vccd1 vccd1 _13257_/X
+ sky130_fd_sc_hd__o31a_2
X_10469_ _19585_/Q _10468_/X _11229_/S vssd1 vssd1 vccd1 vccd1 _10470_/B sky130_fd_sc_hd__mux2_4
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12208_ _19556_/Q _09613_/A _11225_/B _19620_/Q vssd1 vssd1 vccd1 vccd1 _12208_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_124_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13188_ _19299_/Q _13188_/B _15981_/A _14525_/B vssd1 vssd1 vccd1 vccd1 _13189_/B
+ sky130_fd_sc_hd__and4b_4
XFILLER_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19804_ _20061_/CLK _19804_/D vssd1 vssd1 vccd1 vccd1 _19804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_269_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12139_ _20653_/Q _20617_/Q _12139_/S vssd1 vssd1 vccd1 vccd1 _12139_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17996_ _20736_/Q _17997_/C _17995_/Y vssd1 vssd1 vccd1 vccd1 _20736_/D sky130_fd_sc_hd__o21a_1
XFILLER_215_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19735_ _21044_/CLK _19735_/D vssd1 vssd1 vccd1 vccd1 _19735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1960 _09515_/Y vssd1 vssd1 vccd1 vccd1 fanout1960/X sky130_fd_sc_hd__buf_4
X_16947_ _19239_/Q _16980_/A2 _16980_/B1 _19108_/Q _16946_/X vssd1 vssd1 vccd1 vccd1
+ _16947_/X sky130_fd_sc_hd__o221a_1
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1971 _18877_/A vssd1 vssd1 vccd1 vccd1 _18891_/A sky130_fd_sc_hd__buf_4
XFILLER_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1982 _18814_/A vssd1 vssd1 vccd1 vccd1 _18801_/A sky130_fd_sc_hd__clkbuf_4
Xfanout1993 _19051_/A vssd1 vssd1 vccd1 vccd1 _18056_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_226_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19666_ _20561_/CLK _19666_/D vssd1 vssd1 vccd1 vccd1 _19666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16878_ _16878_/A _16878_/B vssd1 vssd1 vccd1 vccd1 _16878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18617_ _18505_/X _18621_/A2 _18615_/Y _18616_/Y vssd1 vssd1 vccd1 vccd1 _18618_/B
+ sky130_fd_sc_hd__o211a_1
X_15829_ _20937_/Q _16044_/A2 _15828_/X vssd1 vssd1 vccd1 vccd1 _15829_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19597_ _19621_/CLK _19597_/D vssd1 vssd1 vccd1 vccd1 _19597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_252_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18548_ _20909_/Q _18559_/B _18547_/X _18458_/B vssd1 vssd1 vccd1 vccd1 _18549_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_240_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18479_ _18783_/A _18479_/B vssd1 vssd1 vccd1 vccd1 _20886_/D sky130_fd_sc_hd__nor2_1
XFILLER_221_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20510_ _20646_/CLK _20510_/D vssd1 vssd1 vccd1 vccd1 _20510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20441_ _20451_/CLK _20441_/D vssd1 vssd1 vccd1 vccd1 _20441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20372_ _20491_/CLK _20372_/D vssd1 vssd1 vccd1 vccd1 _20372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09617_ _12519_/C _09734_/B vssd1 vssd1 vccd1 vccd1 _09617_/Y sky130_fd_sc_hd__nor2_2
XFILLER_216_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09548_ _19152_/Q _19151_/Q _19150_/Q _13867_/A vssd1 vssd1 vccd1 vccd1 _12500_/D
+ sky130_fd_sc_hd__and4b_2
XFILLER_231_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09479_ _20952_/Q vssd1 vssd1 vccd1 vccd1 _09479_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11510_ _20134_/Q _20102_/Q _11916_/S vssd1 vssd1 vccd1 vccd1 _11510_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20708_ _20708_/CLK _20708_/D vssd1 vssd1 vccd1 vccd1 _20708_/Q sky130_fd_sc_hd__dfxtp_1
X_12490_ _13863_/A _12490_/B vssd1 vssd1 vccd1 vccd1 _12664_/C sky130_fd_sc_hd__nand2_8
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11441_ _19383_/Q _20674_/Q _12139_/S vssd1 vssd1 vccd1 vccd1 _11441_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20639_ _20671_/CLK _20639_/D vssd1 vssd1 vccd1 vccd1 _20639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _14160_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14161_/B sky130_fd_sc_hd__nor2_1
X_11372_ _20126_/Q _20094_/Q _11377_/S vssd1 vssd1 vccd1 vccd1 _11372_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13111_ _13103_/X _13110_/Y _09488_/A vssd1 vssd1 vccd1 vccd1 _13111_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10323_ _11273_/A1 _19911_/Q _11256_/S _10311_/X vssd1 vssd1 vccd1 vccd1 _10323_/X
+ sky130_fd_sc_hd__o211a_1
X_14091_ _14105_/A _14107_/B _14091_/C vssd1 vssd1 vccd1 vccd1 _14091_/X sky130_fd_sc_hd__or3_1
XFILLER_180_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_166_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21043_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13042_ _20957_/Q _20891_/Q vssd1 vssd1 vccd1 vccd1 _13453_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10254_ _10252_/X _10253_/X _11378_/S vssd1 vssd1 vccd1 vccd1 _10254_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1201 _17324_/C1 vssd1 vssd1 vccd1 vccd1 _17330_/C1 sky130_fd_sc_hd__buf_4
XFILLER_133_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17850_ _17850_/A _17850_/B vssd1 vssd1 vccd1 vccd1 _17851_/C sky130_fd_sc_hd__nor2_1
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1212 _15025_/X vssd1 vssd1 vccd1 vccd1 _16002_/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10185_ _19636_/Q _19942_/Q _19280_/Q _20067_/Q _12346_/S _11391_/C vssd1 vssd1 vccd1
+ vccd1 _10185_/X sky130_fd_sc_hd__mux4_1
Xfanout1223 _13519_/S vssd1 vssd1 vccd1 vccd1 _13607_/B sky130_fd_sc_hd__buf_6
Xfanout1234 _09684_/X vssd1 vssd1 vccd1 vccd1 _12039_/A1 sky130_fd_sc_hd__buf_6
X_16801_ _16726_/X _16800_/Y _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16801_/X sky130_fd_sc_hd__a21o_2
Xfanout1245 _17337_/Y vssd1 vssd1 vccd1 vccd1 _17370_/B1 sky130_fd_sc_hd__buf_6
Xfanout1256 _12930_/X vssd1 vssd1 vccd1 vccd1 _16716_/A sky130_fd_sc_hd__buf_8
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17781_ _20558_/Q _17921_/A1 _17794_/S vssd1 vssd1 vccd1 vccd1 _20558_/D sky130_fd_sc_hd__mux2_1
Xfanout1267 _09607_/X vssd1 vssd1 vccd1 vccd1 _12155_/B1 sky130_fd_sc_hd__buf_6
X_14993_ _20882_/Q _14992_/X _14993_/S vssd1 vssd1 vccd1 vccd1 _14993_/X sky130_fd_sc_hd__mux2_1
Xfanout1278 _16034_/S vssd1 vssd1 vccd1 vccd1 _11649_/S sky130_fd_sc_hd__buf_8
XFILLER_120_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19520_ _19520_/CLK _19520_/D vssd1 vssd1 vccd1 vccd1 _19520_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1289 _09546_/Y vssd1 vssd1 vccd1 vccd1 _12581_/A sky130_fd_sc_hd__buf_6
X_16732_ _16869_/A _16732_/B vssd1 vssd1 vccd1 vccd1 _16732_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13944_ _16187_/A _13944_/B vssd1 vssd1 vccd1 vccd1 _19146_/D sky130_fd_sc_hd__and2_1
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19451_ _20710_/CLK _19451_/D vssd1 vssd1 vccd1 vccd1 _19451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13875_ _19093_/Q _13953_/A2 _13881_/B1 _19159_/Q _16197_/A vssd1 vssd1 vccd1 vccd1
+ _19093_/D sky130_fd_sc_hd__o221a_1
XFILLER_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16663_ _19920_/Q _17107_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19920_/D sky130_fd_sc_hd__mux2_1
X_18402_ _18708_/A _18402_/B vssd1 vssd1 vccd1 vccd1 _20855_/D sky130_fd_sc_hd__and2_1
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12826_ _12823_/Y _12825_/X _15703_/B2 vssd1 vssd1 vccd1 vccd1 _12829_/B sky130_fd_sc_hd__a21oi_4
XFILLER_90_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15614_ _10277_/A _11416_/B _16057_/A2 _15613_/X vssd1 vssd1 vccd1 vccd1 _15614_/X
+ sky130_fd_sc_hd__o22a_1
X_19382_ _20673_/CLK _19382_/D vssd1 vssd1 vccd1 vccd1 _19382_/Q sky130_fd_sc_hd__dfxtp_1
X_16594_ _16598_/A _16594_/B _16594_/C vssd1 vssd1 vccd1 vccd1 _16595_/A sky130_fd_sc_hd__and3_1
XFILLER_131_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18333_ _18477_/B _18341_/B vssd1 vssd1 vccd1 vccd1 _18333_/Y sky130_fd_sc_hd__nand2_1
XFILLER_199_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15545_ _15545_/A _15545_/B vssd1 vssd1 vccd1 vccd1 _15545_/Y sky130_fd_sc_hd__nand2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12755_/X _12756_/Y _12752_/B vssd1 vssd1 vccd1 vccd1 _12757_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_199_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _20575_/Q _11708_/B vssd1 vssd1 vccd1 vccd1 _11708_/X sky130_fd_sc_hd__or2_1
X_15476_ _20733_/Q _16041_/A2 _16041_/B1 _20765_/Q vssd1 vssd1 vccd1 vccd1 _15476_/X
+ sky130_fd_sc_hd__a22o_1
X_18264_ _18299_/A1 _14332_/B _18263_/Y vssd1 vssd1 vccd1 vccd1 _18529_/B sky130_fd_sc_hd__o21ai_4
X_12688_ _13511_/A _13511_/B vssd1 vssd1 vccd1 vccd1 _13526_/B sky130_fd_sc_hd__and2_1
XFILLER_129_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17215_ _20179_/Q _17949_/A1 _17215_/S vssd1 vssd1 vccd1 vccd1 _20179_/D sky130_fd_sc_hd__mux2_1
X_14427_ _14427_/A _14427_/B _14432_/B vssd1 vssd1 vccd1 vccd1 _14427_/Y sky130_fd_sc_hd__nor3_1
X_11639_ _12003_/A _20041_/Q _19916_/Q _11932_/S0 vssd1 vssd1 vccd1 vccd1 _11639_/X
+ sky130_fd_sc_hd__a22o_1
X_18195_ _18487_/B vssd1 vssd1 vccd1 vccd1 _18195_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14358_ _13205_/A _14357_/X _13262_/Y vssd1 vssd1 vccd1 vccd1 _14359_/C sky130_fd_sc_hd__o21a_1
X_17146_ _20114_/Q _17705_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20114_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13309_ _13309_/A _13309_/B vssd1 vssd1 vccd1 vccd1 _13309_/X sky130_fd_sc_hd__or2_1
X_17077_ _20049_/Q _17111_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20049_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14289_ _19511_/Q _14294_/B vssd1 vssd1 vccd1 vccd1 _14303_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16028_ _16028_/A _16028_/B _16028_/C vssd1 vssd1 vccd1 vccd1 _16028_/X sky130_fd_sc_hd__and3_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17979_ _20731_/Q _17982_/C vssd1 vssd1 vccd1 vccd1 _17985_/C sky130_fd_sc_hd__and2_1
XFILLER_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19718_ _19978_/CLK _19718_/D vssd1 vssd1 vccd1 vccd1 _19718_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_242_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1790 _18198_/B vssd1 vssd1 vccd1 vccd1 _18163_/A sky130_fd_sc_hd__buf_6
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20990_ _20990_/CLK _20990_/D vssd1 vssd1 vccd1 vccd1 _20990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19649_ _20647_/CLK _19649_/D vssd1 vssd1 vccd1 vccd1 _19649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20424_ _20706_/CLK _20424_/D vssd1 vssd1 vccd1 vccd1 _20424_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20355_ _20683_/CLK _20355_/D vssd1 vssd1 vccd1 vccd1 _20355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20286_ _21011_/CLK _20286_/D vssd1 vssd1 vccd1 vccd1 _20286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ _19650_/Q _11994_/S _11966_/X _11995_/S vssd1 vssd1 vccd1 vccd1 _11990_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10941_ _11021_/A _20497_/Q _11035_/S _20529_/Q vssd1 vssd1 vccd1 vccd1 _10941_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_272_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ _13775_/A _13660_/B vssd1 vssd1 vccd1 vccd1 _13660_/X sky130_fd_sc_hd__and2_1
XFILLER_271_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10872_ _19667_/Q _12344_/S _11212_/S vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__o21a_1
XFILLER_189_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _19518_/Q _12872_/B vssd1 vssd1 vccd1 vccd1 _12884_/B sky130_fd_sc_hd__and2_2
XFILLER_213_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13591_/A _13591_/B vssd1 vssd1 vccd1 vccd1 _13591_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15330_ _19533_/Q _15402_/A _15329_/Y _16197_/A vssd1 vssd1 vccd1 vccd1 _19533_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _20878_/Q _12549_/B _12542_/C vssd1 vssd1 vccd1 vccd1 _12550_/B sky130_fd_sc_hd__and3_1
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ _14841_/S _15105_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _15261_/X sky130_fd_sc_hd__o21a_1
X_12473_ _14895_/A _14897_/A vssd1 vssd1 vccd1 vccd1 _14853_/S sky130_fd_sc_hd__nor2_4
X_17000_ _16950_/Y _16999_/X _16875_/B2 vssd1 vssd1 vccd1 vccd1 _17000_/Y sky130_fd_sc_hd__o21bai_4
X_14212_ _14208_/B _14211_/Y _14233_/S vssd1 vssd1 vccd1 vccd1 _14212_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11424_ _11514_/A1 _12138_/A1 _19351_/Q _12129_/S vssd1 vssd1 vccd1 vccd1 _11424_/X
+ sky130_fd_sc_hd__a31o_1
X_15192_ _21015_/Q _20983_/Q _15309_/S vssd1 vssd1 vccd1 vccd1 _15192_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_8 _15419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14143_ _12584_/A _14142_/X _13491_/X vssd1 vssd1 vccd1 vccd1 _14144_/C sky130_fd_sc_hd__a21o_1
X_11355_ _19374_/Q _20665_/Q _11358_/S vssd1 vssd1 vccd1 vccd1 _11355_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _11259_/S _10304_/X _10305_/X vssd1 vssd1 vccd1 vccd1 _10306_/X sky130_fd_sc_hd__o21a_1
X_14074_ _19196_/Q _14106_/A2 _14073_/X _17963_/B1 vssd1 vssd1 vccd1 vccd1 _19196_/D
+ sky130_fd_sc_hd__o211a_1
X_18951_ _21007_/Q _18978_/B vssd1 vssd1 vccd1 vccd1 _18951_/Y sky130_fd_sc_hd__nand2_1
X_11286_ _19798_/Q _11291_/A2 _11284_/X _11291_/B2 _11285_/X vssd1 vssd1 vccd1 vccd1
+ _11286_/X sky130_fd_sc_hd__o221a_1
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17902_ _20673_/Q _17902_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20673_/D sky130_fd_sc_hd__mux2_1
X_13025_ _20966_/Q _20900_/Q vssd1 vssd1 vccd1 vccd1 _13025_/Y sky130_fd_sc_hd__nor2_2
X_10237_ _19282_/Q _20069_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _10237_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18882_ _20997_/Q _18978_/B vssd1 vssd1 vccd1 vccd1 _18882_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1020 _12583_/Y vssd1 vssd1 vccd1 vccd1 _18785_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_266_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1031 _17006_/A1 vssd1 vssd1 vccd1 vccd1 _16981_/A1 sky130_fd_sc_hd__buf_4
Xfanout1042 _11152_/X vssd1 vssd1 vccd1 vccd1 _17887_/A1 sky130_fd_sc_hd__buf_6
X_17833_ _20608_/Q _17871_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20608_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10168_ _12429_/A1 _10166_/X _10167_/X vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__o21a_1
Xfanout1053 _10894_/X vssd1 vssd1 vccd1 vccd1 _17890_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1064 _10728_/X vssd1 vssd1 vccd1 vccd1 _17926_/A1 sky130_fd_sc_hd__buf_6
XFILLER_255_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1075 _17885_/B vssd1 vssd1 vccd1 vccd1 _17574_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_120_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1086 _17916_/A1 vssd1 vssd1 vccd1 vccd1 _17950_/A1 sky130_fd_sc_hd__buf_4
XFILLER_281_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1097 _12156_/X vssd1 vssd1 vccd1 vccd1 _17914_/A1 sky130_fd_sc_hd__buf_4
X_17764_ _20543_/Q _17870_/A1 _17772_/S vssd1 vssd1 vccd1 vccd1 _20543_/D sky130_fd_sc_hd__mux2_1
X_14976_ _15314_/B _14979_/B vssd1 vssd1 vccd1 vccd1 _14978_/B sky130_fd_sc_hd__nor2_2
X_10099_ _20409_/Q _20345_/Q _20637_/Q _20601_/Q _10092_/S _10405_/C vssd1 vssd1 vccd1
+ vccd1 _10099_/X sky130_fd_sc_hd__mux4_1
XFILLER_212_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19503_ _19506_/CLK _19503_/D vssd1 vssd1 vccd1 vccd1 _19503_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_63_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20664_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16715_ _16715_/A vssd1 vssd1 vccd1 vccd1 _17219_/C sky130_fd_sc_hd__inv_2
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13927_ _19131_/Q _13906_/B _13932_/B1 _13388_/D vssd1 vssd1 vccd1 vccd1 _19131_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_223_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17695_ _20479_/Q _17695_/A1 _17703_/S vssd1 vssd1 vccd1 vccd1 _20479_/D sky130_fd_sc_hd__mux2_1
XFILLER_212_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19434_ _20561_/CLK _19434_/D vssd1 vssd1 vccd1 vccd1 _19434_/Q sky130_fd_sc_hd__dfxtp_1
X_16646_ _19903_/Q _17649_/A1 _16670_/S vssd1 vssd1 vccd1 vccd1 _19903_/D sky130_fd_sc_hd__mux2_1
XFILLER_228_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13858_ _16598_/A _16594_/B _19661_/Q _09648_/Y vssd1 vssd1 vccd1 vccd1 _13860_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_50_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19365_ _20720_/CLK _19365_/D vssd1 vssd1 vccd1 vccd1 _19365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12809_ _13253_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _13389_/A sky130_fd_sc_hd__and2_2
XFILLER_250_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16577_ _16591_/A _16577_/B vssd1 vssd1 vccd1 vccd1 _19854_/D sky130_fd_sc_hd__or2_1
XFILLER_210_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13789_ _16240_/A1 _13610_/X _13612_/X _13438_/Y vssd1 vssd1 vccd1 vccd1 _13789_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18316_ _20817_/Q _18315_/Y _18316_/S vssd1 vssd1 vccd1 vccd1 _18317_/B sky130_fd_sc_hd__mux2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ _15528_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _15528_/Y sky130_fd_sc_hd__nand2_1
X_19296_ _20662_/CLK _19296_/D vssd1 vssd1 vccd1 vccd1 _19296_/Q sky130_fd_sc_hd__dfxtp_1
X_18247_ _18720_/A _18247_/B vssd1 vssd1 vccd1 vccd1 _20803_/D sky130_fd_sc_hd__and2_1
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15459_ _14808_/Y _15456_/X _15457_/Y _15458_/Y _15442_/Y vssd1 vssd1 vccd1 vccd1
+ _15459_/X sky130_fd_sc_hd__o311a_1
XFILLER_163_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18178_ _19531_/Q _18198_/B vssd1 vssd1 vccd1 vccd1 _18178_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_144_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17129_ _20097_/Q _17163_/A1 _17132_/S vssd1 vssd1 vccd1 vccd1 _20097_/D sky130_fd_sc_hd__mux2_1
XFILLER_274_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09951_ _19418_/Q _11891_/B vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__or2_1
X_20140_ _20579_/CLK _20140_/D vssd1 vssd1 vccd1 vccd1 _20140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20071_ _20446_/CLK _20071_/D vssd1 vssd1 vccd1 vccd1 _20071_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _19683_/Q _20171_/Q _11527_/S vssd1 vssd1 vccd1 vccd1 _09882_/X sky130_fd_sc_hd__mux2_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20973_ _21041_/CLK _20973_/D vssd1 vssd1 vccd1 vccd1 _20973_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_409 _17676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_272_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20407_ _20635_/CLK _20407_/D vssd1 vssd1 vccd1 vccd1 _20407_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_135_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11140_ _11140_/A _11140_/B vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__or2_4
X_20338_ _20630_/CLK _20338_/D vssd1 vssd1 vccd1 vccd1 _20338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11071_ _12306_/A1 _20691_/Q _11074_/S _11070_/X vssd1 vssd1 vccd1 vccd1 _11071_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20269_ _21016_/CLK _20269_/D vssd1 vssd1 vccd1 vccd1 _20269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput101 dout0[62] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_hd__clkbuf_2
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput112 dout1[14] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_hd__clkbuf_2
X_10022_ _09612_/X _09636_/B _10020_/Y vssd1 vssd1 vccd1 vccd1 _11234_/B sky130_fd_sc_hd__a21o_4
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput123 dout1[24] vssd1 vssd1 vccd1 vccd1 input123/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput134 dout1[34] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__clkbuf_2
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 dout1[44] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__buf_2
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput156 dout1[54] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__clkbuf_2
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput167 dout1[6] vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_hd__clkbuf_2
X_14830_ _10803_/B _12115_/B _14882_/B vssd1 vssd1 vccd1 vccd1 _14830_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput178 irq[1] vssd1 vssd1 vccd1 vccd1 _12540_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 jtag_tms vssd1 vssd1 vccd1 vccd1 _17452_/A sky130_fd_sc_hd__buf_6
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11973_ _11969_/X _11972_/X _12129_/S vssd1 vssd1 vccd1 vccd1 _11973_/X sky130_fd_sc_hd__mux2_1
X_14761_ _19505_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14761_/X sky130_fd_sc_hd__or2_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16500_ _19807_/Q _17686_/A1 _16517_/S vssd1 vssd1 vccd1 vccd1 _19807_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10924_ _19869_/Q _19770_/Q _10924_/S vssd1 vssd1 vccd1 vccd1 _10924_/X sky130_fd_sc_hd__mux2_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _13712_/A _13730_/B vssd1 vssd1 vccd1 vccd1 _13752_/B sky130_fd_sc_hd__or2_1
X_17480_ _20275_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17480_/Y sky130_fd_sc_hd__nand2_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _19451_/Q _17941_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19451_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _19757_/Q _16434_/C _18863_/A vssd1 vssd1 vccd1 vccd1 _16431_/Y sky130_fd_sc_hd__a21oi_1
X_10855_ _19628_/Q _19934_/Q _19272_/Q _20059_/Q _12334_/S0 _12337_/C vssd1 vssd1
+ vccd1 vccd1 _10855_/X sky130_fd_sc_hd__mux4_1
X_13643_ _13663_/A _13663_/B _13666_/B vssd1 vssd1 vccd1 vccd1 _13643_/X sky130_fd_sc_hd__and3_4
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19150_ _19620_/CLK _19150_/D vssd1 vssd1 vccd1 vccd1 _19150_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13574_ _19222_/Q _19221_/Q _13545_/B _19223_/Q vssd1 vssd1 vccd1 vccd1 _13575_/B
+ sky130_fd_sc_hd__a31o_1
X_16362_ _19730_/Q _19731_/Q _16362_/C vssd1 vssd1 vccd1 vccd1 _16364_/B sky130_fd_sc_hd__and3_4
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _20156_/Q _11379_/B vssd1 vssd1 vccd1 vccd1 _10786_/X sky130_fd_sc_hd__or2_1
XFILLER_201_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18101_ _20775_/Q _20774_/Q _18101_/C vssd1 vssd1 vccd1 vccd1 _18103_/B sky130_fd_sc_hd__and3_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15313_ _20856_/Q _14971_/B _15311_/X _15312_/Y _14971_/C vssd1 vssd1 vccd1 vccd1
+ _15313_/X sky130_fd_sc_hd__a221o_1
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ _13350_/A _13107_/B vssd1 vssd1 vccd1 vccd1 _12525_/Y sky130_fd_sc_hd__nor2_8
X_19081_ _20426_/Q vssd1 vssd1 vccd1 vccd1 _20426_/D sky130_fd_sc_hd__clkbuf_2
X_16293_ _16293_/A _16293_/B vssd1 vssd1 vccd1 vccd1 _19705_/D sky130_fd_sc_hd__nor2_1
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_181_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20300_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18032_ _20749_/Q _18028_/B _18031_/Y vssd1 vssd1 vccd1 vccd1 _20749_/D sky130_fd_sc_hd__o21a_1
XFILLER_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ _16050_/A1 _15243_/X _15229_/X vssd1 vssd1 vccd1 vccd1 _15246_/B sky130_fd_sc_hd__a21oi_1
X_12456_ _12464_/A _12468_/B _12464_/C vssd1 vssd1 vccd1 vccd1 _16054_/B sky130_fd_sc_hd__o21a_4
Xclkbuf_leaf_110_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19992_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11407_ _10645_/A _11772_/B _11406_/X vssd1 vssd1 vccd1 vccd1 _11407_/X sky130_fd_sc_hd__a21bo_1
X_15175_ _15611_/S _15175_/B vssd1 vssd1 vccd1 vccd1 _15175_/Y sky130_fd_sc_hd__nor2_1
X_12387_ _20655_/Q _20619_/Q _12389_/S vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14126_ _14204_/A _16068_/B _14126_/C vssd1 vssd1 vccd1 vccd1 _14126_/X sky130_fd_sc_hd__or3_1
X_11338_ _11338_/A1 _11335_/X _11337_/X vssd1 vssd1 vccd1 vccd1 _11338_/X sky130_fd_sc_hd__a21o_1
XFILLER_181_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19983_ _20862_/CLK _19983_/D vssd1 vssd1 vccd1 vccd1 _19983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14057_ _14107_/A _14069_/B _14057_/C vssd1 vssd1 vccd1 vccd1 _14057_/X sky130_fd_sc_hd__or3_1
X_18934_ _18955_/A _18934_/B vssd1 vssd1 vccd1 vccd1 _18934_/Y sky130_fd_sc_hd__nand2_1
X_11269_ _19267_/Q _09688_/B _09688_/A vssd1 vssd1 vccd1 vccd1 _11269_/X sky130_fd_sc_hd__a21o_1
XFILLER_239_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13008_ _20975_/Q _20909_/Q vssd1 vssd1 vccd1 vccd1 _13134_/B sky130_fd_sc_hd__nand2_1
XFILLER_228_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18865_ _18968_/A _18865_/B vssd1 vssd1 vccd1 vccd1 _18865_/Y sky130_fd_sc_hd__nand2_1
XFILLER_255_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17816_ _20591_/Q _17888_/A1 _17844_/S vssd1 vssd1 vccd1 vccd1 _20591_/D sky130_fd_sc_hd__mux2_1
XFILLER_283_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18796_ _19089_/Q _18785_/A2 _12591_/X _13539_/B vssd1 vssd1 vccd1 vccd1 _18796_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17747_ _20526_/Q _17887_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20526_/D sky130_fd_sc_hd__mux2_1
XFILLER_282_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14959_ _15314_/B _14959_/B vssd1 vssd1 vccd1 vccd1 _14997_/C sky130_fd_sc_hd__nor2_1
XFILLER_282_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17678_ _20462_/Q _17678_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20462_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19417_ _20716_/CLK _19417_/D vssd1 vssd1 vccd1 vccd1 _19417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16629_ _19888_/Q _17666_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19888_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19348_ _20703_/CLK _19348_/D vssd1 vssd1 vccd1 vccd1 _19348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19279_ _20472_/CLK _19279_/D vssd1 vssd1 vccd1 vccd1 _19279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20123_ _20155_/CLK _20123_/D vssd1 vssd1 vccd1 vccd1 _20123_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout802 _17505_/A1 vssd1 vssd1 vccd1 vccd1 _17525_/A1 sky130_fd_sc_hd__buf_4
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ _12020_/C1 _09933_/X _11872_/A vssd1 vssd1 vccd1 vccd1 _09934_/Y sky130_fd_sc_hd__a21oi_2
Xfanout813 _13798_/A1 vssd1 vssd1 vccd1 vccd1 _13776_/B1 sky130_fd_sc_hd__buf_8
Xfanout824 _15013_/Y vssd1 vssd1 vccd1 vccd1 _15482_/A2 sky130_fd_sc_hd__buf_4
XFILLER_259_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout835 _18690_/Y vssd1 vssd1 vccd1 vccd1 _18749_/S sky130_fd_sc_hd__buf_6
Xfanout846 _18324_/Y vssd1 vssd1 vccd1 vccd1 _18357_/B sky130_fd_sc_hd__buf_4
Xfanout857 _15015_/X vssd1 vssd1 vccd1 vccd1 _15998_/A2 sky130_fd_sc_hd__buf_8
X_20054_ _20315_/CLK _20054_/D vssd1 vssd1 vccd1 vccd1 _20054_/Q sky130_fd_sc_hd__dfxtp_1
X_09865_ _19548_/Q _12155_/A2 _12155_/B1 _19612_/Q vssd1 vssd1 vccd1 vccd1 _09865_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout868 _15309_/S vssd1 vssd1 vccd1 vccd1 _15508_/S sky130_fd_sc_hd__clkbuf_16
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout879 _16039_/B vssd1 vssd1 vccd1 vccd1 _15933_/B sky130_fd_sc_hd__clkbuf_4
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _19420_/Q _10426_/S _09795_/X _12051_/C1 vssd1 vssd1 vccd1 vccd1 _09796_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_285_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_206 _20216_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_228 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_239 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20956_ _21022_/CLK _20956_/D vssd1 vssd1 vccd1 vccd1 _20956_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _21019_/CLK _20887_/D vssd1 vssd1 vccd1 vccd1 _20887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _10455_/B _10640_/B vssd1 vssd1 vccd1 vccd1 _10640_/X sky130_fd_sc_hd__and2b_1
XFILLER_201_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10571_ _19775_/Q _12043_/B vssd1 vssd1 vccd1 vccd1 _10571_/X sky130_fd_sc_hd__or2_1
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12310_ _12304_/X _12306_/X _12309_/X _11345_/S _12310_/C1 vssd1 vssd1 vccd1 vccd1
+ _12310_/X sky130_fd_sc_hd__o221a_1
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ _13290_/A _13290_/B _13290_/C vssd1 vssd1 vccd1 vccd1 _13290_/X sky130_fd_sc_hd__and3_1
XFILLER_213_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12241_ _12239_/X _12240_/X _12241_/S vssd1 vssd1 vccd1 vccd1 _12241_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12172_ _11849_/S _12169_/X _12171_/X _12183_/C1 vssd1 vssd1 vccd1 vccd1 _12172_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_268_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ _12347_/A1 _19336_/Q _20691_/Q _11126_/B _12347_/C1 vssd1 vssd1 vccd1 vccd1
+ _11123_/X sky130_fd_sc_hd__a221o_1
X_16980_ _19243_/Q _16980_/A2 _16980_/B1 _19112_/Q _16979_/X vssd1 vssd1 vccd1 vccd1
+ _16980_/X sky130_fd_sc_hd__o221a_1
XFILLER_3_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ _15545_/A _11054_/B vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__nand2_2
X_15931_ _15931_/A _16037_/B vssd1 vssd1 vccd1 vccd1 _15931_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10005_ _20138_/Q _20106_/Q _11944_/S vssd1 vssd1 vccd1 vccd1 _10005_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18650_ _20936_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18650_/Y sky130_fd_sc_hd__nand2_1
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _15973_/A1 _15861_/X _15849_/Y vssd1 vssd1 vccd1 vccd1 _15862_/X sky130_fd_sc_hd__a21bo_1
XFILLER_77_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17601_ _20359_/Q _17878_/A1 _17601_/S vssd1 vssd1 vccd1 vccd1 _20359_/D sky130_fd_sc_hd__mux2_1
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14813_ _14811_/X _14812_/X _15058_/S vssd1 vssd1 vccd1 vccd1 _14813_/X sky130_fd_sc_hd__mux2_1
XFILLER_218_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _19498_/Q _18760_/B vssd1 vssd1 vccd1 vccd1 _18581_/Y sky130_fd_sc_hd__nand2_2
XFILLER_264_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _13414_/A _12565_/B _15791_/X _15792_/X vssd1 vssd1 vccd1 vccd1 _15793_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_280_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17532_ _17532_/A _17532_/B vssd1 vssd1 vccd1 vccd1 _20298_/D sky130_fd_sc_hd__nor2_1
XFILLER_205_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _19119_/Q _14764_/A2 _14743_/X _14758_/C1 vssd1 vssd1 vccd1 vccd1 _19496_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_217_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _11956_/A _15887_/S vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__nor2_4
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10907_ _11008_/A1 _19306_/Q _09623_/B _10152_/S vssd1 vssd1 vccd1 vccd1 _10907_/X
+ sky130_fd_sc_hd__o31a_1
X_17463_ _17487_/A1 _17462_/Y _18598_/A vssd1 vssd1 vccd1 vccd1 _20266_/D sky130_fd_sc_hd__a21oi_1
X_14675_ _19434_/Q _17924_/A1 _14685_/S vssd1 vssd1 vccd1 vccd1 _19434_/D sky130_fd_sc_hd__mux2_1
X_11887_ _20486_/Q _20326_/Q _11891_/B vssd1 vssd1 vccd1 vccd1 _11887_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19202_ _20426_/CLK _19202_/D vssd1 vssd1 vccd1 vccd1 _19202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16414_ _19750_/Q _16412_/B _16413_/Y vssd1 vssd1 vccd1 vccd1 _19750_/D sky130_fd_sc_hd__o21a_1
X_10838_ _12309_/S _10837_/X _10836_/X _12399_/A1 vssd1 vssd1 vccd1 vccd1 _10838_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13626_ _13626_/A1 _13412_/A _15816_/A _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13626_/X
+ sky130_fd_sc_hd__a22o_4
X_17394_ _20245_/Q _17337_/B _17530_/A2 _20294_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17394_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ _19511_/CLK _19133_/D vssd1 vssd1 vccd1 vccd1 _19133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16345_ _19724_/Q _16346_/C _19725_/Q vssd1 vssd1 vccd1 vccd1 _16347_/B sky130_fd_sc_hd__a21oi_1
X_10769_ _19804_/Q _12412_/A2 _10767_/X _12412_/B2 _10768_/X vssd1 vssd1 vccd1 vccd1
+ _10769_/X sky130_fd_sc_hd__o221a_1
X_13557_ _13544_/A _13544_/B _12698_/C vssd1 vssd1 vccd1 vccd1 _13558_/B sky130_fd_sc_hd__a21oi_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _13897_/A _12508_/B _12517_/B _09695_/Y vssd1 vssd1 vccd1 vccd1 _12509_/C
+ sky130_fd_sc_hd__or4b_2
X_19064_ _20409_/Q vssd1 vssd1 vccd1 vccd1 _20409_/D sky130_fd_sc_hd__clkbuf_2
X_16276_ _19692_/Q _17950_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19692_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13488_ _12652_/B _13484_/Y _13487_/Y vssd1 vssd1 vccd1 vccd1 _13488_/X sky130_fd_sc_hd__a21o_1
XFILLER_173_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18015_ _20743_/Q _18013_/B _18014_/Y vssd1 vssd1 vccd1 vccd1 _20743_/D sky130_fd_sc_hd__o21a_1
X_15227_ _13523_/A _12471_/X _14837_/S _15224_/Y _15222_/X vssd1 vssd1 vccd1 vccd1
+ _15227_/X sky130_fd_sc_hd__o221a_1
X_12439_ _12202_/A _12202_/B _13183_/A _13182_/A _13178_/A vssd1 vssd1 vccd1 vccd1
+ _12450_/A sky130_fd_sc_hd__a2111o_4
Xoutput405 _13798_/X vssd1 vssd1 vccd1 vccd1 din0[7] sky130_fd_sc_hd__buf_4
Xoutput416 _19976_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[15] sky130_fd_sc_hd__buf_4
XFILLER_218_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput427 _19986_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[25] sky130_fd_sc_hd__buf_4
Xoutput438 _19967_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[6] sky130_fd_sc_hd__buf_4
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15158_ _15167_/S _15158_/B vssd1 vssd1 vccd1 vccd1 _15158_/X sky130_fd_sc_hd__or2_1
Xoutput449 _20261_/Q vssd1 vssd1 vccd1 vccd1 probe_jtagInstruction[4] sky130_fd_sc_hd__buf_4
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _14003_/S _14081_/A _14522_/A vssd1 vssd1 vccd1 vccd1 _19214_/D sky130_fd_sc_hd__a21oi_1
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15089_ _17275_/A _15482_/A2 _15088_/X vssd1 vssd1 vccd1 vccd1 _15089_/X sky130_fd_sc_hd__a21o_1
X_19966_ _19978_/CLK _19966_/D vssd1 vssd1 vccd1 vccd1 _19966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18917_ _18532_/X _18971_/B _18915_/X _18916_/Y vssd1 vssd1 vccd1 vccd1 _18918_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_256_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19897_ _20315_/CLK _19897_/D vssd1 vssd1 vccd1 vccd1 _19897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09650_ _11228_/A1 _14041_/A2 _09647_/X _09649_/X vssd1 vssd1 vccd1 vccd1 _09650_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_41_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18848_ _18502_/X _18861_/B _18846_/X _18847_/Y vssd1 vssd1 vccd1 vccd1 _18849_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_267_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09581_ _09578_/X _12972_/B _09580_/X _09604_/A _19089_/Q vssd1 vssd1 vccd1 vccd1
+ _09585_/C sky130_fd_sc_hd__o32ai_4
XFILLER_243_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18779_ _19119_/Q _18830_/A _18778_/X vssd1 vssd1 vccd1 vccd1 _18779_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_209_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20810_ _21043_/CLK _20810_/D vssd1 vssd1 vccd1 vccd1 _20810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20741_ _20742_/CLK _20741_/D vssd1 vssd1 vccd1 vccd1 _20741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20672_ _20672_/CLK _20672_/D vssd1 vssd1 vccd1 vccd1 _20672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1608 _12301_/S vssd1 vssd1 vccd1 vccd1 _12241_/S sky130_fd_sc_hd__clkbuf_4
Xfanout610 _14567_/X vssd1 vssd1 vccd1 vccd1 _14599_/S sky130_fd_sc_hd__buf_12
XFILLER_266_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout621 _14205_/A2 vssd1 vssd1 vccd1 vccd1 _14256_/A2 sky130_fd_sc_hd__buf_6
Xfanout1619 fanout1630/X vssd1 vssd1 vccd1 vccd1 _10585_/S sky130_fd_sc_hd__buf_6
X_20106_ _20481_/CLK _20106_/D vssd1 vssd1 vccd1 vccd1 _20106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout632 _13863_/Y vssd1 vssd1 vccd1 vccd1 _13889_/B1 sky130_fd_sc_hd__buf_6
X_09917_ _09915_/X _09916_/X _11849_/S vssd1 vssd1 vccd1 vccd1 _09917_/X sky130_fd_sc_hd__mux2_1
Xfanout643 _16170_/S vssd1 vssd1 vccd1 vccd1 _16196_/S sky130_fd_sc_hd__buf_4
Xfanout654 _14810_/X vssd1 vssd1 vccd1 vccd1 _16036_/A2 sky130_fd_sc_hd__buf_4
Xfanout665 _14115_/Y vssd1 vssd1 vccd1 vccd1 _14204_/B sky130_fd_sc_hd__buf_2
Xfanout676 _13902_/B vssd1 vssd1 vccd1 vccd1 _17851_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_247_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20037_ _20692_/CLK _20037_/D vssd1 vssd1 vccd1 vccd1 _20037_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout687 _14040_/A2 vssd1 vssd1 vccd1 vccd1 _14043_/A2 sky130_fd_sc_hd__buf_4
XFILLER_37_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09848_ _09829_/A _19484_/Q _19452_/Q _10397_/S _12100_/B1 vssd1 vssd1 vccd1 vccd1
+ _09848_/X sky130_fd_sc_hd__a221o_1
Xfanout698 _14107_/A vssd1 vssd1 vccd1 vccd1 _14099_/A sky130_fd_sc_hd__buf_4
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _17909_/A1 _12194_/A1 _12194_/B2 _09778_/X vssd1 vssd1 vccd1 vccd1 _15822_/A
+ sky130_fd_sc_hd__a22o_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11810_ _19953_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__or2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _13586_/A _12790_/B _12790_/C _12790_/D vssd1 vssd1 vccd1 vccd1 _12791_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11741_/A vssd1 vssd1 vccd1 vccd1 _11743_/A sky130_fd_sc_hd__clkinv_2
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20939_ _21009_/CLK _20939_/D vssd1 vssd1 vccd1 vccd1 _20939_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _18692_/A _14460_/B vssd1 vssd1 vccd1 vccd1 _19254_/D sky130_fd_sc_hd__and2_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _12051_/A1 _20511_/Q _12056_/S _11654_/X vssd1 vssd1 vccd1 vccd1 _11672_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10623_ _10621_/X _10622_/X _12023_/S vssd1 vssd1 vccd1 vccd1 _10623_/X sky130_fd_sc_hd__mux2_1
X_13411_ _13411_/A _13411_/B vssd1 vssd1 vccd1 vccd1 _13412_/D sky130_fd_sc_hd__or2_1
X_14391_ _20293_/Q _14431_/A2 _14431_/B1 input234/X vssd1 vssd1 vccd1 vccd1 _14392_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_139_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16130_ _10288_/X _16132_/A2 _16129_/X vssd1 vssd1 vccd1 vccd1 _19589_/D sky130_fd_sc_hd__o21a_1
X_13342_ _20963_/Q _13355_/B _13340_/Y _13341_/X vssd1 vssd1 vccd1 vccd1 _13342_/X
+ sky130_fd_sc_hd__a22o_1
X_10554_ _10032_/Y _11150_/B _09638_/Y vssd1 vssd1 vccd1 vccd1 _10554_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13273_ _13272_/B _13270_/X _13271_/Y _13272_/Y _18560_/A vssd1 vssd1 vccd1 vccd1
+ _13273_/X sky130_fd_sc_hd__o311a_1
X_16061_ _15544_/A _16052_/X _16060_/X _15527_/B vssd1 vssd1 vccd1 vccd1 _16061_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_182_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10485_ _19875_/Q _19776_/Q _10485_/S vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15012_ _15314_/B _15012_/B _15021_/C vssd1 vssd1 vccd1 vccd1 _15142_/S sky130_fd_sc_hd__or3b_4
X_12224_ _12222_/X _12223_/X _12376_/S vssd1 vssd1 vccd1 vccd1 _12224_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19820_ _20479_/CLK _19820_/D vssd1 vssd1 vccd1 vccd1 _19820_/Q sky130_fd_sc_hd__dfxtp_1
X_12155_ _19555_/Q _12155_/A2 _12155_/B1 _19619_/Q vssd1 vssd1 vccd1 vccd1 _12155_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11106_ _19800_/Q _12412_/A2 _11104_/X _12412_/B2 _11105_/X vssd1 vssd1 vccd1 vccd1
+ _11106_/X sky130_fd_sc_hd__o221a_1
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19751_ _21017_/CLK _19751_/D vssd1 vssd1 vccd1 vccd1 _19751_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16963_ _20423_/Q _16963_/A2 _16963_/B1 vssd1 vssd1 vccd1 vccd1 _16963_/X sky130_fd_sc_hd__a21o_1
X_12086_ _20423_/Q _20359_/Q _20651_/Q _20615_/Q _10628_/S _12084_/C vssd1 vssd1 vccd1
+ vccd1 _12086_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18702_ _18702_/A _18702_/B vssd1 vssd1 vccd1 vccd1 _20951_/D sky130_fd_sc_hd__and2_1
XFILLER_277_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11037_ _12429_/A1 _11035_/X _11036_/X vssd1 vssd1 vccd1 vccd1 _11037_/Y sky130_fd_sc_hd__o21ai_1
X_15914_ _20812_/Q _15941_/A2 _15907_/X _15941_/B2 _15913_/X vssd1 vssd1 vccd1 vccd1
+ _15914_/X sky130_fd_sc_hd__a221o_4
XFILLER_231_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19682_ _20481_/CLK _19682_/D vssd1 vssd1 vccd1 vccd1 _19682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16894_ _16885_/A _16893_/X _16866_/B2 vssd1 vssd1 vccd1 vccd1 _16894_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18633_ _18517_/X _18688_/A2 _18631_/Y _18632_/Y vssd1 vssd1 vccd1 vccd1 _18634_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_280_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _11878_/B _15984_/A2 _15984_/B1 vssd1 vssd1 vccd1 vccd1 _15845_/Y sky130_fd_sc_hd__a21oi_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18564_ _18564_/A vssd1 vssd1 vccd1 vccd1 _18565_/B sky130_fd_sc_hd__inv_2
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _20967_/Q _16045_/A2 _16016_/S _20839_/Q _15775_/X vssd1 vssd1 vccd1 vccd1
+ _15776_/X sky130_fd_sc_hd__a221o_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _19228_/Q _19227_/Q _19226_/Q vssd1 vssd1 vccd1 vccd1 _12990_/B sky130_fd_sc_hd__and3_1
XFILLER_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17515_ _17525_/A1 _17514_/Y _17430_/A vssd1 vssd1 vccd1 vccd1 _20292_/D sky130_fd_sc_hd__a21oi_1
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14727_ _19484_/Q _17802_/A1 _14733_/S vssd1 vssd1 vccd1 vccd1 _19484_/D sky130_fd_sc_hd__mux2_1
X_18495_ _18598_/A _18495_/B vssd1 vssd1 vccd1 vccd1 _20891_/D sky130_fd_sc_hd__nor2_1
X_11939_ _20486_/Q _11616_/B _11948_/A1 vssd1 vssd1 vccd1 vccd1 _11939_/X sky130_fd_sc_hd__a21o_1
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_570 _19089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_581 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_592 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17446_ _17446_/A _17446_/B vssd1 vssd1 vccd1 vccd1 _17446_/Y sky130_fd_sc_hd__nor2_1
XFILLER_221_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14658_ _19420_/Q _17802_/A1 _14662_/S vssd1 vssd1 vccd1 vccd1 _19420_/D sky130_fd_sc_hd__mux2_1
XFILLER_221_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13609_ _13609_/A _13609_/B vssd1 vssd1 vccd1 vccd1 _13609_/Y sky130_fd_sc_hd__nand2_1
X_17377_ _20237_/Q _17381_/A2 _17376_/X _14482_/A vssd1 vssd1 vccd1 vccd1 _20237_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14589_ _19355_/Q _17941_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19355_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19116_ _21044_/CLK _19116_/D vssd1 vssd1 vccd1 vccd1 _19116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16328_ _19718_/Q _16330_/C _16327_/Y vssd1 vssd1 vccd1 vccd1 _19718_/D sky130_fd_sc_hd__o21a_1
XFILLER_174_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19047_ _21042_/Q _19049_/A2 _19046_/X _18740_/A vssd1 vssd1 vccd1 vccd1 _21042_/D
+ sky130_fd_sc_hd__o211a_1
X_16259_ _19675_/Q _17199_/A1 _16275_/S vssd1 vssd1 vccd1 vccd1 _19675_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19949_ _20717_/CLK _19949_/D vssd1 vssd1 vccd1 vccd1 _19949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09702_ _19685_/Q _20173_/Q _11889_/S vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__mux2_1
XFILLER_261_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09633_ _19550_/Q _12155_/A2 _12155_/B1 _19614_/Q vssd1 vssd1 vccd1 vccd1 _09633_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09564_ _12464_/A _14112_/B _12468_/B vssd1 vssd1 vccd1 vccd1 _14897_/A sky130_fd_sc_hd__or3b_4
XFILLER_270_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_213_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20710_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_271_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _09666_/B vssd1 vssd1 vccd1 vccd1 _09495_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20724_ _20794_/CLK _20724_/D vssd1 vssd1 vccd1 vccd1 _20724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20655_ _20655_/CLK _20655_/D vssd1 vssd1 vccd1 vccd1 _20655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20586_ _20586_/CLK _20586_/D vssd1 vssd1 vccd1 vccd1 _20586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ _10268_/X _10269_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _10270_/X sky130_fd_sc_hd__mux2_1
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1405 _10345_/S vssd1 vssd1 vccd1 vccd1 _10518_/S sky130_fd_sc_hd__buf_6
Xfanout1416 fanout1422/X vssd1 vssd1 vccd1 vccd1 _12417_/S sky130_fd_sc_hd__buf_4
XFILLER_48_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1427 _12248_/B1 vssd1 vssd1 vccd1 vccd1 _12334_/S0 sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1438 _15129_/A0 vssd1 vssd1 vccd1 vccd1 _11291_/B2 sky130_fd_sc_hd__buf_6
Xfanout1449 _10611_/B vssd1 vssd1 vccd1 vccd1 _10405_/C sky130_fd_sc_hd__buf_6
XFILLER_87_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13960_ _14041_/A1 _13960_/A2 _10890_/X _14041_/B1 _19835_/Q vssd1 vssd1 vccd1 vccd1
+ _14053_/C sky130_fd_sc_hd__o32a_1
XFILLER_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout495 _17885_/X vssd1 vssd1 vccd1 vccd1 _17916_/S sky130_fd_sc_hd__buf_6
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12911_ _12911_/A _12911_/B vssd1 vssd1 vccd1 vccd1 _12912_/B sky130_fd_sc_hd__or2_1
XFILLER_101_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13891_ _19109_/Q _19050_/S _13896_/B1 _12513_/B _14458_/A vssd1 vssd1 vccd1 vccd1
+ _19109_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ _15630_/A _16037_/B vssd1 vssd1 vccd1 vccd1 _15630_/X sky130_fd_sc_hd__or2_1
X_12842_ _12866_/A _12864_/B _13300_/B _12842_/D vssd1 vssd1 vccd1 vccd1 _13248_/A
+ sky130_fd_sc_hd__nand4b_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15561_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15561_/Y sky130_fd_sc_hd__nand2_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12781_/B _12773_/B vssd1 vssd1 vccd1 vccd1 _12773_/X sky130_fd_sc_hd__or2_1
XFILLER_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17300_ _20205_/Q _17327_/A2 _17330_/C1 vssd1 vssd1 vccd1 vccd1 _17300_/X sky130_fd_sc_hd__a21o_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _19290_/Q _17107_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19290_/D sky130_fd_sc_hd__mux2_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _18538_/B vssd1 vssd1 vccd1 vccd1 _18280_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _12107_/A1 _17904_/A1 _11723_/Y _09750_/Y vssd1 vssd1 vccd1 vccd1 _15686_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_15492_ _15492_/A _15492_/B vssd1 vssd1 vccd1 vccd1 _15492_/Y sky130_fd_sc_hd__nand2_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17231_/A _17235_/B vssd1 vssd1 vccd1 vccd1 _17336_/B sky130_fd_sc_hd__or2_4
X_14443_ _20244_/Q _14443_/B _17337_/A vssd1 vssd1 vccd1 vccd1 _17528_/B sky130_fd_sc_hd__or3_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11655_ _19947_/Q _12044_/B vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__or2_1
XFILLER_156_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_88_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19704_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17162_ _20128_/Q _17930_/A1 _17166_/S vssd1 vssd1 vccd1 vccd1 _20128_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _09834_/A _19311_/Q _10405_/C _12023_/S vssd1 vssd1 vccd1 vccd1 _10606_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_127_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14374_ _14372_/Y _14374_/B vssd1 vssd1 vccd1 vccd1 _14376_/A sky130_fd_sc_hd__and2b_1
X_11586_ _19948_/Q _11895_/B vssd1 vssd1 vccd1 vccd1 _11586_/X sky130_fd_sc_hd__or2_1
XFILLER_196_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16113_ _19581_/Q _16131_/A2 _16129_/B1 vssd1 vssd1 vccd1 vccd1 _16113_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10537_ _10525_/X _10536_/X _11396_/S vssd1 vssd1 vccd1 vccd1 _10537_/X sky130_fd_sc_hd__mux2_2
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13325_ _13350_/A _13300_/C _13321_/Y _13324_/X vssd1 vssd1 vccd1 vccd1 _13325_/X
+ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_17_wb_clk_i _20408_/CLK vssd1 vssd1 vccd1 vccd1 _20647_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17093_ _20063_/Q _17929_/A1 _17111_/S vssd1 vssd1 vccd1 vccd1 _20063_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16044_ _20945_/Q _16044_/A2 _16043_/X vssd1 vssd1 vccd1 vccd1 _16044_/X sky130_fd_sc_hd__o21a_1
XFILLER_109_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10468_ _11242_/A1 _14038_/A2 _10467_/X _11242_/B1 _19857_/Q vssd1 vssd1 vccd1 vccd1
+ _10468_/X sky130_fd_sc_hd__o32a_1
X_13256_ _20937_/Q _13363_/B _13323_/C _13255_/Y _18667_/B vssd1 vssd1 vccd1 vccd1
+ _13256_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_269_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _12288_/C _12207_/B vssd1 vssd1 vccd1 vccd1 _12207_/Y sky130_fd_sc_hd__nand2_2
X_13187_ _13188_/B _13631_/B vssd1 vssd1 vccd1 vccd1 _13437_/A sky130_fd_sc_hd__nor2_1
X_10399_ _19673_/Q _20161_/Q _10400_/S vssd1 vssd1 vccd1 vccd1 _10399_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19803_ _20662_/CLK _19803_/D vssd1 vssd1 vccd1 vccd1 _19803_/Q sky130_fd_sc_hd__dfxtp_1
X_12138_ _12138_/A1 _20521_/Q _12143_/S _12130_/X vssd1 vssd1 vccd1 vccd1 _12138_/X
+ sky130_fd_sc_hd__o211a_1
X_17995_ _17998_/A _17995_/B vssd1 vssd1 vccd1 vccd1 _17995_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1950 _17331_/C1 vssd1 vssd1 vccd1 vccd1 _17274_/C1 sky130_fd_sc_hd__buf_4
X_19734_ _21020_/CLK _19734_/D vssd1 vssd1 vccd1 vccd1 _19734_/Q sky130_fd_sc_hd__dfxtp_2
X_16946_ _20421_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16946_/X sky130_fd_sc_hd__a21o_1
X_12069_ _20048_/Q _19923_/Q _12070_/S vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__mux2_1
Xfanout1961 _17532_/A vssd1 vssd1 vccd1 vccd1 _17430_/A sky130_fd_sc_hd__buf_6
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1972 _18877_/A vssd1 vssd1 vccd1 vccd1 _18104_/A sky130_fd_sc_hd__buf_4
XFILLER_93_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1983 _17952_/A vssd1 vssd1 vccd1 vccd1 _18814_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_265_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1994 fanout2002/X vssd1 vssd1 vccd1 vccd1 _19051_/A sky130_fd_sc_hd__clkbuf_4
X_19665_ _20692_/CLK _19665_/D vssd1 vssd1 vccd1 vccd1 _19665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16877_ _19976_/Q _16876_/A _16876_/Y _18126_/A vssd1 vssd1 vccd1 vccd1 _19976_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18616_ _19507_/Q _18616_/B vssd1 vssd1 vccd1 vccd1 _18616_/Y sky130_fd_sc_hd__nand2_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _20905_/Q _16043_/A2 _16043_/B1 _15827_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _15828_/X sky130_fd_sc_hd__a221o_1
X_19596_ _19621_/CLK _19596_/D vssd1 vssd1 vccd1 vccd1 _19596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18547_ _18560_/A _18547_/B vssd1 vssd1 vccd1 vccd1 _18547_/X sky130_fd_sc_hd__or2_1
XFILLER_280_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15759_ _11281_/A _15978_/A2 _13417_/A _15949_/A vssd1 vssd1 vccd1 vccd1 _15760_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_206_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18478_ _20886_/Q fanout753/X _18477_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18479_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17429_ _20259_/Q _20252_/Q _17433_/S vssd1 vssd1 vccd1 vccd1 _17430_/B sky130_fd_sc_hd__mux2_1
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20440_ _20568_/CLK _20440_/D vssd1 vssd1 vccd1 vccd1 _20440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20371_ _20467_/CLK _20371_/D vssd1 vssd1 vccd1 vccd1 _20371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09616_ _17538_/C _09689_/A vssd1 vssd1 vccd1 vccd1 _09616_/Y sky130_fd_sc_hd__nor2_1
XFILLER_56_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09547_ _12580_/A _09556_/A vssd1 vssd1 vccd1 vccd1 _09547_/X sky130_fd_sc_hd__or2_4
XFILLER_271_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09478_ _20981_/Q vssd1 vssd1 vccd1 vccd1 _09478_/Y sky130_fd_sc_hd__inv_2
XPHY_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20707_ _20715_/CLK _20707_/D vssd1 vssd1 vccd1 vccd1 _20707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11440_ _20414_/Q _12148_/S _11426_/X _09901_/S vssd1 vssd1 vccd1 vccd1 _11440_/X
+ sky130_fd_sc_hd__o211a_1
X_20638_ _20638_/CLK _20638_/D vssd1 vssd1 vccd1 vccd1 _20638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11371_ _12357_/A1 _11369_/X _11370_/X vssd1 vssd1 vccd1 vccd1 _11371_/X sky130_fd_sc_hd__o21a_1
XFILLER_109_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20569_ _20701_/CLK _20569_/D vssd1 vssd1 vccd1 vccd1 _20569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10322_ _10320_/X _10321_/X _10322_/S vssd1 vssd1 vccd1 vccd1 _10322_/X sky130_fd_sc_hd__mux2_1
X_13110_ _13105_/X _13108_/X _13109_/X vssd1 vssd1 vccd1 vccd1 _13110_/Y sky130_fd_sc_hd__a21oi_1
X_14090_ _19204_/Q _14106_/A2 _14089_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1 _19204_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13041_ _20957_/Q _20891_/Q vssd1 vssd1 vccd1 vccd1 _13453_/A sky130_fd_sc_hd__or2_2
X_10253_ _19880_/Q _19781_/Q _11042_/B vssd1 vssd1 vccd1 vccd1 _10253_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1202 _17233_/Y vssd1 vssd1 vccd1 vccd1 _17324_/C1 sky130_fd_sc_hd__clkbuf_4
X_10184_ _19811_/Q _11392_/A2 _10182_/X _09738_/A _10183_/X vssd1 vssd1 vccd1 vccd1
+ _10184_/X sky130_fd_sc_hd__o221a_1
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1213 _16052_/A1 vssd1 vssd1 vccd1 vccd1 _16024_/A1 sky130_fd_sc_hd__buf_4
Xfanout1224 _13519_/S vssd1 vssd1 vccd1 vccd1 _13564_/B sky130_fd_sc_hd__buf_4
XFILLER_79_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1235 _09684_/X vssd1 vssd1 vccd1 vccd1 _12366_/A1 sky130_fd_sc_hd__buf_2
X_16800_ _16800_/A vssd1 vssd1 vccd1 vccd1 _16800_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_94_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1246 _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17400_/C1 sky130_fd_sc_hd__buf_4
XFILLER_121_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17780_ _20557_/Q _17780_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20557_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14992_ _20980_/Q _14956_/Y _15508_/S _21012_/Q _14991_/X vssd1 vssd1 vccd1 vccd1
+ _14992_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_135_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _19219_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout1257 _16063_/A2 vssd1 vssd1 vccd1 vccd1 _15978_/A2 sky130_fd_sc_hd__buf_4
XFILLER_93_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1268 _18152_/C vssd1 vssd1 vccd1 vccd1 _11225_/B sky130_fd_sc_hd__buf_4
Xfanout1279 _16034_/S vssd1 vssd1 vccd1 vccd1 _11726_/S sky130_fd_sc_hd__buf_6
XFILLER_247_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16731_ _19961_/Q _16822_/A _16730_/Y _18801_/A vssd1 vssd1 vccd1 vccd1 _19961_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_120_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13943_ _19146_/Q _13141_/X _13943_/S vssd1 vssd1 vccd1 vccd1 _13944_/B sky130_fd_sc_hd__mux2_1
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19450_ _20712_/CLK _19450_/D vssd1 vssd1 vccd1 vccd1 _19450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16662_ _19919_/Q _17874_/A1 _16666_/S vssd1 vssd1 vccd1 vccd1 _19919_/D sky130_fd_sc_hd__mux2_1
X_13874_ _19092_/Q _13953_/A2 _13881_/B1 _19158_/Q _16197_/A vssd1 vssd1 vccd1 vccd1
+ _19092_/D sky130_fd_sc_hd__o221a_1
XFILLER_46_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18401_ _20855_/Q _18185_/Y _18419_/S vssd1 vssd1 vccd1 vccd1 _18402_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15613_ _16058_/A2 _15264_/B _15613_/S vssd1 vssd1 vccd1 vccd1 _15613_/X sky130_fd_sc_hd__mux2_1
X_19381_ _20672_/CLK _19381_/D vssd1 vssd1 vccd1 vccd1 _19381_/Q sky130_fd_sc_hd__dfxtp_1
X_12825_ split8/X _12847_/A2 _15526_/A _12824_/X vssd1 vssd1 vccd1 vccd1 _12825_/X
+ sky130_fd_sc_hd__a211o_1
X_16593_ _16593_/A _16593_/B vssd1 vssd1 vccd1 vccd1 _19862_/D sky130_fd_sc_hd__or2_1
XFILLER_216_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18332_ _20821_/Q _18341_/B _18331_/Y _18698_/A vssd1 vssd1 vccd1 vccd1 _20821_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15544_ _15544_/A _15544_/B vssd1 vssd1 vccd1 vccd1 _15544_/X sky130_fd_sc_hd__or2_1
XFILLER_203_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _15473_/A _12784_/B vssd1 vssd1 vccd1 vccd1 _12756_/Y sky130_fd_sc_hd__nand2_1
XFILLER_188_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18263_ _19548_/Q _18308_/B vssd1 vssd1 vccd1 vccd1 _18263_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _09839_/A _11696_/X _11700_/X _11706_/X vssd1 vssd1 vccd1 vccd1 _11723_/A
+ sky130_fd_sc_hd__a31o_1
X_15475_ _19713_/Q _15475_/A2 _15475_/B1 _19745_/Q vssd1 vssd1 vccd1 vccd1 _15475_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12687_ _13526_/A _12692_/C vssd1 vssd1 vccd1 vccd1 _13511_/B sky130_fd_sc_hd__nor2_1
XFILLER_202_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17214_ _20178_/Q _17705_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20178_/D sky130_fd_sc_hd__mux2_1
X_14426_ _14426_/A _14432_/A _14426_/C _14426_/D vssd1 vssd1 vccd1 vccd1 _14432_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_175_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18194_ _18213_/B _14188_/B _18193_/Y vssd1 vssd1 vccd1 vccd1 _18487_/B sky130_fd_sc_hd__o21ai_4
X_11638_ _11641_/S _11635_/X _11637_/X vssd1 vssd1 vccd1 vccd1 _11638_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17145_ _20113_/Q _17704_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20113_/D sky130_fd_sc_hd__mux2_1
X_14357_ _14352_/B _14356_/Y _14417_/S vssd1 vssd1 vccd1 vccd1 _14357_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11569_ _12194_/A1 _11534_/X _11568_/Y _09750_/Y vssd1 vssd1 vccd1 vccd1 _15630_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_156_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13308_ _13373_/A _19234_/Q _14776_/C1 _13307_/Y vssd1 vssd1 vccd1 vccd1 _13361_/A
+ sky130_fd_sc_hd__o211a_1
X_17076_ _20048_/Q _17178_/A1 _17076_/S vssd1 vssd1 vccd1 vccd1 _20048_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14288_ _20283_/Q _14330_/A2 _14330_/B1 input223/X vssd1 vssd1 vccd1 vccd1 _14294_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_143_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16027_ _12436_/A _12443_/B _16057_/A2 _16026_/X vssd1 vssd1 vccd1 vccd1 _16027_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13239_ _13373_/A _13239_/B _13239_/C vssd1 vssd1 vccd1 vccd1 _13239_/X sky130_fd_sc_hd__and3_1
XFILLER_171_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17978_ _20730_/Q _17975_/A _17977_/Y vssd1 vssd1 vccd1 vccd1 _20730_/D sky130_fd_sc_hd__o21a_1
XFILLER_78_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19717_ _20862_/CLK _19717_/D vssd1 vssd1 vccd1 vccd1 _19717_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1780 _20262_/Q vssd1 vssd1 vccd1 vccd1 _17423_/D sky130_fd_sc_hd__buf_2
X_16929_ _20419_/Q _16963_/A2 _16963_/B1 vssd1 vssd1 vccd1 vccd1 _16929_/X sky130_fd_sc_hd__a21o_1
XFILLER_284_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1791 _18199_/A1 vssd1 vssd1 vccd1 vccd1 _18198_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_266_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19648_ _20682_/CLK _19648_/D vssd1 vssd1 vccd1 vccd1 _19648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19579_ _19590_/CLK _19579_/D vssd1 vssd1 vccd1 vccd1 _19579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20423_ _20666_/CLK _20423_/D vssd1 vssd1 vccd1 vccd1 _20423_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_181_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20354_ _20646_/CLK _20354_/D vssd1 vssd1 vccd1 vccd1 _20354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20285_ _21043_/CLK _20285_/D vssd1 vssd1 vccd1 vccd1 _20285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10940_ _10938_/X _10939_/X _11033_/S vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10871_ _20155_/Q _11379_/B vssd1 vssd1 vccd1 vccd1 _10871_/X sky130_fd_sc_hd__or2_1
XFILLER_231_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _19517_/Q _19516_/Q _12804_/B vssd1 vssd1 vccd1 vccd1 _12872_/B sky130_fd_sc_hd__and3_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13590_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13591_/B sky130_fd_sc_hd__nor2_1
XFILLER_243_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12541_ _20879_/Q _12549_/B _12541_/C vssd1 vssd1 vccd1 vccd1 _12553_/B sky130_fd_sc_hd__and3_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _13539_/B _15127_/B _15220_/X _15259_/Y vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12472_ _12463_/A _15264_/B _12469_/X _12463_/Y vssd1 vssd1 vccd1 vccd1 _12472_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_185_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14211_ _14211_/A _14211_/B vssd1 vssd1 vccd1 vccd1 _14211_/Y sky130_fd_sc_hd__xnor2_1
X_11423_ _19415_/Q _12124_/S _11422_/X _11423_/C1 vssd1 vssd1 vccd1 vccd1 _11423_/X
+ sky130_fd_sc_hd__o211a_1
X_15191_ input283/X _14930_/X _15142_/S vssd1 vssd1 vccd1 vccd1 _15191_/X sky130_fd_sc_hd__a21o_1
XFILLER_137_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_9 _15419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _20405_/Q _11358_/S _11349_/X _12301_/S vssd1 vssd1 vccd1 vccd1 _11354_/X
+ sky130_fd_sc_hd__o211a_1
X_14142_ _14139_/B _14141_/Y _14202_/S vssd1 vssd1 vccd1 vccd1 _14142_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10305_ _11273_/A1 _19348_/Q _20703_/Q _10485_/S _12519_/C vssd1 vssd1 vccd1 vccd1
+ _10305_/X sky130_fd_sc_hd__a221o_1
XFILLER_141_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14073_ _14099_/A _14073_/B _14073_/C vssd1 vssd1 vccd1 vccd1 _14073_/X sky130_fd_sc_hd__or3_1
X_11285_ _11290_/A _19302_/Q _11290_/C vssd1 vssd1 vccd1 vccd1 _11285_/X sky130_fd_sc_hd__or3_1
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18950_ _18671_/Y _18977_/A2 _18948_/Y _18949_/Y vssd1 vssd1 vccd1 vccd1 _18950_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17901_ _20672_/Q _17901_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20672_/D sky130_fd_sc_hd__mux2_1
X_10236_ _11258_/A1 _19912_/Q _10235_/S _10224_/X vssd1 vssd1 vccd1 vccd1 _10236_/X
+ sky130_fd_sc_hd__o211a_1
X_13024_ _20967_/Q _20901_/Q vssd1 vssd1 vccd1 vccd1 _13270_/B sky130_fd_sc_hd__nand2_1
X_18881_ _18632_/Y _18970_/A2 _18879_/Y _18880_/Y vssd1 vssd1 vccd1 vccd1 _18881_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1010 _15259_/B vssd1 vssd1 vccd1 vccd1 _15127_/B sky130_fd_sc_hd__clkbuf_8
Xfanout1021 _16963_/B1 vssd1 vssd1 vccd1 vccd1 _16979_/B1 sky130_fd_sc_hd__buf_4
X_17832_ _20607_/Q _17870_/A1 _17840_/S vssd1 vssd1 vccd1 vccd1 _20607_/D sky130_fd_sc_hd__mux2_1
XFILLER_126_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10167_ _10262_/A _19347_/Q _20702_/Q _11042_/B _11378_/S vssd1 vssd1 vccd1 vccd1
+ _10167_/X sky130_fd_sc_hd__a221o_1
Xfanout1032 _14902_/X vssd1 vssd1 vccd1 vccd1 _17006_/A1 sky130_fd_sc_hd__buf_4
Xfanout1043 _16608_/A1 vssd1 vssd1 vccd1 vccd1 _17922_/A1 sky130_fd_sc_hd__buf_4
Xfanout1054 _10894_/X vssd1 vssd1 vccd1 vccd1 _17750_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_67_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1065 _11397_/B2 vssd1 vssd1 vccd1 vccd1 _12194_/B2 sky130_fd_sc_hd__buf_6
XFILLER_254_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17763_ _20542_/Q _17869_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20542_/D sky130_fd_sc_hd__mux2_1
Xfanout1076 _18949_/B1 vssd1 vssd1 vccd1 vccd1 _18767_/B sky130_fd_sc_hd__buf_6
X_14975_ _14987_/A _14979_/B vssd1 vssd1 vccd1 vccd1 _14975_/Y sky130_fd_sc_hd__nor2_1
Xfanout1087 _12367_/X vssd1 vssd1 vccd1 vccd1 _17916_/A1 sky130_fd_sc_hd__buf_8
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10098_ _19378_/Q _10603_/B _10096_/X _12085_/B2 _10097_/X vssd1 vssd1 vccd1 vccd1
+ _10098_/X sky130_fd_sc_hd__o221a_1
XFILLER_187_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1098 _17948_/A1 vssd1 vssd1 vccd1 vccd1 _17112_/A1 sky130_fd_sc_hd__buf_4
XFILLER_94_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16714_ _16719_/A _16714_/B _16714_/C _16714_/D vssd1 vssd1 vccd1 vccd1 _16715_/A
+ sky130_fd_sc_hd__or4_2
X_19502_ _21023_/CLK _19502_/D vssd1 vssd1 vccd1 vccd1 _19502_/Q sky130_fd_sc_hd__dfxtp_4
X_13926_ _19130_/Q _13906_/B _13903_/Y _13388_/A vssd1 vssd1 vccd1 vccd1 _19130_/D
+ sky130_fd_sc_hd__o22a_1
X_17694_ _20478_/Q _17903_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20478_/D sky130_fd_sc_hd__mux2_1
XFILLER_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19433_ _20565_/CLK _19433_/D vssd1 vssd1 vccd1 vccd1 _19433_/Q sky130_fd_sc_hd__dfxtp_1
X_16645_ _19902_/Q _17891_/A1 _16670_/S vssd1 vssd1 vccd1 vccd1 _19902_/D sky130_fd_sc_hd__mux2_1
XFILLER_263_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13857_ _13463_/B _13446_/B _09516_/Y _19659_/Q vssd1 vssd1 vccd1 vccd1 _13860_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19364_ _20719_/CLK _19364_/D vssd1 vssd1 vccd1 vccd1 _19364_/Q sky130_fd_sc_hd__dfxtp_1
X_12808_ _12906_/A _12808_/B vssd1 vssd1 vccd1 vccd1 _12809_/B sky130_fd_sc_hd__or2_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16576_ _19854_/Q _16576_/A2 _16576_/B1 input25/X vssd1 vssd1 vccd1 vccd1 _16577_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13788_ _13612_/A _13438_/Y _13596_/X _13595_/Y _16240_/A1 vssd1 vssd1 vccd1 vccd1
+ _13788_/X sky130_fd_sc_hd__a32o_4
XFILLER_43_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18315_ _18560_/B vssd1 vssd1 vccd1 vccd1 _18315_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_203_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15527_ _15527_/A _15527_/B vssd1 vssd1 vccd1 vccd1 _15527_/Y sky130_fd_sc_hd__nand2_1
XFILLER_231_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_32_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20660_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19295_ _20446_/CLK _19295_/D vssd1 vssd1 vccd1 vccd1 _19295_/Q sky130_fd_sc_hd__dfxtp_1
X_12739_ _12739_/A vssd1 vssd1 vccd1 vccd1 _12739_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18246_ _20803_/Q _18245_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18247_/B sky130_fd_sc_hd__mux2_1
XFILLER_124_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15458_ _15433_/X _15434_/X _15441_/X _15520_/B2 vssd1 vssd1 vccd1 vccd1 _15458_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14409_ _14437_/A _14437_/B _14409_/C vssd1 vssd1 vccd1 vccd1 _14409_/X sky130_fd_sc_hd__or3_1
X_18177_ _18422_/A _18177_/B vssd1 vssd1 vccd1 vccd1 _20789_/D sky130_fd_sc_hd__and2_1
X_15389_ _20954_/Q _15322_/C _15388_/X _15322_/B vssd1 vssd1 vccd1 vccd1 _15389_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17128_ _20096_/Q _17930_/A1 _17132_/S vssd1 vssd1 vccd1 vccd1 _20096_/D sky130_fd_sc_hd__mux2_1
XFILLER_237_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09950_ _19949_/Q _11895_/B vssd1 vssd1 vccd1 vccd1 _09950_/X sky130_fd_sc_hd__or2_1
X_17059_ _20031_/Q _17686_/A1 _17076_/S vssd1 vssd1 vccd1 vccd1 _20031_/D sky130_fd_sc_hd__mux2_1
X_20070_ _20573_/CLK _20070_/D vssd1 vssd1 vccd1 vccd1 _20070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09881_ _12120_/A1 _19483_/Q _19451_/Q _11916_/S _11892_/C1 vssd1 vssd1 vccd1 vccd1
+ _09881_/X sky130_fd_sc_hd__a221o_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20972_ _21041_/CLK _20972_/D vssd1 vssd1 vccd1 vccd1 _20972_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20406_ _20666_/CLK _20406_/D vssd1 vssd1 vccd1 vccd1 _20406_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20337_ _20667_/CLK _20337_/D vssd1 vssd1 vccd1 vccd1 _20337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11070_ _12306_/A1 _12371_/A1 _19336_/Q _12302_/S vssd1 vssd1 vccd1 vccd1 _11070_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_277_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20268_ _20268_/CLK _20268_/D vssd1 vssd1 vccd1 vccd1 _20268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10021_ _09612_/X _09636_/B _10020_/Y vssd1 vssd1 vccd1 vccd1 _10021_/Y sky130_fd_sc_hd__a21oi_1
Xinput102 dout0[63] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_hd__clkbuf_2
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput113 dout1[15] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20199_ _20727_/CLK _20199_/D vssd1 vssd1 vccd1 vccd1 _20199_/Q sky130_fd_sc_hd__dfxtp_1
Xinput124 dout1[25] vssd1 vssd1 vccd1 vccd1 input124/X sky130_fd_sc_hd__clkbuf_2
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput135 dout1[35] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__clkbuf_2
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput146 dout1[45] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__clkbuf_2
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput157 dout1[55] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__clkbuf_2
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 dout1[7] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput179 irq[2] vssd1 vssd1 vccd1 vccd1 _12548_/C sky130_fd_sc_hd__clkbuf_4
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _19127_/Q _14764_/A2 _14759_/X _18352_/C1 vssd1 vssd1 vccd1 vccd1 _19504_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11972_ _11970_/X _11971_/X _11995_/S vssd1 vssd1 vccd1 vccd1 _11972_/X sky130_fd_sc_hd__mux2_1
XFILLER_263_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13711_ _13780_/A _13711_/B vssd1 vssd1 vccd1 vccd1 _13711_/X sky130_fd_sc_hd__and2_1
X_10923_ _10920_/X _10921_/X _10922_/X _11170_/B1 _12302_/S vssd1 vssd1 vccd1 vccd1
+ _10923_/X sky130_fd_sc_hd__o221a_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _19450_/Q _17940_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19450_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16430_ _19756_/Q _16428_/B _16429_/Y vssd1 vssd1 vccd1 vccd1 _19756_/D sky130_fd_sc_hd__o21a_1
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _13642_/A vssd1 vssd1 vccd1 vccd1 _13666_/B sky130_fd_sc_hd__inv_6
X_10854_ _19803_/Q _12255_/A2 _10852_/X _09738_/A _10853_/X vssd1 vssd1 vccd1 vccd1
+ _10854_/X sky130_fd_sc_hd__o221a_1
XFILLER_147_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _19730_/Q _16362_/C _19731_/Q vssd1 vssd1 vccd1 vccd1 _16363_/B sky130_fd_sc_hd__a21oi_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _12664_/C _13572_/X _12982_/B vssd1 vssd1 vccd1 vccd1 _13573_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_9_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _12265_/A _10784_/Y _10781_/Y _12431_/A1 vssd1 vssd1 vccd1 vccd1 _10785_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18100_ _20774_/Q _18101_/C _20775_/Q vssd1 vssd1 vccd1 vccd1 _18102_/B sky130_fd_sc_hd__a21oi_1
X_15312_ _09479_/Y _14972_/B _14971_/B vssd1 vssd1 vccd1 vccd1 _15312_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12524_ _18763_/A1 _09498_/Y _18598_/A _12523_/X vssd1 vssd1 vccd1 vccd1 _13479_/A
+ sky130_fd_sc_hd__a211oi_4
X_19080_ _20425_/Q vssd1 vssd1 vccd1 vccd1 _20425_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _19705_/Q _16294_/C _16381_/B1 vssd1 vssd1 vccd1 vccd1 _16293_/B sky130_fd_sc_hd__o21ai_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18031_ _18112_/A _18036_/C vssd1 vssd1 vccd1 vccd1 _18031_/Y sky130_fd_sc_hd__nor2_1
X_15243_ _15021_/A _15230_/X _15242_/X vssd1 vssd1 vccd1 vccd1 _15243_/X sky130_fd_sc_hd__a21o_4
X_12455_ _12464_/A _12510_/C _13863_/A vssd1 vssd1 vccd1 vccd1 _12455_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_157_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11406_ _13459_/A _13611_/A _11766_/B vssd1 vssd1 vccd1 vccd1 _11406_/X sky130_fd_sc_hd__or3_1
X_15174_ _15155_/S _15038_/X _15173_/Y vssd1 vssd1 vccd1 vccd1 _15174_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12386_ _12396_/A1 _20523_/Q _12391_/S _12378_/X vssd1 vssd1 vccd1 vccd1 _12386_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14125_ _14122_/Y _14124_/X _13552_/A _12529_/X vssd1 vssd1 vccd1 vccd1 _14126_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11337_ _19470_/Q _09695_/Y _11336_/X _12377_/S vssd1 vssd1 vccd1 vccd1 _11337_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19982_ _20862_/CLK _19982_/D vssd1 vssd1 vccd1 vccd1 _19982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_150_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21023_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14056_ _19187_/Q _14108_/A2 _14055_/X _14458_/A vssd1 vssd1 vccd1 vccd1 _19187_/D
+ sky130_fd_sc_hd__o211a_1
X_18933_ _19109_/Q _18954_/A2 _18967_/B1 _13439_/C vssd1 vssd1 vccd1 vccd1 _18934_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ _11268_/A _20054_/Q _11268_/C vssd1 vssd1 vccd1 vccd1 _11268_/X sky130_fd_sc_hd__and3_1
XFILLER_141_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _20975_/Q _20909_/Q vssd1 vssd1 vccd1 vccd1 _13007_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10219_ _11336_/A _10217_/X _10218_/X vssd1 vssd1 vccd1 vccd1 _10219_/X sky130_fd_sc_hd__o21a_1
X_11199_ _11197_/X _11198_/X _12414_/S vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18864_ _19099_/Q _18864_/A2 _18864_/B1 _13426_/A vssd1 vssd1 vccd1 vccd1 _18865_/B
+ sky130_fd_sc_hd__a22o_1
X_17815_ _20590_/Q _17887_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20590_/D sky130_fd_sc_hd__mux2_1
X_18795_ _18795_/A _18795_/B vssd1 vssd1 vccd1 vccd1 _20984_/D sky130_fd_sc_hd__nor2_1
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17746_ _20525_/Q _17886_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20525_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14958_ _14958_/A _14973_/B _14966_/C vssd1 vssd1 vccd1 vccd1 _14959_/B sky130_fd_sc_hd__or3_1
XFILLER_242_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _13909_/A _13919_/S vssd1 vssd1 vccd1 vccd1 _13909_/Y sky130_fd_sc_hd__nand2_1
X_17677_ _20461_/Q _17780_/A1 _17706_/S vssd1 vssd1 vccd1 vccd1 _20461_/D sky130_fd_sc_hd__mux2_1
X_14889_ _14841_/S _14888_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _14889_/X sky130_fd_sc_hd__o21a_2
XFILLER_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19416_ _20716_/CLK _19416_/D vssd1 vssd1 vccd1 vccd1 _19416_/Q sky130_fd_sc_hd__dfxtp_1
X_16628_ _19887_/Q _17802_/A1 _16632_/S vssd1 vssd1 vccd1 vccd1 _19887_/D sky130_fd_sc_hd__mux2_1
XFILLER_196_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16559_ _16593_/A _16559_/B vssd1 vssd1 vccd1 vccd1 _19845_/D sky130_fd_sc_hd__or2_1
X_19347_ _20702_/CLK _19347_/D vssd1 vssd1 vccd1 vccd1 _19347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19278_ _20669_/CLK _19278_/D vssd1 vssd1 vccd1 vccd1 _19278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18229_ _18223_/B _14259_/B _18228_/Y vssd1 vssd1 vccd1 vccd1 _18508_/B sky130_fd_sc_hd__o21ai_4
XFILLER_175_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20122_ _20561_/CLK _20122_/D vssd1 vssd1 vccd1 vccd1 _20122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09933_ _09929_/X _09932_/X _11949_/S vssd1 vssd1 vccd1 vccd1 _09933_/X sky130_fd_sc_hd__mux2_1
Xfanout803 _17461_/X vssd1 vssd1 vccd1 vccd1 _17505_/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout814 _12563_/Y vssd1 vssd1 vccd1 vccd1 _13798_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout825 _14884_/X vssd1 vssd1 vccd1 vccd1 _15610_/B1 sky130_fd_sc_hd__clkbuf_16
X_20053_ _20085_/CLK _20053_/D vssd1 vssd1 vccd1 vccd1 _20053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout836 _18690_/Y vssd1 vssd1 vccd1 vccd1 _18719_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout847 _18343_/B vssd1 vssd1 vccd1 vccd1 _18349_/B sky130_fd_sc_hd__buf_6
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _11761_/A vssd1 vssd1 vccd1 vccd1 _13414_/A sky130_fd_sc_hd__inv_2
XFILLER_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout858 _15995_/A2 vssd1 vssd1 vccd1 vccd1 _16044_/A2 sky130_fd_sc_hd__buf_6
XFILLER_113_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout869 _14957_/X vssd1 vssd1 vccd1 vccd1 _15309_/S sky130_fd_sc_hd__buf_8
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09795_ _20579_/Q _12043_/B vssd1 vssd1 vccd1 vccd1 _09795_/X sky130_fd_sc_hd__or2_1
XFILLER_280_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_207 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_229 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20955_ _21019_/CLK _20955_/D vssd1 vssd1 vccd1 vccd1 _20955_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20949_/CLK _20886_/D vssd1 vssd1 vccd1 vccd1 _20886_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_81_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10570_ _12136_/B1 _10565_/X _10567_/X _10569_/X _12046_/B1 vssd1 vssd1 vccd1 vccd1
+ _10570_/X sky130_fd_sc_hd__o221a_1
XFILLER_194_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ _19296_/Q _20083_/Q _12316_/S vssd1 vssd1 vccd1 vccd1 _12240_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ _12189_/A _12171_/B vssd1 vssd1 vccd1 vccd1 _12171_/X sky130_fd_sc_hd__or2_1
XFILLER_163_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11122_ _11118_/A _11121_/Y _11118_/Y _11384_/S vssd1 vssd1 vccd1 vccd1 _11122_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11053_ _15545_/A _11054_/B vssd1 vssd1 vccd1 vccd1 _11053_/Y sky130_fd_sc_hd__nor2_2
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15930_ _15219_/Y _15925_/Y _15926_/Y _15929_/X vssd1 vssd1 vccd1 vccd1 _15930_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10004_ _19682_/Q _20170_/Q _11944_/S vssd1 vssd1 vccd1 vccd1 _10004_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15861_ _15882_/A1 _15850_/X _15851_/X _15860_/X vssd1 vssd1 vccd1 vccd1 _15861_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _20358_/Q _17911_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20358_/D sky130_fd_sc_hd__mux2_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _11412_/B _11737_/B _14815_/S vssd1 vssd1 vccd1 vccd1 _14812_/X sky130_fd_sc_hd__mux2_1
XFILLER_280_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _20918_/Q _18592_/B vssd1 vssd1 vccd1 vccd1 _18580_/Y sky130_fd_sc_hd__nand2_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _15258_/A _15406_/Y _15409_/B _14822_/S vssd1 vssd1 vccd1 vccd1 _15792_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_224_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17531_ _14483_/S _17528_/C _17537_/A vssd1 vssd1 vccd1 vccd1 _17532_/B sky130_fd_sc_hd__o21a_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _19496_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14743_/X sky130_fd_sc_hd__or2_1
XFILLER_83_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _11955_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _15887_/S sky130_fd_sc_hd__and2_4
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _11008_/A1 _19901_/Q _10924_/S _20026_/Q vssd1 vssd1 vccd1 vccd1 _10906_/X
+ sky130_fd_sc_hd__o22a_1
X_17462_ _20266_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17462_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14674_ _19433_/Q _17923_/A1 _14685_/S vssd1 vssd1 vccd1 vccd1 _19433_/D sky130_fd_sc_hd__mux2_1
XFILLER_260_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11886_ _12156_/A1 _11885_/X _11884_/X vssd1 vssd1 vccd1 vccd1 _11886_/X sky130_fd_sc_hd__a21o_1
X_19201_ _20659_/CLK _19201_/D vssd1 vssd1 vccd1 vccd1 _19201_/Q sky130_fd_sc_hd__dfxtp_1
X_16413_ _16451_/A _16418_/C vssd1 vssd1 vccd1 vccd1 _16413_/Y sky130_fd_sc_hd__nor2_1
X_13625_ _13481_/A _13411_/A _13414_/Y _16598_/C vssd1 vssd1 vccd1 vccd1 _13625_/Y
+ sky130_fd_sc_hd__o2bb2ai_4
X_10837_ _19371_/Q _20662_/Q _12316_/S vssd1 vssd1 vccd1 vccd1 _10837_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17393_ _20245_/Q _17401_/A2 _17392_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _20245_/D
+ sky130_fd_sc_hd__o211a_1
X_19132_ _19232_/CLK _19132_/D vssd1 vssd1 vccd1 vccd1 _19132_/Q sky130_fd_sc_hd__dfxtp_1
X_16344_ _19724_/Q _16346_/C _16343_/Y vssd1 vssd1 vccd1 vccd1 _19724_/D sky130_fd_sc_hd__o21a_1
XFILLER_186_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13556_ _13582_/A _19222_/Q vssd1 vssd1 vccd1 vccd1 _13556_/Y sky130_fd_sc_hd__nand2_1
X_10768_ _12411_/A _19308_/Q _12406_/C vssd1 vssd1 vccd1 vccd1 _10768_/X sky130_fd_sc_hd__or3_1
XFILLER_146_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ _12517_/C _12519_/A _12584_/B _11367_/A vssd1 vssd1 vccd1 vccd1 _12508_/B
+ sky130_fd_sc_hd__or4b_1
X_19063_ _20408_/Q vssd1 vssd1 vccd1 vccd1 _20408_/D sky130_fd_sc_hd__clkbuf_2
X_16275_ _19691_/Q _17949_/A1 _16275_/S vssd1 vssd1 vccd1 vccd1 _19691_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13487_ _13498_/B _13485_/Y _13486_/Y vssd1 vssd1 vccd1 vccd1 _13487_/Y sky130_fd_sc_hd__o21ai_1
X_10699_ _10697_/X _10698_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _10700_/B sky130_fd_sc_hd__mux2_1
XFILLER_185_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18014_ _18096_/A _18019_/C vssd1 vssd1 vccd1 vccd1 _18014_/Y sky130_fd_sc_hd__nor2_1
XFILLER_218_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15226_ _15226_/A _15226_/B vssd1 vssd1 vccd1 vccd1 _15226_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12438_ _13178_/A vssd1 vssd1 vccd1 vccd1 _12438_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput406 _13799_/X vssd1 vssd1 vccd1 vccd1 din0[8] sky130_fd_sc_hd__buf_4
Xoutput417 _19977_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[16] sky130_fd_sc_hd__buf_4
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput428 _19987_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[26] sky130_fd_sc_hd__buf_4
XFILLER_172_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15157_ _15157_/A vssd1 vssd1 vccd1 vccd1 _15157_/Y sky130_fd_sc_hd__inv_2
X_12369_ _12396_/A1 _19492_/Q _19460_/Q _12368_/S _12371_/C1 vssd1 vssd1 vccd1 vccd1
+ _12369_/X sky130_fd_sc_hd__a221o_1
Xoutput439 _19968_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[7] sky130_fd_sc_hd__buf_4
XFILLER_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14108_ _19213_/Q _14108_/A2 _14107_/X _17963_/B1 vssd1 vssd1 vccd1 vccd1 _19213_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15088_ _15081_/X _15087_/X _15142_/S vssd1 vssd1 vccd1 vccd1 _15088_/X sky130_fd_sc_hd__mux2_1
X_19965_ _20624_/CLK _19965_/D vssd1 vssd1 vccd1 vccd1 _19965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14039_ _19212_/Q _14105_/C _14039_/S vssd1 vssd1 vccd1 vccd1 _14039_/X sky130_fd_sc_hd__mux2_1
X_18916_ _21002_/Q _18971_/B vssd1 vssd1 vccd1 vccd1 _18916_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19896_ _20155_/CLK _19896_/D vssd1 vssd1 vccd1 vccd1 _19896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18847_ _20992_/Q _18861_/B vssd1 vssd1 vccd1 vccd1 _18847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09580_ _19115_/Q _19113_/Q _19112_/Q _19109_/Q vssd1 vssd1 vccd1 vccd1 _09580_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_83_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18778_ _19086_/Q _12589_/B _12592_/C _15127_/A _12533_/B vssd1 vssd1 vccd1 vccd1
+ _18778_/X sky130_fd_sc_hd__a221o_1
XFILLER_83_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17729_ _20510_/Q _17869_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20510_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20740_ _20862_/CLK _20740_/D vssd1 vssd1 vccd1 vccd1 _20740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20671_ _20671_/CLK _20671_/D vssd1 vssd1 vccd1 vccd1 _20671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout600 _14635_/X vssd1 vssd1 vccd1 vccd1 _14662_/S sky130_fd_sc_hd__clkbuf_8
Xfanout1609 _11094_/S vssd1 vssd1 vccd1 vccd1 _12301_/S sky130_fd_sc_hd__buf_6
X_20105_ _20708_/CLK _20105_/D vssd1 vssd1 vccd1 vccd1 _20105_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout611 _14531_/X vssd1 vssd1 vccd1 vccd1 _14560_/S sky130_fd_sc_hd__clkbuf_16
X_09916_ _20418_/Q _20354_/Q _20646_/Q _20610_/Q _12182_/S _11846_/C vssd1 vssd1 vccd1
+ vccd1 _09916_/X sky130_fd_sc_hd__mux4_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout622 _14116_/Y vssd1 vssd1 vccd1 vccd1 _14205_/A2 sky130_fd_sc_hd__buf_6
Xfanout633 _16822_/A vssd1 vssd1 vccd1 vccd1 _16985_/B1 sky130_fd_sc_hd__buf_12
Xfanout644 _16170_/S vssd1 vssd1 vccd1 vccd1 _16194_/S sky130_fd_sc_hd__buf_2
XFILLER_59_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout655 _15402_/A vssd1 vssd1 vccd1 vccd1 _15492_/A sky130_fd_sc_hd__buf_4
Xfanout666 _14108_/A2 vssd1 vssd1 vccd1 vccd1 _14104_/A2 sky130_fd_sc_hd__buf_4
X_20036_ _20315_/CLK _20036_/D vssd1 vssd1 vccd1 vccd1 _20036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout677 _14738_/B vssd1 vssd1 vccd1 vccd1 _13902_/B sky130_fd_sc_hd__buf_6
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09847_ _18765_/B _09842_/X _09846_/Y _15678_/A1 vssd1 vssd1 vccd1 vccd1 _09847_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout688 _14031_/A2 vssd1 vssd1 vccd1 vccd1 _14040_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_246_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout699 _14107_/A vssd1 vssd1 vccd1 vccd1 _14105_/A sky130_fd_sc_hd__buf_2
XFILLER_218_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09769_/X _09777_/Y _12192_/A1 _09761_/X vssd1 vssd1 vccd1 vccd1 _09778_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11742_/A _11742_/B vssd1 vssd1 vccd1 vccd1 _11741_/A sky130_fd_sc_hd__or2_4
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _21004_/CLK _20938_/D vssd1 vssd1 vccd1 vccd1 _20938_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _12059_/A1 _11670_/X _11667_/X _12059_/C1 vssd1 vssd1 vccd1 vccd1 _11671_/X
+ sky130_fd_sc_hd__a211o_1
X_20869_ _21043_/CLK _20869_/D vssd1 vssd1 vccd1 vccd1 _20869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ _14306_/A1 _19230_/Q _14772_/C1 _13409_/X vssd1 vssd1 vccd1 vccd1 _13411_/B
+ sky130_fd_sc_hd__o211a_1
X_10622_ _20127_/Q _20095_/Q _10622_/S vssd1 vssd1 vccd1 vccd1 _10622_/X sky130_fd_sc_hd__mux2_1
X_14390_ _19241_/Q _14398_/A2 _14389_/X _14780_/C1 vssd1 vssd1 vccd1 vccd1 _19241_/D
+ sky130_fd_sc_hd__o211a_1
X_13341_ _13340_/A _13340_/B _13355_/B vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__o21ba_1
X_10553_ _10553_/A _10553_/B _10553_/C _10553_/D vssd1 vssd1 vccd1 vccd1 _11150_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_139_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16060_ _15890_/A _16053_/Y _16059_/X _16056_/X vssd1 vssd1 vccd1 vccd1 _16060_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13272_ _20967_/Q _13272_/B vssd1 vssd1 vccd1 vccd1 _13272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _10482_/X _10483_/X _11256_/S vssd1 vssd1 vccd1 vccd1 _10484_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ _14938_/Y _15021_/C vssd1 vssd1 vccd1 vccd1 _15452_/S sky130_fd_sc_hd__nand2b_4
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12223_ _20147_/Q _20115_/Q _12375_/S vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12154_ _12366_/A1 _10041_/B _10037_/B vssd1 vssd1 vccd1 vccd1 _12154_/X sky130_fd_sc_hd__a21o_4
XFILLER_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _12411_/A _19304_/Q _12411_/C vssd1 vssd1 vccd1 vccd1 _11105_/X sky130_fd_sc_hd__or3_1
XFILLER_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19750_ _19978_/CLK _19750_/D vssd1 vssd1 vccd1 vccd1 _19750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16962_ _19986_/Q _17012_/A2 _16961_/Y _17012_/C1 vssd1 vssd1 vccd1 vccd1 _19986_/D
+ sky130_fd_sc_hd__a211o_1
X_12085_ _19392_/Q _12085_/A2 _12083_/X _12085_/B2 _12084_/X vssd1 vssd1 vccd1 vccd1
+ _12085_/X sky130_fd_sc_hd__o221a_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18701_ _20951_/Q _18185_/Y _18719_/S vssd1 vssd1 vccd1 vccd1 _18702_/B sky130_fd_sc_hd__mux2_1
XFILLER_265_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11036_ _12347_/A1 _19465_/Q _19433_/Q _11377_/S _11212_/S vssd1 vssd1 vccd1 vccd1
+ _11036_/X sky130_fd_sc_hd__a221o_1
XFILLER_209_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15913_ _16046_/A1 _15912_/X _15908_/X vssd1 vssd1 vccd1 vccd1 _15913_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16893_ input51/X input86/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16893_/X sky130_fd_sc_hd__mux2_8
X_19681_ _20708_/CLK _19681_/D vssd1 vssd1 vccd1 vccd1 _19681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15844_ _11883_/D _15925_/B _15219_/Y _15843_/Y vssd1 vssd1 vccd1 vccd1 _15844_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18632_ _19511_/Q _18671_/B vssd1 vssd1 vccd1 vccd1 _18632_/Y sky130_fd_sc_hd__nand2_1
XFILLER_264_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18563_ _18563_/A _18981_/B _18563_/C vssd1 vssd1 vccd1 vccd1 _18563_/X sky130_fd_sc_hd__or3_4
X_15775_ _20935_/Q _16044_/A2 _15774_/X vssd1 vssd1 vccd1 vccd1 _15775_/X sky130_fd_sc_hd__o21a_1
XFILLER_280_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _19225_/Q _19224_/Q _13587_/B vssd1 vssd1 vccd1 vccd1 _13449_/B sky130_fd_sc_hd__and3_1
XFILLER_217_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _19483_/Q _17941_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19483_/D sky130_fd_sc_hd__mux2_1
X_17514_ _20292_/Q _17522_/B vssd1 vssd1 vccd1 vccd1 _17514_/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18494_ _20891_/Q _18474_/S _18493_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18495_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_11938_ _11946_/A1 _20390_/Q _20454_/Q _11947_/S _12016_/C1 vssd1 vssd1 vccd1 vccd1
+ _11938_/X sky130_fd_sc_hd__a221o_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_560 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_571 _19841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_582 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17445_ _17421_/B _17446_/B _17457_/C _17438_/X vssd1 vssd1 vccd1 vccd1 _17445_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _19419_/Q _17801_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19419_/D sky130_fd_sc_hd__mux2_1
XANTENNA_593 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ _11946_/A1 _20389_/Q _20453_/Q _11944_/S vssd1 vssd1 vccd1 vccd1 _11869_/X
+ sky130_fd_sc_hd__a22o_1
X_13608_ _18604_/B _13606_/X _13607_/Y _13598_/Y _13603_/X vssd1 vssd1 vccd1 vccd1
+ _13609_/B sky130_fd_sc_hd__a32o_1
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17376_ _20236_/Q _17378_/A2 _17382_/B1 _20285_/Q _17380_/C1 vssd1 vssd1 vccd1 vccd1
+ _17376_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14588_ _19354_/Q _17940_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19354_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19115_ _20721_/CLK _19115_/D vssd1 vssd1 vccd1 vccd1 _19115_/Q sky130_fd_sc_hd__dfxtp_4
X_16327_ _19718_/Q _16330_/C _16451_/A vssd1 vssd1 vccd1 vccd1 _16327_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_199_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13539_ _13631_/B _13539_/B vssd1 vssd1 vccd1 vccd1 _13539_/Y sky130_fd_sc_hd__nor2_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19046_ _18310_/Y _19046_/A2 _19048_/B1 _12551_/B _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19046_/X sky130_fd_sc_hd__a221o_1
X_16258_ _19674_/Q _17689_/A1 _16275_/S vssd1 vssd1 vccd1 vccd1 _19674_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15209_ _11019_/Y _15208_/X _15402_/A vssd1 vssd1 vccd1 vccd1 _15209_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ _16189_/A _16189_/B vssd1 vssd1 vccd1 vccd1 _19618_/D sky130_fd_sc_hd__and2_1
XFILLER_160_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19948_ _20480_/CLK _19948_/D vssd1 vssd1 vccd1 vccd1 _19948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09701_ _11983_/A1 _19485_/Q _19453_/Q _11889_/S _11892_/C1 vssd1 vssd1 vccd1 vccd1
+ _09701_/X sky130_fd_sc_hd__a221o_1
XFILLER_96_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19879_ _20557_/CLK _19879_/D vssd1 vssd1 vccd1 vccd1 _19879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_261_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09632_ _09630_/X _09632_/B vssd1 vssd1 vccd1 vccd1 _09632_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09563_ _12464_/A _12468_/B _11268_/C vssd1 vssd1 vccd1 vccd1 _14898_/A sky130_fd_sc_hd__and3b_4
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09494_ _19121_/Q vssd1 vssd1 vccd1 vccd1 _09494_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20723_ _20794_/CLK _20723_/D vssd1 vssd1 vccd1 vccd1 _20723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20654_ _20686_/CLK _20654_/D vssd1 vssd1 vccd1 vccd1 _20654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20585_ _20585_/CLK _20585_/D vssd1 vssd1 vccd1 vccd1 _20585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1406 _10345_/S vssd1 vssd1 vccd1 vccd1 _11292_/S0 sky130_fd_sc_hd__buf_6
Xfanout1417 fanout1422/X vssd1 vssd1 vccd1 vccd1 _11377_/S sky130_fd_sc_hd__buf_6
Xfanout1428 _12248_/B1 vssd1 vssd1 vccd1 vccd1 _12339_/S0 sky130_fd_sc_hd__buf_6
XFILLER_278_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1439 _09735_/Y vssd1 vssd1 vccd1 vccd1 _15129_/A0 sky130_fd_sc_hd__buf_6
XFILLER_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20019_ _20273_/CLK _20019_/D vssd1 vssd1 vccd1 vccd1 _20019_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12910_ _13116_/A _13116_/B _13116_/C _12629_/Y vssd1 vssd1 vccd1 vccd1 _13106_/C
+ sky130_fd_sc_hd__a211o_1
Xfanout496 _17851_/X vssd1 vssd1 vccd1 vccd1 _17880_/S sky130_fd_sc_hd__buf_12
XFILLER_207_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13890_ _19108_/Q _14040_/A2 _13896_/B1 _10831_/S _13890_/C1 vssd1 vssd1 vccd1 vccd1
+ _19108_/D sky130_fd_sc_hd__o221a_1
XFILLER_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12841_ _13300_/B _12842_/D vssd1 vssd1 vccd1 vccd1 _13321_/A sky130_fd_sc_hd__nand2_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _19540_/Q _15591_/A _15558_/X _15559_/X _16167_/C1 vssd1 vssd1 vccd1 vccd1
+ _19540_/D sky130_fd_sc_hd__o221a_1
XFILLER_243_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _19501_/Q _12639_/A _19502_/Q vssd1 vssd1 vccd1 vccd1 _12773_/B sky130_fd_sc_hd__a21oi_1
XFILLER_215_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _19289_/Q _17874_/A1 _14516_/S vssd1 vssd1 vccd1 vccd1 _19289_/D sky130_fd_sc_hd__mux2_1
XFILLER_215_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11723_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11723_/Y sky130_fd_sc_hd__nand2_2
XFILLER_9_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _19505_/Q _15589_/S _15490_/X vssd1 vssd1 vccd1 vccd1 _15492_/B sky130_fd_sc_hd__o21ai_4
XFILLER_261_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17230_ _17441_/A _17423_/D _17441_/C vssd1 vssd1 vccd1 vccd1 _17230_/Y sky130_fd_sc_hd__nand3_4
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14442_ _14443_/B _17337_/A vssd1 vssd1 vccd1 vccd1 _17526_/B sky130_fd_sc_hd__nor2_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11654_ _20543_/Q _11682_/S vssd1 vssd1 vccd1 vccd1 _11654_/X sky130_fd_sc_hd__or2_1
XFILLER_168_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10605_ _09834_/A _19906_/Q _10622_/S _20031_/Q vssd1 vssd1 vccd1 vccd1 _10605_/X
+ sky130_fd_sc_hd__o22a_1
X_17161_ _20127_/Q _17686_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20127_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14373_ _19519_/Q _14373_/B vssd1 vssd1 vccd1 vccd1 _14374_/B sky130_fd_sc_hd__nand2_1
XFILLER_168_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11585_ _20544_/Q _11965_/B vssd1 vssd1 vccd1 vccd1 _11585_/X sky130_fd_sc_hd__or2_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16112_ _09867_/X _16132_/A2 _16111_/X vssd1 vssd1 vccd1 vccd1 _19580_/D sky130_fd_sc_hd__o21a_1
XFILLER_155_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13324_ _20932_/Q _13350_/B _13323_/X _18671_/B vssd1 vssd1 vccd1 vccd1 _13324_/X
+ sky130_fd_sc_hd__a211o_1
X_17092_ _20062_/Q _17894_/A1 _17114_/S vssd1 vssd1 vccd1 vccd1 _20062_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _10530_/X _10535_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _10536_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16043_ _20913_/Q _16043_/A2 _16043_/B1 _16040_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _16043_/X sky130_fd_sc_hd__a221o_1
X_13255_ _19238_/Q _13255_/B vssd1 vssd1 vccd1 vccd1 _13255_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ input125/X input160/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__mux2_8
XFILLER_124_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12206_ _13432_/A _12206_/B _12206_/C vssd1 vssd1 vccd1 vccd1 _12207_/B sky130_fd_sc_hd__or3_1
XFILLER_142_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20563_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13186_ _19299_/Q _13631_/B vssd1 vssd1 vccd1 vccd1 _16066_/B sky130_fd_sc_hd__or2_4
X_10398_ _15649_/A1 _10397_/X _10396_/X vssd1 vssd1 vccd1 vccd1 _10398_/X sky130_fd_sc_hd__o21a_1
X_19802_ _20667_/CLK _19802_/D vssd1 vssd1 vccd1 vccd1 _19802_/Q sky130_fd_sc_hd__dfxtp_1
X_12137_ _12137_/A1 _12129_/X _12135_/X _12136_/Y _12137_/C1 vssd1 vssd1 vccd1 vccd1
+ _12137_/X sky130_fd_sc_hd__a221o_1
X_17994_ _20736_/Q _17997_/C vssd1 vssd1 vccd1 vccd1 _17995_/B sky130_fd_sc_hd__and2_1
XFILLER_97_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1940 _13890_/C1 vssd1 vssd1 vccd1 vccd1 _16107_/B1 sky130_fd_sc_hd__buf_4
X_19733_ _21020_/CLK _19733_/D vssd1 vssd1 vccd1 vccd1 _19733_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16945_ _20624_/Q _16945_/B _16945_/C vssd1 vssd1 vccd1 vccd1 _16945_/X sky130_fd_sc_hd__and3_4
X_12068_ _09806_/S _12067_/X _12066_/X _12068_/C1 vssd1 vssd1 vccd1 vccd1 _12068_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout1951 _16381_/B1 vssd1 vssd1 vccd1 vccd1 _17331_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_238_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1962 _18960_/A vssd1 vssd1 vccd1 vccd1 _18932_/A sky130_fd_sc_hd__buf_4
XFILLER_226_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1973 _18877_/A vssd1 vssd1 vccd1 vccd1 _18096_/A sky130_fd_sc_hd__buf_2
Xfanout1984 _18808_/A vssd1 vssd1 vccd1 vccd1 _18783_/A sky130_fd_sc_hd__buf_4
X_11019_ _19497_/Q _11189_/B vssd1 vssd1 vccd1 vccd1 _11019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19664_ _20563_/CLK _19664_/D vssd1 vssd1 vccd1 vccd1 _19664_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1995 _18704_/A vssd1 vssd1 vccd1 vccd1 _18126_/A sky130_fd_sc_hd__buf_4
X_16876_ _16876_/A _16876_/B vssd1 vssd1 vccd1 vccd1 _16876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_237_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18615_ _20927_/Q _18619_/B vssd1 vssd1 vccd1 vccd1 _18615_/Y sky130_fd_sc_hd__nand2_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _21035_/Q _21003_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _15827_/X sky130_fd_sc_hd__mux2_1
X_19595_ _19621_/CLK _19595_/D vssd1 vssd1 vccd1 vccd1 _19595_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18546_ _18966_/A _18546_/B vssd1 vssd1 vccd1 vccd1 _20908_/D sky130_fd_sc_hd__nor2_1
X_15758_ _15948_/A1 _12811_/X _15757_/X _12832_/B vssd1 vssd1 vccd1 vccd1 _15760_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14709_ _19466_/Q _17924_/A1 _14719_/S vssd1 vssd1 vccd1 vccd1 _19466_/D sky130_fd_sc_hd__mux2_1
X_15689_ _20740_/Q _16041_/A2 _16041_/B1 _20772_/Q vssd1 vssd1 vccd1 vccd1 _15689_/X
+ sky130_fd_sc_hd__a22o_4
X_18477_ _18570_/B _18477_/B vssd1 vssd1 vccd1 vccd1 _18477_/X sky130_fd_sc_hd__or2_1
XANTENNA_390 _16860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17428_ _17432_/A _17428_/B vssd1 vssd1 vccd1 vccd1 _20258_/D sky130_fd_sc_hd__and2_1
XFILLER_220_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17359_ _20228_/Q _17363_/A2 _17358_/X _18700_/A vssd1 vssd1 vccd1 vccd1 _20228_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20370_ _20630_/CLK _20370_/D vssd1 vssd1 vccd1 vccd1 _20370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19029_ _21033_/Q _19049_/A2 _19028_/X _18740_/A vssd1 vssd1 vccd1 vccd1 _21033_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09615_ _12513_/D _10979_/C vssd1 vssd1 vccd1 vccd1 _09615_/Y sky130_fd_sc_hd__nand2_8
XFILLER_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09546_ _12580_/A _09556_/A vssd1 vssd1 vccd1 vccd1 _09546_/Y sky130_fd_sc_hd__nor2_4
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09477_ _09609_/A vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__inv_2
XPHY_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20706_ _20706_/CLK _20706_/D vssd1 vssd1 vccd1 vccd1 _20706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20637_ _20668_/CLK _20637_/D vssd1 vssd1 vccd1 vccd1 _20637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11370_ _12347_/A1 _19342_/Q _20697_/Q _11377_/S _12347_/C1 vssd1 vssd1 vccd1 vccd1
+ _11370_/X sky130_fd_sc_hd__a221o_1
XFILLER_137_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20568_ _20568_/CLK _20568_/D vssd1 vssd1 vccd1 vccd1 _20568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10321_ _19812_/Q _19316_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10321_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20499_ _20688_/CLK _20499_/D vssd1 vssd1 vccd1 vccd1 _20499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ _20958_/Q _20892_/Q vssd1 vssd1 vccd1 vccd1 _13315_/B sky130_fd_sc_hd__nand2_2
X_10252_ _10262_/A _19477_/Q _19445_/Q _11042_/B vssd1 vssd1 vccd1 vccd1 _10252_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ _11391_/A _19315_/Q _11391_/C vssd1 vssd1 vccd1 vccd1 _10183_/X sky130_fd_sc_hd__or3_1
XFILLER_278_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1203 _17331_/A2 vssd1 vssd1 vccd1 vccd1 _17268_/A2 sky130_fd_sc_hd__buf_4
Xfanout1214 _16133_/C vssd1 vssd1 vccd1 vccd1 _16052_/A1 sky130_fd_sc_hd__buf_4
XFILLER_267_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1225 _13305_/B vssd1 vssd1 vccd1 vccd1 _13519_/S sky130_fd_sc_hd__buf_4
Xfanout1236 _09683_/X vssd1 vssd1 vccd1 vccd1 split7/A sky130_fd_sc_hd__buf_12
XFILLER_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14991_ _14957_/B _15021_/B _14997_/C vssd1 vssd1 vccd1 vccd1 _14991_/X sky130_fd_sc_hd__o21a_1
Xfanout1247 _17336_/Y vssd1 vssd1 vccd1 vccd1 _17380_/C1 sky130_fd_sc_hd__buf_6
XFILLER_94_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1258 _12581_/B vssd1 vssd1 vccd1 vccd1 _16063_/A2 sky130_fd_sc_hd__buf_6
Xfanout1269 _09613_/B vssd1 vssd1 vccd1 vccd1 _18152_/C sky130_fd_sc_hd__clkbuf_4
X_16730_ _16822_/A _16730_/B vssd1 vssd1 vccd1 vccd1 _16730_/Y sky130_fd_sc_hd__nor2_1
X_13942_ _19145_/Q _13941_/B _13941_/Y _18752_/A vssd1 vssd1 vccd1 vccd1 _19145_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16661_ _19918_/Q _17835_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19918_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13873_ _19091_/Q _13953_/A2 _13881_/B1 _19157_/Q _16197_/A vssd1 vssd1 vccd1 vccd1
+ _19091_/D sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_175_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21008_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18400_ _18708_/A _18400_/B vssd1 vssd1 vccd1 vccd1 _20854_/D sky130_fd_sc_hd__and2_1
X_15612_ _14889_/X _15611_/X _15612_/S vssd1 vssd1 vccd1 vccd1 _15626_/B sky130_fd_sc_hd__mux2_2
XFILLER_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12824_ _19513_/Q _12835_/A vssd1 vssd1 vccd1 vccd1 _12824_/X sky130_fd_sc_hd__xor2_2
XFILLER_90_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16592_ _19862_/Q _16592_/A2 _16592_/B1 input34/X vssd1 vssd1 vccd1 vccd1 _16593_/B
+ sky130_fd_sc_hd__o22a_1
X_19380_ _20671_/CLK _19380_/D vssd1 vssd1 vccd1 vccd1 _19380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_262_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20856_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_222_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18331_ _18471_/B _18341_/B vssd1 vssd1 vccd1 vccd1 _18331_/Y sky130_fd_sc_hd__nand2_1
X_15543_ _16052_/A1 _15529_/X _15542_/Y _13426_/C _16052_/B2 vssd1 vssd1 vccd1 vccd1
+ _15544_/B sky130_fd_sc_hd__a32o_1
XFILLER_199_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12755_ _14803_/A1 _12582_/C _12784_/B _12754_/X vssd1 vssd1 vccd1 vccd1 _12755_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18728_/A _18262_/B vssd1 vssd1 vccd1 vccd1 _20806_/D sky130_fd_sc_hd__and2_1
X_11706_ _12105_/A _12023_/S _11703_/X _11705_/X vssd1 vssd1 vccd1 vccd1 _11706_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_202_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15474_ _15283_/A _15473_/Y _15096_/B vssd1 vssd1 vccd1 vccd1 _15474_/X sky130_fd_sc_hd__a21o_1
XFILLER_203_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12686_ _12686_/A _12686_/B _12686_/C vssd1 vssd1 vccd1 vccd1 _12692_/C sky130_fd_sc_hd__and3_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14425_ _14432_/A _14426_/C _14426_/D _14426_/A vssd1 vssd1 vccd1 vccd1 _14427_/B
+ sky130_fd_sc_hd__o22a_1
X_17213_ _20177_/Q _17704_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20177_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18193_ _19534_/Q _18213_/B vssd1 vssd1 vccd1 vccd1 _18193_/Y sky130_fd_sc_hd__nand2b_2
X_11637_ _12003_/C _11636_/X _11933_/S vssd1 vssd1 vccd1 vccd1 _11637_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17144_ _20112_/Q _17178_/A1 _17144_/S vssd1 vssd1 vccd1 vccd1 _20112_/D sky130_fd_sc_hd__mux2_1
X_14356_ _14356_/A _14361_/B vssd1 vssd1 vccd1 vccd1 _14356_/Y sky130_fd_sc_hd__nor2_1
X_11568_ _11568_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11568_/Y sky130_fd_sc_hd__nand2_4
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13307_ _13302_/X _13306_/X _13373_/A vssd1 vssd1 vccd1 vccd1 _13307_/Y sky130_fd_sc_hd__o21ai_2
X_10519_ _10517_/X _10518_/X _11304_/S vssd1 vssd1 vccd1 vccd1 _10519_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17075_ _20047_/Q _17945_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20047_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14287_ _19231_/Q _14398_/A2 _14286_/X _14776_/C1 vssd1 vssd1 vccd1 vccd1 _19231_/D
+ sky130_fd_sc_hd__o211a_1
X_11499_ _20541_/Q _12133_/S vssd1 vssd1 vccd1 vccd1 _11499_/X sky130_fd_sc_hd__or2_1
XFILLER_226_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16026_ _15264_/B _16058_/A2 _16026_/S vssd1 vssd1 vccd1 vccd1 _16026_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13238_ _20971_/Q _13370_/B _13237_/Y _18767_/A vssd1 vssd1 vccd1 vccd1 _13239_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13169_ _09941_/B _13415_/B _09941_/A vssd1 vssd1 vccd1 vccd1 _13414_/B sky130_fd_sc_hd__a21boi_4
XFILLER_112_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17977_ _18064_/A _17982_/C vssd1 vssd1 vccd1 vccd1 _17977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19716_ _20863_/CLK _19716_/D vssd1 vssd1 vccd1 vccd1 _19716_/Q sky130_fd_sc_hd__dfxtp_1
X_16928_ _19982_/Q _17012_/A2 _16927_/Y _18094_/A vssd1 vssd1 vccd1 vccd1 _19982_/D
+ sky130_fd_sc_hd__a211o_1
Xfanout1770 output482/A vssd1 vssd1 vccd1 vccd1 _13275_/A1 sky130_fd_sc_hd__buf_4
Xfanout1781 _20255_/Q vssd1 vssd1 vccd1 vccd1 _17402_/A sky130_fd_sc_hd__buf_6
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1792 _18199_/A1 vssd1 vssd1 vccd1 vccd1 _18148_/S sky130_fd_sc_hd__buf_6
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19647_ _20649_/CLK _19647_/D vssd1 vssd1 vccd1 vccd1 _19647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16859_ _19974_/Q _16887_/A _16858_/Y _16896_/C1 vssd1 vssd1 vccd1 vccd1 _19974_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_37_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19578_ _20341_/CLK _19578_/D vssd1 vssd1 vccd1 vccd1 _19578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18529_ _18651_/B _18529_/B vssd1 vssd1 vccd1 vccd1 _18529_/X sky130_fd_sc_hd__or2_2
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20422_ _20706_/CLK _20422_/D vssd1 vssd1 vccd1 vccd1 _20422_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_119_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20353_ _20353_/CLK _20353_/D vssd1 vssd1 vccd1 vccd1 _20353_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20284_ _21030_/CLK _20284_/D vssd1 vssd1 vccd1 vccd1 _20284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20580_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_275_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10870_ _10866_/A _10869_/Y _10866_/Y _12504_/A vssd1 vssd1 vccd1 vccd1 _10870_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_189_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _17452_/A vssd1 vssd1 vccd1 vccd1 _17457_/A sky130_fd_sc_hd__inv_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12540_ _20867_/Q _12548_/B _12540_/C vssd1 vssd1 vccd1 vccd1 _12552_/C sky130_fd_sc_hd__and3_2
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ _16054_/B _12471_/B vssd1 vssd1 vccd1 vccd1 _12471_/X sky130_fd_sc_hd__or2_4
XFILLER_185_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14210_ _14197_/Y _14201_/B _14199_/B vssd1 vssd1 vccd1 vccd1 _14211_/B sky130_fd_sc_hd__o21ai_4
X_11422_ _20574_/Q _11895_/B vssd1 vssd1 vccd1 vccd1 _11422_/X sky130_fd_sc_hd__or2_1
X_15190_ _20725_/Q _16041_/A2 _16041_/B1 _20757_/Q vssd1 vssd1 vccd1 vccd1 _15190_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14141_ _14141_/A _14141_/B vssd1 vssd1 vccd1 vccd1 _14141_/Y sky130_fd_sc_hd__xnor2_1
X_11353_ _12301_/S _11352_/X _11351_/X _11353_/C1 vssd1 vssd1 vccd1 vccd1 _11353_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_192_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10304_ _19412_/Q _20571_/Q _10485_/S vssd1 vssd1 vccd1 vccd1 _10304_/X sky130_fd_sc_hd__mux2_1
X_14072_ _19195_/Q _14104_/A2 _14071_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1 _19195_/D
+ sky130_fd_sc_hd__o211a_1
X_11284_ _11026_/A _19897_/Q _11292_/S0 _20022_/Q vssd1 vssd1 vccd1 vccd1 _11284_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_141_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17900_ _20671_/Q _17900_/A1 _17912_/S vssd1 vssd1 vccd1 vccd1 _20671_/D sky130_fd_sc_hd__mux2_1
X_13023_ _20967_/Q _20901_/Q vssd1 vssd1 vccd1 vccd1 _13270_/A sky130_fd_sc_hd__or2_2
X_10235_ _10233_/X _10234_/X _10235_/S vssd1 vssd1 vccd1 vccd1 _10235_/X sky130_fd_sc_hd__mux2_1
XFILLER_279_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18880_ _19134_/Q _18949_/A2 _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18880_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_133_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1000 _16000_/A1 vssd1 vssd1 vccd1 vccd1 _15882_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_121_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1011 _14881_/X vssd1 vssd1 vccd1 vccd1 _15259_/B sky130_fd_sc_hd__buf_4
XFILLER_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1022 _17004_/B1 vssd1 vssd1 vccd1 vccd1 _16870_/B1 sky130_fd_sc_hd__buf_4
X_17831_ _20606_/Q _17869_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20606_/D sky130_fd_sc_hd__mux2_1
X_10166_ _19411_/Q _20570_/Q _11042_/B vssd1 vssd1 vccd1 vccd1 _10166_/X sky130_fd_sc_hd__mux2_1
Xfanout1033 _16878_/A vssd1 vssd1 vccd1 vccd1 _16869_/A sky130_fd_sc_hd__buf_4
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1044 _16608_/A1 vssd1 vssd1 vccd1 vccd1 _17679_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_282_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1055 _17924_/A1 vssd1 vssd1 vccd1 vccd1 _17647_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 _11397_/B2 vssd1 vssd1 vccd1 vccd1 _12433_/B2 sky130_fd_sc_hd__buf_12
Xfanout1077 _18949_/B1 vssd1 vssd1 vccd1 vccd1 _18880_/B1 sky130_fd_sc_hd__buf_6
X_17762_ _20541_/Q _17902_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20541_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1088 _17674_/A1 vssd1 vssd1 vccd1 vccd1 _17708_/A1 sky130_fd_sc_hd__clkbuf_4
X_14974_ _15022_/A _14981_/A _15022_/B _14981_/B vssd1 vssd1 vccd1 vccd1 _14979_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_208_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10097_ _12084_/A _20669_/Q _12084_/C vssd1 vssd1 vccd1 vccd1 _10097_/X sky130_fd_sc_hd__or3_1
XFILLER_208_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19501_ _19696_/CLK _19501_/D vssd1 vssd1 vccd1 vccd1 _19501_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1099 _12156_/X vssd1 vssd1 vccd1 vccd1 _17948_/A1 sky130_fd_sc_hd__buf_4
X_16713_ _16945_/C _17219_/B vssd1 vssd1 vccd1 vccd1 _16713_/X sky130_fd_sc_hd__and2_2
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13925_ _19129_/Q _13921_/B _13932_/B1 _13361_/B vssd1 vssd1 vccd1 vccd1 _19129_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_267_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17693_ _20477_/Q _17693_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20477_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19432_ _20563_/CLK _19432_/D vssd1 vssd1 vccd1 vccd1 _19432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_262_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16644_ _19901_/Q _17750_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19901_/D sky130_fd_sc_hd__mux2_1
X_13856_ _19659_/Q _16232_/B _13854_/Y _13242_/B vssd1 vssd1 vccd1 vccd1 _16133_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_222_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ _12906_/A _12808_/B vssd1 vssd1 vccd1 vccd1 _13253_/A sky130_fd_sc_hd__nand2_1
X_19363_ _20718_/CLK _19363_/D vssd1 vssd1 vccd1 vccd1 _19363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16575_ _16593_/A _16575_/B vssd1 vssd1 vccd1 vccd1 _19853_/D sky130_fd_sc_hd__or2_1
X_13787_ _13612_/A _13438_/Y _15369_/A _13583_/Y _13244_/X vssd1 vssd1 vccd1 vccd1
+ _13787_/X sky130_fd_sc_hd__a32o_4
XFILLER_188_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10999_ _20400_/Q _11009_/A2 _10996_/X _10997_/X _10998_/X vssd1 vssd1 vccd1 vccd1
+ _10999_/X sky130_fd_sc_hd__o221a_1
XFILLER_16_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18314_ _18313_/B _14435_/A _18313_/Y vssd1 vssd1 vccd1 vccd1 _18560_/B sky130_fd_sc_hd__o21ai_4
XFILLER_204_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ _15526_/A _15526_/B vssd1 vssd1 vccd1 vccd1 _15526_/Y sky130_fd_sc_hd__nor2_2
X_12738_ _15528_/A _12738_/B vssd1 vssd1 vccd1 vccd1 _12739_/A sky130_fd_sc_hd__nor2_1
XFILLER_203_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _20081_/CLK _19294_/D vssd1 vssd1 vccd1 vccd1 _19294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18245_ _18517_/B vssd1 vssd1 vccd1 vccd1 _18245_/Y sky130_fd_sc_hd__inv_2
X_15457_ _15283_/A _15443_/Y _15457_/B1 vssd1 vssd1 vccd1 vccd1 _15457_/Y sky130_fd_sc_hd__a21oi_1
X_12669_ _12667_/X _12668_/X _12708_/B vssd1 vssd1 vccd1 vccd1 _12674_/B sky130_fd_sc_hd__a21o_1
X_14408_ _09488_/A _13119_/X _13124_/B _14407_/X vssd1 vssd1 vccd1 vccd1 _14409_/C
+ sky130_fd_sc_hd__a31o_1
X_18176_ _20789_/Q _18175_/Y _18236_/S vssd1 vssd1 vccd1 vccd1 _18177_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_72_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20633_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15388_ _15387_/X _20826_/Q _15388_/S vssd1 vssd1 vccd1 vccd1 _15388_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14339_ _19236_/Q _14438_/A2 _14338_/X _14794_/C1 vssd1 vssd1 vccd1 vccd1 _19236_/D
+ sky130_fd_sc_hd__o211a_1
X_17127_ _20095_/Q _17686_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20095_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17058_ _20030_/Q _17058_/A1 _17080_/S vssd1 vssd1 vccd1 vccd1 _20030_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16009_ _16009_/A _16009_/B vssd1 vssd1 vccd1 vccd1 _16009_/X sky130_fd_sc_hd__and2_1
XFILLER_103_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09880_ _19886_/Q _19787_/Q _11916_/S vssd1 vssd1 vccd1 vccd1 _09880_/X sky130_fd_sc_hd__mux2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20971_ _21040_/CLK _20971_/D vssd1 vssd1 vccd1 vccd1 _20971_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20405_ _21044_/CLK _20405_/D vssd1 vssd1 vccd1 vccd1 _20405_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_147_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20336_ _20690_/CLK _20336_/D vssd1 vssd1 vccd1 vccd1 _20336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20267_ _21022_/CLK _20267_/D vssd1 vssd1 vccd1 vccd1 _20267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10020_ _11235_/A _10020_/B vssd1 vssd1 vccd1 vccd1 _10020_/Y sky130_fd_sc_hd__nor2_2
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput103 dout0[6] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_hd__clkbuf_2
X_20198_ _20688_/CLK _20198_/D vssd1 vssd1 vccd1 vccd1 _20198_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput114 dout1[16] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput125 dout1[26] vssd1 vssd1 vccd1 vccd1 input125/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput136 dout1[36] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__clkbuf_2
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput147 dout1[46] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput158 dout1[56] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__clkbuf_2
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput169 dout1[8] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11971_ _19689_/Q _20177_/Q _11978_/S vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__mux2_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13710_ _13776_/B1 _13747_/B _13709_/X vssd1 vssd1 vccd1 vccd1 _13711_/B sky130_fd_sc_hd__a21oi_4
X_10922_ _20369_/Q _20433_/Q _10983_/S vssd1 vssd1 vccd1 vccd1 _10922_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _19449_/Q _17939_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19449_/D sky130_fd_sc_hd__mux2_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13641_ _13653_/A _13641_/B vssd1 vssd1 vccd1 vccd1 _13642_/A sky130_fd_sc_hd__nand2_2
X_10853_ _12337_/A _19307_/Q _12337_/C vssd1 vssd1 vccd1 vccd1 _10853_/X sky130_fd_sc_hd__or3_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _19730_/Q _16362_/C _16359_/Y vssd1 vssd1 vccd1 vccd1 _19730_/D sky130_fd_sc_hd__o21a_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13586_/C _13572_/B vssd1 vssd1 vccd1 vccd1 _13572_/X sky130_fd_sc_hd__or2_1
X_10784_ _12420_/B1 _10782_/X _10783_/X vssd1 vssd1 vccd1 vccd1 _10784_/Y sky130_fd_sc_hd__o21ai_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _20824_/Q _14965_/X _14972_/B _15310_/X vssd1 vssd1 vccd1 vccd1 _15311_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_197_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12523_ _14110_/A _12521_/Y _12522_/Y _13552_/A vssd1 vssd1 vccd1 vccd1 _12523_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_158_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _19705_/Q _16294_/C vssd1 vssd1 vccd1 vccd1 _16293_/A sky130_fd_sc_hd__and2_1
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _19706_/Q _15241_/X _15454_/S vssd1 vssd1 vccd1 vccd1 _15242_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18030_ _20749_/Q _20748_/Q _18030_/C vssd1 vssd1 vccd1 vccd1 _18036_/C sky130_fd_sc_hd__and3_4
X_12454_ _12454_/A _12454_/B _12454_/C vssd1 vssd1 vccd1 vccd1 _12454_/Y sky130_fd_sc_hd__nor3_1
XFILLER_200_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11405_ _11405_/A _11772_/B vssd1 vssd1 vccd1 vccd1 _11405_/X sky130_fd_sc_hd__or2_1
X_15173_ _15155_/S _15036_/X _15254_/S vssd1 vssd1 vccd1 vccd1 _15173_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ _09502_/A _12377_/X _12383_/X _12384_/Y _12385_/C1 vssd1 vssd1 vccd1 vccd1
+ _12385_/X sky130_fd_sc_hd__a221o_2
XFILLER_153_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14124_ _19494_/Q _14123_/B _14202_/S _13552_/A vssd1 vssd1 vccd1 vccd1 _14124_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11336_ _11336_/A _19438_/Q _11342_/S vssd1 vssd1 vccd1 vccd1 _11336_/X sky130_fd_sc_hd__and3_1
X_19981_ _20014_/CLK _19981_/D vssd1 vssd1 vccd1 vccd1 _19981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14055_ _14107_/A _14107_/B _14055_/C vssd1 vssd1 vccd1 vccd1 _14055_/X sky130_fd_sc_hd__or3_1
XFILLER_137_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18932_ _18932_/A _18932_/B vssd1 vssd1 vccd1 vccd1 _21004_/D sky130_fd_sc_hd__nor2_1
XFILLER_180_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11267_ _19366_/Q _09689_/D _11265_/X _11274_/B2 _11266_/X vssd1 vssd1 vccd1 vccd1
+ _11267_/X sky130_fd_sc_hd__o221a_1
XFILLER_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13006_ _20976_/Q _20910_/Q vssd1 vssd1 vccd1 vccd1 _13091_/B sky130_fd_sc_hd__or2_1
XFILLER_279_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10218_ _11258_/A1 _19349_/Q _20704_/Q _10217_/S _11338_/A1 vssd1 vssd1 vccd1 vccd1
+ _10218_/X sky130_fd_sc_hd__a221o_1
XFILLER_239_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18863_ _18863_/A _18863_/B vssd1 vssd1 vccd1 vccd1 _20994_/D sky130_fd_sc_hd__nor2_1
XFILLER_122_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11198_ _20398_/Q _20334_/Q _20626_/Q _20590_/Q _12339_/S0 _12254_/C vssd1 vssd1
+ vccd1 vccd1 _11198_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_190_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19609_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17814_ _20589_/Q _17852_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20589_/D sky130_fd_sc_hd__mux2_1
X_10149_ _11170_/B1 _10148_/X _10147_/X _09688_/A vssd1 vssd1 vccd1 vccd1 _10149_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18794_ _18477_/X _18819_/B _18792_/X _18793_/Y vssd1 vssd1 vccd1 vccd1 _18795_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17745_ _17745_/A _17851_/B _17745_/C vssd1 vssd1 vccd1 vccd1 _17745_/X sky130_fd_sc_hd__and3_4
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14957_ _15308_/C _14957_/B vssd1 vssd1 vccd1 vccd1 _14957_/X sky130_fd_sc_hd__and2_1
XFILLER_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13908_ _19119_/Q _13921_/B _13907_/Y _14758_/C1 vssd1 vssd1 vccd1 vccd1 _19119_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_236_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17676_ _17745_/A _17676_/B _17676_/C vssd1 vssd1 vccd1 vccd1 _17676_/X sky130_fd_sc_hd__and3_4
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14888_ _14885_/B _14887_/X _15357_/S vssd1 vssd1 vccd1 vccd1 _14888_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19415_ _20574_/CLK _19415_/D vssd1 vssd1 vccd1 vccd1 _19415_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_262_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16627_ _19886_/Q _17801_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19886_/D sky130_fd_sc_hd__mux2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13839_ _20261_/Q _20260_/Q _20259_/Q _13839_/D vssd1 vssd1 vccd1 vccd1 _13839_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_223_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19346_ _20701_/CLK _19346_/D vssd1 vssd1 vccd1 vccd1 _19346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16558_ _19845_/Q _16576_/A2 _16576_/B1 input15/X vssd1 vssd1 vccd1 vccd1 _16559_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15509_ _20894_/Q _15937_/A2 _15566_/B1 _15508_/X _15937_/C1 vssd1 vssd1 vccd1 vccd1
+ _15509_/X sky130_fd_sc_hd__a221o_1
X_19277_ _20671_/CLK _19277_/D vssd1 vssd1 vccd1 vccd1 _19277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16489_ _16672_/A _17744_/A vssd1 vssd1 vccd1 vccd1 _16490_/C sky130_fd_sc_hd__nor2_1
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18228_ _19541_/Q _18248_/B vssd1 vssd1 vccd1 vccd1 _18228_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ _18163_/A _14123_/B _18158_/Y vssd1 vssd1 vccd1 vccd1 _18459_/B sky130_fd_sc_hd__o21ai_4
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20121_ _20565_/CLK _20121_/D vssd1 vssd1 vccd1 vccd1 _20121_/Q sky130_fd_sc_hd__dfxtp_1
X_09932_ _11948_/A1 _09931_/X _09930_/X vssd1 vssd1 vccd1 vccd1 _09932_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout804 _17495_/A1 vssd1 vssd1 vccd1 vccd1 _17487_/A1 sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_207_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20677_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout815 _13740_/B vssd1 vssd1 vccd1 vccd1 _13655_/A sky130_fd_sc_hd__buf_8
X_20052_ _20084_/CLK _20052_/D vssd1 vssd1 vccd1 vccd1 _20052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout826 _14884_/X vssd1 vssd1 vccd1 vccd1 _15548_/B1 sky130_fd_sc_hd__buf_4
Xfanout837 _18690_/Y vssd1 vssd1 vccd1 vccd1 _18707_/S sky130_fd_sc_hd__buf_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _09863_/A _09863_/B vssd1 vssd1 vccd1 vccd1 _11761_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout848 _18343_/B vssd1 vssd1 vccd1 vccd1 _18341_/B sky130_fd_sc_hd__buf_6
XFILLER_259_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 _15337_/A2 vssd1 vssd1 vccd1 vccd1 _15995_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_133_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09794_ _12060_/A1 _19484_/Q _19452_/Q _10426_/S _12051_/C1 vssd1 vssd1 vccd1 vccd1
+ _09794_/X sky130_fd_sc_hd__a221o_1
XFILLER_246_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_208 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20954_ _21018_/CLK _20954_/D vssd1 vssd1 vccd1 vccd1 _20954_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_219 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20885_ _21019_/CLK _20885_/D vssd1 vssd1 vccd1 vccd1 _20885_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12170_ _20489_/Q _20329_/Q _12174_/S vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__mux2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ _12357_/A1 _11119_/X _11120_/X vssd1 vssd1 vccd1 vccd1 _11121_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20319_ _20479_/CLK _20319_/D vssd1 vssd1 vccd1 vccd1 _20319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11052_ _15407_/S _11054_/B vssd1 vssd1 vccd1 vccd1 _11052_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10003_ _09776_/S _09998_/Y _10002_/Y _12020_/C1 vssd1 vssd1 vccd1 vccd1 _10003_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_277_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _19758_/Q _15999_/A2 _15859_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15860_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14811_ _11411_/B _11733_/B _14815_/S vssd1 vssd1 vccd1 vccd1 _14811_/X sky130_fd_sc_hd__mux2_1
XFILLER_264_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _09862_/A _15984_/A2 _15984_/B1 _09863_/A _15890_/A vssd1 vssd1 vccd1 vccd1
+ _15791_/X sky130_fd_sc_hd__a221o_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _20299_/Q _17530_/A2 _17529_/X vssd1 vssd1 vccd1 vccd1 _17537_/B sky130_fd_sc_hd__a21o_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14742_ _19118_/Q _14802_/A2 _14741_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _19495_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11954_ _11955_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__nor2_1
XFILLER_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _19627_/Q _09689_/D _10902_/X _10903_/X _10904_/X vssd1 vssd1 vccd1 vccd1
+ _10905_/X sky130_fd_sc_hd__o221a_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14673_ _19432_/Q _17922_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19432_/D sky130_fd_sc_hd__mux2_1
X_17461_ _17461_/A _17461_/B vssd1 vssd1 vccd1 vccd1 _17461_/X sky130_fd_sc_hd__or2_4
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11885_ _12039_/A1 _10558_/B split7/X vssd1 vssd1 vccd1 vccd1 _11885_/X sky130_fd_sc_hd__a21o_4
XFILLER_45_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19200_ _19560_/CLK _19200_/D vssd1 vssd1 vccd1 vccd1 _19200_/Q sky130_fd_sc_hd__dfxtp_1
X_16412_ _19750_/Q _16412_/B vssd1 vssd1 vccd1 vccd1 _16418_/C sky130_fd_sc_hd__and2_2
X_13624_ _13626_/A1 _13412_/B _15762_/A _13624_/B2 vssd1 vssd1 vccd1 vccd1 _13624_/X
+ sky130_fd_sc_hd__a22o_2
X_10836_ _20402_/Q _11161_/S _10822_/X _12324_/S vssd1 vssd1 vccd1 vccd1 _10836_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17392_ _20244_/Q _17337_/B _17530_/A2 _20293_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17392_/X sky130_fd_sc_hd__a221o_1
XFILLER_73_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19131_ _19232_/CLK _19131_/D vssd1 vssd1 vccd1 vccd1 _19131_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16343_ _19724_/Q _16346_/C _18863_/A vssd1 vssd1 vccd1 vccd1 _16343_/Y sky130_fd_sc_hd__a21oi_1
X_13555_ _13624_/B2 _13542_/X _13554_/Y _19661_/D vssd1 vssd1 vccd1 vccd1 _13555_/X
+ sky130_fd_sc_hd__a22o_4
X_10767_ _12411_/A _19903_/Q _12272_/B2 _20028_/Q vssd1 vssd1 vccd1 vccd1 _10767_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ _12513_/C _12513_/D _12511_/B _12506_/D vssd1 vssd1 vccd1 vccd1 _12585_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19062_ _20407_/Q vssd1 vssd1 vccd1 vccd1 _20407_/D sky130_fd_sc_hd__clkbuf_2
X_16274_ _19690_/Q _17705_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19690_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13486_ _20916_/Q _13602_/A1 _18760_/B vssd1 vssd1 vccd1 vccd1 _13486_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ _20468_/Q _20308_/Q _12268_/S vssd1 vssd1 vccd1 vccd1 _10698_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15225_ _10933_/Y _11320_/B _15500_/A0 _14878_/B vssd1 vssd1 vccd1 vccd1 _15226_/B
+ sky130_fd_sc_hd__a31o_1
X_18013_ _20743_/Q _18013_/B vssd1 vssd1 vccd1 vccd1 _18019_/C sky130_fd_sc_hd__and2_2
X_12437_ _12437_/A _16026_/S vssd1 vssd1 vccd1 vccd1 _13178_/A sky130_fd_sc_hd__nor2_8
Xoutput407 _13800_/X vssd1 vssd1 vccd1 vccd1 din0[9] sky130_fd_sc_hd__buf_4
XFILLER_172_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15156_ _14887_/X _15155_/X _15357_/S vssd1 vssd1 vccd1 vccd1 _15157_/A sky130_fd_sc_hd__mux2_2
X_12368_ _19895_/Q _19796_/Q _12368_/S vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__mux2_1
Xoutput418 _19978_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[17] sky130_fd_sc_hd__buf_4
Xoutput429 _19988_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[27] sky130_fd_sc_hd__buf_4
XFILLER_271_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14107_ _14107_/A _14107_/B _14107_/C vssd1 vssd1 vccd1 vccd1 _14107_/X sky130_fd_sc_hd__or3_1
XFILLER_259_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11319_ _11319_/A _13523_/A _11779_/B vssd1 vssd1 vccd1 vccd1 _11319_/X sky130_fd_sc_hd__and3_1
XFILLER_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15087_ _20787_/Q _15016_/A _15021_/X input2/X _15086_/X vssd1 vssd1 vccd1 vccd1
+ _15087_/X sky130_fd_sc_hd__a221o_2
X_19964_ _20268_/CLK _19964_/D vssd1 vssd1 vccd1 vccd1 _19964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12299_ _20149_/Q _20117_/Q _12300_/S vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14038_ _14041_/A1 _14038_/A2 _10287_/X _14038_/B1 _19861_/Q vssd1 vssd1 vccd1 vccd1
+ _14105_/C sky130_fd_sc_hd__o32a_1
X_18915_ _18651_/Y _18970_/A2 _18914_/X _18901_/S vssd1 vssd1 vccd1 vccd1 _18915_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19895_ _20719_/CLK _19895_/D vssd1 vssd1 vccd1 vccd1 _19895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18846_ _18612_/Y _18867_/A2 _18844_/Y _18845_/Y vssd1 vssd1 vccd1 vccd1 _18846_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_268_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18777_ _18775_/X _18776_/X _18808_/A vssd1 vssd1 vccd1 vccd1 _20981_/D sky130_fd_sc_hd__a21oi_1
XFILLER_209_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15989_ _19731_/Q _15989_/A2 _15989_/B1 _19763_/Q vssd1 vssd1 vccd1 vccd1 _15989_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17728_ _20509_/Q _17902_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20509_/D sky130_fd_sc_hd__mux2_1
XFILLER_282_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17659_ _20445_/Q _17693_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20445_/D sky130_fd_sc_hd__mux2_1
XFILLER_211_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20670_ _20670_/CLK _20670_/D vssd1 vssd1 vccd1 vccd1 _20670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19329_ _19956_/CLK _19329_/D vssd1 vssd1 vccd1 vccd1 _19329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout601 _14650_/S vssd1 vssd1 vccd1 vccd1 _14667_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_99_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout612 _14531_/X vssd1 vssd1 vccd1 vccd1 _14558_/S sky130_fd_sc_hd__buf_6
X_20104_ _20715_/CLK _20104_/D vssd1 vssd1 vccd1 vccd1 _20104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09915_ _19387_/Q _12009_/A2 _09913_/X _12183_/C1 _09914_/X vssd1 vssd1 vccd1 vccd1
+ _09915_/X sky130_fd_sc_hd__o221a_1
XFILLER_104_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout623 _13903_/Y vssd1 vssd1 vccd1 vccd1 _13946_/B1 sky130_fd_sc_hd__buf_6
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout634 _16707_/X vssd1 vssd1 vccd1 vccd1 _16822_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_99_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout645 _16133_/X vssd1 vssd1 vccd1 vccd1 _16170_/S sky130_fd_sc_hd__buf_8
Xfanout656 _15591_/A vssd1 vssd1 vccd1 vccd1 _15402_/A sky130_fd_sc_hd__buf_4
XFILLER_113_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout667 _14108_/A2 vssd1 vssd1 vccd1 vccd1 _14106_/A2 sky130_fd_sc_hd__buf_2
X_20035_ _20694_/CLK _20035_/D vssd1 vssd1 vccd1 vccd1 _20035_/Q sky130_fd_sc_hd__dfxtp_1
X_09846_ _12828_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_258_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout678 _13862_/X vssd1 vssd1 vccd1 vccd1 _14738_/B sky130_fd_sc_hd__buf_6
XFILLER_101_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout689 _13862_/X vssd1 vssd1 vccd1 vccd1 _14031_/A2 sky130_fd_sc_hd__buf_4
XFILLER_218_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _12850_/A1 _09776_/X _11872_/A vssd1 vssd1 vccd1 vccd1 _09777_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_73_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20937_ _21004_/CLK _20937_/D vssd1 vssd1 vccd1 vccd1 _20937_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11670_ _11668_/X _11669_/X _11670_/S vssd1 vssd1 vccd1 vccd1 _11670_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ _21030_/CLK _20868_/D vssd1 vssd1 vccd1 vccd1 _20868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ _19671_/Q _20159_/Q _10621_/S vssd1 vssd1 vccd1 vccd1 _10621_/X sky130_fd_sc_hd__mux2_1
X_20799_ _20856_/CLK _20799_/D vssd1 vssd1 vccd1 vccd1 _20799_/Q sky130_fd_sc_hd__dfxtp_1
X_13340_ _13340_/A _13340_/B vssd1 vssd1 vccd1 vccd1 _13340_/Y sky130_fd_sc_hd__nand2_1
X_10552_ _19576_/Q _10551_/X _11243_/S vssd1 vssd1 vccd1 vccd1 _10553_/D sky130_fd_sc_hd__mux2_4
XFILLER_195_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13271_ _13270_/A _13270_/B _13270_/C vssd1 vssd1 vccd1 vccd1 _13271_/Y sky130_fd_sc_hd__a21oi_1
X_10483_ _20375_/Q _20439_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _10483_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_129_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21019_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15010_ _15022_/A _15022_/B _15022_/C vssd1 vssd1 vccd1 vccd1 _15021_/C sky130_fd_sc_hd__nor3_4
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12222_ _19691_/Q _20179_/Q _12368_/S vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _12153_/A1 _12152_/X _12153_/B1 vssd1 vssd1 vccd1 vccd1 _12153_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11104_ _12411_/A _19899_/Q _12272_/B2 _20024_/Q vssd1 vssd1 vccd1 vccd1 _11104_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16961_ _16958_/Y _16960_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16961_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12084_ _12084_/A _20683_/Q _12084_/C vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__or3_1
XFILLER_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18700_ _18700_/A _18700_/B vssd1 vssd1 vccd1 vccd1 _20950_/D sky130_fd_sc_hd__and2_1
XFILLER_238_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11035_ _19868_/Q _19769_/Q _11035_/S vssd1 vssd1 vccd1 vccd1 _11035_/X sky130_fd_sc_hd__mux2_1
X_15912_ _20972_/Q _15939_/A2 _15996_/B1 _20844_/Q _15911_/X vssd1 vssd1 vccd1 vccd1
+ _15912_/X sky130_fd_sc_hd__a221o_1
X_19680_ _20715_/CLK _19680_/D vssd1 vssd1 vccd1 vccd1 _19680_/Q sky130_fd_sc_hd__dfxtp_1
X_16892_ _16932_/A1 _16891_/X _16932_/B1 vssd1 vssd1 vccd1 vccd1 _16892_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18631_ _20931_/Q _18686_/B vssd1 vssd1 vccd1 vccd1 _18631_/Y sky130_fd_sc_hd__nand2_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _15843_/A _15925_/B vssd1 vssd1 vccd1 vccd1 _15843_/Y sky130_fd_sc_hd__nand2_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ _18980_/A _18562_/B vssd1 vssd1 vccd1 vccd1 _20913_/D sky130_fd_sc_hd__nor2_1
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _19223_/Q _19222_/Q _19221_/Q _13545_/B vssd1 vssd1 vccd1 vccd1 _13587_/B
+ sky130_fd_sc_hd__and4_4
X_15774_ _20903_/Q _16043_/A2 _16043_/B1 _15773_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _15774_/X sky130_fd_sc_hd__a221o_1
XFILLER_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17513_ _17525_/A1 _17512_/Y _17430_/A vssd1 vssd1 vccd1 vccd1 _20291_/D sky130_fd_sc_hd__a21oi_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14725_ _19482_/Q _17940_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19482_/D sky130_fd_sc_hd__mux2_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18493_ _18604_/B _18493_/B vssd1 vssd1 vccd1 vccd1 _18493_/X sky130_fd_sc_hd__or2_2
X_11937_ _11948_/A1 _11936_/X _11935_/X vssd1 vssd1 vccd1 vccd1 _11937_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_550 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_561 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_572 _19841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17444_ _17402_/A _17442_/A _17434_/A _17443_/X vssd1 vssd1 vccd1 vccd1 _20262_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_583 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14656_ _19418_/Q _17800_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19418_/D sky130_fd_sc_hd__mux2_1
X_11868_ _20325_/Q _11616_/B _11867_/X vssd1 vssd1 vccd1 vccd1 _11868_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_594 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10819_ _19403_/Q _12300_/S _10818_/X _09695_/A vssd1 vssd1 vccd1 vccd1 _10819_/X
+ sky130_fd_sc_hd__o211a_1
X_13607_ _20956_/Q _13607_/B vssd1 vssd1 vccd1 vccd1 _13607_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17375_ _20236_/Q _17381_/A2 _17374_/X _14482_/A vssd1 vssd1 vccd1 vccd1 _20236_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11799_ _09783_/A _11799_/B vssd1 vssd1 vccd1 vccd1 _11799_/Y sky130_fd_sc_hd__nand2b_1
X_14587_ _19353_/Q _17939_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19353_/D sky130_fd_sc_hd__mux2_1
X_19114_ _20721_/CLK _19114_/D vssd1 vssd1 vccd1 vccd1 _19114_/Q sky130_fd_sc_hd__dfxtp_4
X_16326_ _16330_/C _16326_/B vssd1 vssd1 vccd1 vccd1 _19717_/D sky130_fd_sc_hd__nor2_1
X_13538_ _15264_/A _13538_/B vssd1 vssd1 vccd1 vccd1 _13539_/B sky130_fd_sc_hd__xnor2_4
XFILLER_158_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19045_ _21041_/Q _19015_/B _19044_/X _18754_/A vssd1 vssd1 vccd1 vccd1 _21041_/D
+ sky130_fd_sc_hd__o211a_1
X_13469_ _13790_/A _13473_/B split2/A vssd1 vssd1 vccd1 vccd1 _13469_/Y sky130_fd_sc_hd__a21oi_4
X_16257_ _19673_/Q _17931_/A1 _16275_/S vssd1 vssd1 vccd1 vccd1 _19673_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15208_ _15208_/A _15208_/B _15208_/C vssd1 vssd1 vccd1 vccd1 _15208_/X sky130_fd_sc_hd__and3_1
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16188_ _19618_/Q _15943_/X _16190_/S vssd1 vssd1 vccd1 vccd1 _16189_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15139_ _20852_/Q _15322_/B _15137_/X _15138_/Y vssd1 vssd1 vccd1 vccd1 _15139_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19947_ _20081_/CLK _19947_/D vssd1 vssd1 vccd1 vccd1 _19947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _19888_/Q _19789_/Q _11889_/S vssd1 vssd1 vccd1 vccd1 _09700_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19878_ _20570_/CLK _19878_/D vssd1 vssd1 vccd1 vccd1 _19878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09631_ _09630_/X _09632_/B vssd1 vssd1 vccd1 vccd1 _09631_/X sky130_fd_sc_hd__and2b_4
XFILLER_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18829_ _19094_/Q _12589_/B _12592_/C _15442_/B vssd1 vssd1 vccd1 vccd1 _18830_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_283_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ _12513_/A _12513_/B _12588_/A _09560_/X _14894_/A vssd1 vssd1 vccd1 vccd1
+ _09562_/X sky130_fd_sc_hd__o32a_2
XFILLER_283_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09493_ _19122_/Q vssd1 vssd1 vccd1 vccd1 _09493_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20722_ _20794_/CLK _20722_/D vssd1 vssd1 vccd1 vccd1 _20722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20653_ _20685_/CLK _20653_/D vssd1 vssd1 vccd1 vccd1 _20653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20584_ _20716_/CLK _20584_/D vssd1 vssd1 vccd1 vccd1 _20584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1407 fanout1430/X vssd1 vssd1 vccd1 vccd1 _10345_/S sky130_fd_sc_hd__buf_4
Xfanout1418 fanout1422/X vssd1 vssd1 vccd1 vccd1 _11126_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_266_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1429 fanout1430/X vssd1 vssd1 vccd1 vccd1 _12248_/B1 sky130_fd_sc_hd__buf_4
XFILLER_24_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20018_ _20862_/CLK _20018_/D vssd1 vssd1 vccd1 vccd1 _20018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09829_ _09829_/A _19324_/Q _12084_/C vssd1 vssd1 vccd1 vccd1 _09829_/X sky130_fd_sc_hd__or3_1
Xfanout497 _17851_/X vssd1 vssd1 vccd1 vccd1 _17878_/S sky130_fd_sc_hd__buf_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12840_ _12839_/A _12839_/B _12839_/C _12839_/D vssd1 vssd1 vccd1 vccd1 _12842_/D
+ sky130_fd_sc_hd__o22ai_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12759_/X _12771_/B _12771_/C _12771_/D vssd1 vssd1 vccd1 vccd1 _12791_/C
+ sky130_fd_sc_hd__nand4b_2
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14510_ _19288_/Q _17835_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19288_/D sky130_fd_sc_hd__mux2_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _09839_/A _11711_/X _11715_/X _11721_/X vssd1 vssd1 vccd1 vccd1 _11723_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15442_/A _13459_/Y _15472_/Y _15489_/X vssd1 vssd1 vccd1 vccd1 _15490_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_199_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14441_ _17402_/A _17335_/B vssd1 vssd1 vccd1 vccd1 _17337_/A sky130_fd_sc_hd__nand2_4
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11653_ _20351_/Q _12043_/B vssd1 vssd1 vccd1 vccd1 _11653_/X sky130_fd_sc_hd__or2_1
XFILLER_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ _19938_/Q _10405_/C _11693_/B _12091_/S vssd1 vssd1 vccd1 vccd1 _10604_/X
+ sky130_fd_sc_hd__o31a_1
X_17160_ _20126_/Q _17788_/A1 _17166_/S vssd1 vssd1 vccd1 vccd1 _20126_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14372_ _19519_/Q _14373_/B vssd1 vssd1 vccd1 vccd1 _14372_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ _20352_/Q _11897_/B vssd1 vssd1 vccd1 vccd1 _11584_/X sky130_fd_sc_hd__or2_1
XFILLER_7_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16111_ _19580_/Q _16127_/A2 _16131_/B1 vssd1 vssd1 vccd1 vccd1 _16111_/X sky130_fd_sc_hd__o21a_1
XFILLER_155_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ _13296_/B _13323_/B _13323_/C vssd1 vssd1 vccd1 vccd1 _13323_/X sky130_fd_sc_hd__and3b_1
X_10535_ _10533_/X _10534_/X _11033_/S vssd1 vssd1 vccd1 vccd1 _10535_/X sky130_fd_sc_hd__mux2_1
X_17091_ _20061_/Q _17859_/A1 _17114_/S vssd1 vssd1 vccd1 vccd1 _20061_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13254_ _13253_/A _13253_/C _13253_/B vssd1 vssd1 vccd1 vccd1 _13254_/Y sky130_fd_sc_hd__a21oi_1
X_16042_ _20881_/Q _16042_/A2 fanout819/X vssd1 vssd1 vccd1 vccd1 _16042_/X sky130_fd_sc_hd__o21ba_1
XFILLER_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10466_ _10032_/Y _10465_/Y _09638_/Y vssd1 vssd1 vccd1 vccd1 _10466_/X sky130_fd_sc_hd__a21o_1
XFILLER_182_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12205_ _12206_/B _12206_/C _13432_/A vssd1 vssd1 vccd1 vccd1 _12288_/C sky130_fd_sc_hd__o21ai_2
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _13653_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13631_/B sky130_fd_sc_hd__nand2_8
XFILLER_135_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10397_ _19409_/Q _20568_/Q _10397_/S vssd1 vssd1 vccd1 vccd1 _10397_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_wb_clk_i ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_269_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19801_ _20660_/CLK _19801_/D vssd1 vssd1 vccd1 vccd1 _19801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12136_ _12135_/A _12122_/Y _12136_/B1 vssd1 vssd1 vccd1 vccd1 _12136_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_285_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17993_ _20735_/Q _17989_/B _17992_/Y vssd1 vssd1 vccd1 vccd1 _20735_/D sky130_fd_sc_hd__o21a_1
XFILLER_2_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19732_ _20816_/CLK _19732_/D vssd1 vssd1 vccd1 vccd1 _19732_/Q sky130_fd_sc_hd__dfxtp_1
X_16944_ _19984_/Q _16876_/A _16943_/Y _17012_/C1 vssd1 vssd1 vccd1 vccd1 _19984_/D
+ sky130_fd_sc_hd__a211o_1
Xfanout1930 _18476_/A vssd1 vssd1 vccd1 vccd1 _18710_/A sky130_fd_sc_hd__buf_4
X_12067_ _19824_/Q _19328_/Q _12070_/S vssd1 vssd1 vccd1 vccd1 _12067_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_97_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20727_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1941 _13890_/C1 vssd1 vssd1 vccd1 vccd1 _16131_/B1 sky130_fd_sc_hd__buf_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1952 fanout1960/X vssd1 vssd1 vccd1 vccd1 _16381_/B1 sky130_fd_sc_hd__buf_2
XFILLER_277_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1963 _18960_/A vssd1 vssd1 vccd1 vccd1 _18973_/A sky130_fd_sc_hd__buf_2
X_11018_ _15545_/A vssd1 vssd1 vccd1 vccd1 _11018_/Y sky130_fd_sc_hd__inv_2
X_19663_ _20561_/CLK _19663_/D vssd1 vssd1 vccd1 vccd1 _19663_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1974 _13595_/A vssd1 vssd1 vccd1 vccd1 _18877_/A sky130_fd_sc_hd__buf_4
XFILLER_237_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1985 _16896_/C1 vssd1 vssd1 vccd1 vccd1 _16451_/A sky130_fd_sc_hd__buf_4
X_16875_ _17008_/B1 _16872_/X _16874_/X _16875_/B2 vssd1 vssd1 vccd1 vccd1 _16876_/B
+ sky130_fd_sc_hd__o2bb2a_4
Xclkbuf_leaf_26_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20635_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1996 fanout2002/X vssd1 vssd1 vccd1 vccd1 _18704_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18614_ _18856_/A _18614_/B vssd1 vssd1 vccd1 vccd1 _20926_/D sky130_fd_sc_hd__nor2_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _20873_/Q _16018_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15826_/X sky130_fd_sc_hd__o21ba_1
X_19594_ _19621_/CLK _19594_/D vssd1 vssd1 vccd1 vccd1 _19594_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18545_ _20908_/Q fanout750/X _18544_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18546_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_234_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15757_ _15526_/B _15740_/Y _15756_/X _15526_/Y vssd1 vssd1 vccd1 vccd1 _15757_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12969_ _19115_/Q _19098_/Q _19096_/Q vssd1 vssd1 vccd1 vccd1 _12972_/C sky130_fd_sc_hd__or3_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14708_ _19465_/Q _17189_/A1 _14719_/S vssd1 vssd1 vccd1 vccd1 _19465_/D sky130_fd_sc_hd__mux2_1
XFILLER_261_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18476_ _18476_/A _18476_/B vssd1 vssd1 vccd1 vccd1 _20885_/D sky130_fd_sc_hd__and2_1
X_15688_ _19720_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15688_/X sky130_fd_sc_hd__or2_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_380 _15649_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_391 _16869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17427_ _20258_/Q _20251_/Q _17433_/S vssd1 vssd1 vccd1 vccd1 _17428_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14639_ _19401_/Q _17923_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19401_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17358_ _20227_/Q _17364_/A2 _17362_/B1 _20276_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17358_/X sky130_fd_sc_hd__a221o_1
XFILLER_193_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16309_ _19711_/Q _16308_/B _18414_/A vssd1 vssd1 vccd1 vccd1 _16310_/B sky130_fd_sc_hd__o21ai_1
X_17289_ _20202_/Q _17331_/A2 _17287_/X _17288_/X _17331_/C1 vssd1 vssd1 vccd1 vccd1
+ _20202_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19028_ _18265_/Y _19046_/A2 _19048_/B1 _12551_/A _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19028_/X sky130_fd_sc_hd__a221o_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09614_ _12513_/D _11261_/C vssd1 vssd1 vccd1 vccd1 _09614_/X sky130_fd_sc_hd__and2_4
XFILLER_284_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ _19154_/Q _12579_/C vssd1 vssd1 vccd1 vccd1 _09556_/A sky130_fd_sc_hd__nand2_2
XFILLER_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20705_ _20710_/CLK _20705_/D vssd1 vssd1 vccd1 vccd1 _20705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20636_ _20683_/CLK _20636_/D vssd1 vssd1 vccd1 vccd1 _20636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20567_ _20701_/CLK _20567_/D vssd1 vssd1 vccd1 vccd1 _20567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _19637_/Q _19943_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20498_ _20662_/CLK _20498_/D vssd1 vssd1 vccd1 vccd1 _20498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10251_ _10247_/X _10250_/X _11375_/S vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10182_ _11391_/A _19910_/Q _12346_/S _20035_/Q vssd1 vssd1 vccd1 vccd1 _10182_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1204 _17331_/A2 vssd1 vssd1 vccd1 vccd1 _17280_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_278_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1215 _14807_/X vssd1 vssd1 vccd1 vccd1 _16133_/C sky130_fd_sc_hd__buf_8
Xfanout1226 _15527_/A vssd1 vssd1 vccd1 vccd1 _12486_/B sky130_fd_sc_hd__clkbuf_8
Xfanout1237 _09683_/X vssd1 vssd1 vccd1 vccd1 _10037_/B sky130_fd_sc_hd__buf_6
X_14990_ _15308_/B _14997_/C vssd1 vssd1 vccd1 vccd1 _14993_/S sky130_fd_sc_hd__nand2_1
XFILLER_120_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1248 _17370_/C1 vssd1 vssd1 vccd1 vccd1 _17362_/C1 sky130_fd_sc_hd__buf_6
XFILLER_259_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1259 _12730_/A2 vssd1 vssd1 vccd1 vccd1 _12847_/A2 sky130_fd_sc_hd__buf_8
XFILLER_247_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13941_ _13941_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _13941_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16660_ _19917_/Q _17872_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19917_/D sky130_fd_sc_hd__mux2_1
XFILLER_235_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13872_ _19090_/Q _14527_/A2 _13896_/B1 _19156_/Q _16193_/A vssd1 vssd1 vccd1 vccd1
+ _19090_/D sky130_fd_sc_hd__o221a_1
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15611_ _15352_/X _15356_/Y _15611_/S vssd1 vssd1 vccd1 vccd1 _15611_/X sky130_fd_sc_hd__mux2_1
XFILLER_216_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12823_ _15713_/A _15526_/A vssd1 vssd1 vccd1 vccd1 _12823_/Y sky130_fd_sc_hd__nand2_1
XFILLER_250_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16591_ _16591_/A _16591_/B vssd1 vssd1 vccd1 vccd1 _19861_/D sky130_fd_sc_hd__or2_1
XFILLER_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18330_ _20820_/Q _18341_/B _18329_/Y _18396_/A vssd1 vssd1 vccd1 vccd1 _20820_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15542_ _15644_/A1 _16851_/B _15528_/Y vssd1 vssd1 vccd1 vccd1 _15542_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12754_/A _12754_/B vssd1 vssd1 vccd1 vccd1 _12754_/X sky130_fd_sc_hd__or2_1
XFILLER_215_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _20806_/Q _18260_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18262_/B sky130_fd_sc_hd__mux2_1
XFILLER_98_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11705_ _12105_/A _12091_/S _11704_/X _10409_/A vssd1 vssd1 vccd1 vccd1 _11705_/X
+ sky130_fd_sc_hd__a31o_1
X_12685_ _12686_/B _12686_/C _12686_/A vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__a21oi_4
XFILLER_15_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15473_ _15473_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _15473_/Y sky130_fd_sc_hd__nand2_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_144_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19695_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17212_ _20176_/Q _17946_/A1 _17212_/S vssd1 vssd1 vccd1 vccd1 _20176_/D sky130_fd_sc_hd__mux2_1
X_14424_ _14424_/A _14424_/B vssd1 vssd1 vccd1 vccd1 _14426_/D sky130_fd_sc_hd__nor2_1
X_11636_ _09752_/A _19353_/Q _20708_/Q _12013_/S vssd1 vssd1 vccd1 vccd1 _11636_/X
+ sky130_fd_sc_hd__a22o_1
X_18192_ _18418_/A _18192_/B vssd1 vssd1 vccd1 vccd1 _20792_/D sky130_fd_sc_hd__and2_1
XFILLER_187_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17143_ _20111_/Q _17805_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20111_/D sky130_fd_sc_hd__mux2_1
X_14355_ _14354_/A _14354_/B _14354_/C vssd1 vssd1 vccd1 vccd1 _14361_/B sky130_fd_sc_hd__a21oi_1
X_11567_ _12192_/A1 _11556_/X _11560_/X _11566_/X vssd1 vssd1 vccd1 vccd1 _11568_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10518_ _19875_/Q _19776_/Q _10518_/S vssd1 vssd1 vccd1 vccd1 _10518_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13306_ _13355_/B _13303_/X _13304_/Y _13305_/Y _18671_/B vssd1 vssd1 vccd1 vccd1
+ _13306_/X sky130_fd_sc_hd__o311a_1
XFILLER_157_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17074_ _20046_/Q _17910_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20046_/D sky130_fd_sc_hd__mux2_1
X_14286_ _14397_/A _14397_/B _14286_/C vssd1 vssd1 vccd1 vccd1 _14286_/X sky130_fd_sc_hd__or3_1
XFILLER_171_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ _20349_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _11498_/X sky130_fd_sc_hd__or2_1
X_13237_ _13015_/X _13016_/Y _13084_/Y _13397_/B _13236_/Y vssd1 vssd1 vccd1 vccd1
+ _13237_/Y sky130_fd_sc_hd__a311oi_4
X_16025_ _16053_/A _16025_/B vssd1 vssd1 vccd1 vccd1 _16025_/Y sky130_fd_sc_hd__nor2_1
X_10449_ _13670_/A1 split4/A _10448_/X _12075_/C1 vssd1 vssd1 vccd1 vccd1 _13680_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_226_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ _13167_/A _11743_/B _13167_/B _11741_/A vssd1 vssd1 vccd1 vccd1 _13415_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_151_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12119_ _12035_/A _12033_/Y _12118_/X vssd1 vssd1 vccd1 vccd1 _12202_/B sky130_fd_sc_hd__o21a_1
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17976_ _20730_/Q _20729_/Q _17976_/C vssd1 vssd1 vccd1 vccd1 _17982_/C sky130_fd_sc_hd__and3_1
X_13099_ _09488_/A _19246_/Q _14802_/C1 vssd1 vssd1 vccd1 vccd1 _13100_/B sky130_fd_sc_hd__o21a_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19715_ _20863_/CLK _19715_/D vssd1 vssd1 vccd1 vccd1 _19715_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_242_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16927_ _16924_/Y _16926_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16927_/Y sky130_fd_sc_hd__a21oi_4
Xfanout1760 _09488_/Y vssd1 vssd1 vccd1 vccd1 _13139_/A sky130_fd_sc_hd__buf_6
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1771 _14244_/A1 vssd1 vssd1 vccd1 vccd1 _14275_/A1 sky130_fd_sc_hd__buf_4
Xfanout1782 _20255_/Q vssd1 vssd1 vccd1 vccd1 _17460_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_238_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1793 _18149_/S vssd1 vssd1 vccd1 vccd1 _14917_/A sky130_fd_sc_hd__buf_2
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19646_ _20077_/CLK _19646_/D vssd1 vssd1 vccd1 vccd1 _19646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16858_ _16887_/A _16858_/B vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15809_ _16002_/A1 _15795_/Y _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15809_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19577_ _19577_/CLK _19577_/D vssd1 vssd1 vccd1 vccd1 _19577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16789_ input103/X input74/X _16799_/S vssd1 vssd1 vccd1 vccd1 _16790_/A sky130_fd_sc_hd__mux2_2
XFILLER_281_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18528_ _18960_/A _18528_/B vssd1 vssd1 vccd1 vccd1 _20902_/D sky130_fd_sc_hd__nor2_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18459_ _18570_/B _18459_/B vssd1 vssd1 vccd1 vccd1 _18459_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20421_ _20421_/CLK _20421_/D vssd1 vssd1 vccd1 vccd1 _20421_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20352_ _20676_/CLK _20352_/D vssd1 vssd1 vccd1 vccd1 _20352_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20283_ _21030_/CLK _20283_/D vssd1 vssd1 vccd1 vccd1 _20283_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09528_ input49/X vssd1 vssd1 vccd1 vccd1 _09528_/Y sky130_fd_sc_hd__inv_2
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12470_ _16054_/B _12471_/B vssd1 vssd1 vccd1 vccd1 _12470_/Y sky130_fd_sc_hd__nor2_4
XFILLER_177_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _12138_/A1 _19479_/Q _19447_/Q _12124_/S _11423_/C1 vssd1 vssd1 vccd1 vccd1
+ _11421_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20619_ _20655_/CLK _20619_/D vssd1 vssd1 vccd1 vccd1 _20619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14140_ _14138_/Y _14140_/B vssd1 vssd1 vccd1 vccd1 _14141_/B sky130_fd_sc_hd__and2b_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11352_ _20633_/Q _20597_/Q _11358_/S vssd1 vssd1 vccd1 vccd1 _11352_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10303_ _20132_/Q _20100_/Q _10303_/S vssd1 vssd1 vccd1 vccd1 _10303_/X sky130_fd_sc_hd__mux2_1
X_14071_ _14099_/A _14099_/B _14071_/C vssd1 vssd1 vccd1 vccd1 _14071_/X sky130_fd_sc_hd__or3_1
XFILLER_152_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11283_ _11280_/Y _11281_/Y _11313_/B vssd1 vssd1 vccd1 vccd1 _15035_/S sky130_fd_sc_hd__a21o_4
X_13022_ _20968_/Q _20902_/Q vssd1 vssd1 vccd1 vccd1 _13394_/B sky130_fd_sc_hd__nand2_2
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10234_ _19813_/Q _19317_/Q _10986_/B vssd1 vssd1 vccd1 vccd1 _10234_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1001 _14904_/X vssd1 vssd1 vccd1 vccd1 _16000_/A1 sky130_fd_sc_hd__buf_8
XFILLER_3_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17830_ _20605_/Q _17902_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20605_/D sky130_fd_sc_hd__mux2_1
Xfanout1012 _16028_/C vssd1 vssd1 vccd1 vccd1 _15981_/B sky130_fd_sc_hd__buf_4
XFILLER_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10165_ _12464_/A _11726_/S _10164_/Y vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__o21a_2
Xfanout1023 _16963_/B1 vssd1 vssd1 vccd1 vccd1 _17004_/B1 sky130_fd_sc_hd__buf_6
Xfanout1034 _14901_/Y vssd1 vssd1 vccd1 vccd1 _16878_/A sky130_fd_sc_hd__buf_6
XFILLER_79_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1045 _16608_/A1 vssd1 vssd1 vccd1 vccd1 _17888_/A1 sky130_fd_sc_hd__buf_2
XFILLER_255_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1056 _10894_/X vssd1 vssd1 vccd1 vccd1 _17924_/A1 sky130_fd_sc_hd__clkbuf_2
X_17761_ _20540_/Q _17901_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20540_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14973_ _14973_/A _14973_/B _14973_/C vssd1 vssd1 vccd1 vccd1 _14981_/B sky130_fd_sc_hd__or3_1
Xfanout1067 _09749_/X vssd1 vssd1 vccd1 vccd1 _11397_/B2 sky130_fd_sc_hd__buf_6
X_10096_ _12084_/A _20505_/Q _10092_/S _20537_/Q vssd1 vssd1 vccd1 vccd1 _10096_/X
+ sky130_fd_sc_hd__o22a_1
Xfanout1078 _13193_/Y vssd1 vssd1 vccd1 vccd1 _18949_/B1 sky130_fd_sc_hd__buf_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1089 _17917_/A1 vssd1 vssd1 vccd1 vccd1 _17674_/A1 sky130_fd_sc_hd__buf_4
X_19500_ _21021_/CLK _19500_/D vssd1 vssd1 vccd1 vccd1 _19500_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16712_ _20621_/Q _16945_/B vssd1 vssd1 vccd1 vccd1 _17219_/B sky130_fd_sc_hd__and2_4
XFILLER_48_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13924_ _19128_/Q _13921_/B _13932_/B1 _13458_/Y vssd1 vssd1 vccd1 vccd1 _19128_/D
+ sky130_fd_sc_hd__o22a_1
X_17692_ _20476_/Q _17692_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20476_/D sky130_fd_sc_hd__mux2_1
XFILLER_247_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19431_ _20561_/CLK _19431_/D vssd1 vssd1 vccd1 vccd1 _19431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16643_ _19900_/Q _17855_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19900_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13855_ _19659_/Q _16232_/B _13854_/Y vssd1 vssd1 vccd1 vccd1 _13855_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_263_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19362_ _20585_/CLK _19362_/D vssd1 vssd1 vccd1 vccd1 _19362_/Q sky130_fd_sc_hd__dfxtp_1
X_12806_ _19516_/Q _12916_/A2 _12805_/X _12916_/B2 vssd1 vssd1 vccd1 vccd1 _12808_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_90_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16574_ _19853_/Q _16578_/A2 _16578_/B1 input24/X vssd1 vssd1 vccd1 vccd1 _16575_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10998_ _20336_/Q _09623_/B _11169_/B _11170_/B1 vssd1 vssd1 vccd1 vccd1 _10998_/X
+ sky130_fd_sc_hd__o31a_1
X_13786_ _13612_/A split3/A _13568_/Y _13566_/Y _13244_/X vssd1 vssd1 vccd1 vccd1
+ _13786_/X sky130_fd_sc_hd__a32o_4
XFILLER_231_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18313_ _19558_/Q _18313_/B vssd1 vssd1 vccd1 vccd1 _18313_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_188_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _19539_/Q _15591_/A _15524_/Y _16167_/C1 vssd1 vssd1 vccd1 vccd1 _19539_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12749_/A _12749_/B vssd1 vssd1 vccd1 vccd1 _13309_/A sky130_fd_sc_hd__nor2_1
X_19293_ _20647_/CLK _19293_/D vssd1 vssd1 vccd1 vccd1 _19293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18248_/B _14294_/B _18243_/Y vssd1 vssd1 vccd1 vccd1 _18517_/B sky130_fd_sc_hd__o21ai_4
XFILLER_188_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15456_ _15644_/A1 _16824_/B _15443_/Y vssd1 vssd1 vccd1 vccd1 _15456_/X sky130_fd_sc_hd__o21a_1
X_12668_ _12668_/A _12738_/B vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__or2_1
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14407_ _14427_/A _14405_/X _14406_/X _13139_/A vssd1 vssd1 vccd1 vccd1 _14407_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18175_ _18471_/B vssd1 vssd1 vccd1 vccd1 _18175_/Y sky130_fd_sc_hd__inv_2
X_11619_ _20480_/Q _11641_/S _11213_/B _11617_/X _11618_/X vssd1 vssd1 vccd1 vccd1
+ _11619_/X sky130_fd_sc_hd__a311o_1
X_15387_ _20922_/Q _15567_/A2 _15386_/X vssd1 vssd1 vccd1 vccd1 _15387_/X sky130_fd_sc_hd__o21a_2
XFILLER_184_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12599_ _19500_/Q _12647_/A vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__and2_2
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17126_ _20094_/Q _17788_/A1 _17132_/S vssd1 vssd1 vccd1 vccd1 _20094_/D sky130_fd_sc_hd__mux2_1
XFILLER_274_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14338_ _14437_/A _14437_/B _14338_/C vssd1 vssd1 vccd1 vccd1 _14338_/X sky130_fd_sc_hd__or3_1
XFILLER_171_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17057_ _20029_/Q _17684_/A1 _17080_/S vssd1 vssd1 vccd1 vccd1 _20029_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14269_ _19509_/Q _14269_/B vssd1 vssd1 vccd1 vccd1 _14270_/B sky130_fd_sc_hd__nor2_1
XFILLER_98_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16008_ _19556_/Q _16007_/A _16007_/Y _16189_/A vssd1 vssd1 vccd1 vccd1 _19556_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20704_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17959_ _20724_/Q _20723_/Q _17959_/C vssd1 vssd1 vccd1 vccd1 _17961_/A sky130_fd_sc_hd__and3_1
XFILLER_239_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1590 _09623_/B vssd1 vssd1 vccd1 vccd1 _11270_/A2 sky130_fd_sc_hd__buf_6
X_20970_ _21000_/CLK _20970_/D vssd1 vssd1 vccd1 vccd1 _20970_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_226_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19629_ _20463_/CLK _19629_/D vssd1 vssd1 vccd1 vccd1 _19629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20404_ _20759_/CLK _20404_/D vssd1 vssd1 vccd1 vccd1 _20404_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_215_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20335_ _20686_/CLK _20335_/D vssd1 vssd1 vccd1 vccd1 _20335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20266_ _21015_/CLK _20266_/D vssd1 vssd1 vccd1 vccd1 _20266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput104 dout0[7] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20197_ _20688_/CLK _20197_/D vssd1 vssd1 vccd1 vccd1 _20197_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput115 dout1[17] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput126 dout1[27] vssd1 vssd1 vccd1 vccd1 input126/X sky130_fd_sc_hd__clkbuf_2
XFILLER_277_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 dout1[37] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__clkbuf_2
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput148 dout1[47] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__clkbuf_2
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput159 dout1[57] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _20145_/Q _20113_/Q _11978_/S vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10921_ _20465_/Q _09688_/B _10235_/S vssd1 vssd1 vccd1 vccd1 _10921_/X sky130_fd_sc_hd__a21o_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10852_ _12332_/A _19902_/Q _12334_/S0 _20027_/Q vssd1 vssd1 vccd1 vccd1 _10852_/X
+ sky130_fd_sc_hd__o22a_1
X_13640_ _15954_/A _13189_/B _16239_/B _13478_/B vssd1 vssd1 vccd1 vccd1 _13640_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_60_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10692_/A _19468_/Q _19436_/Q _11116_/S _12419_/C1 vssd1 vssd1 vccd1 vccd1
+ _10783_/X sky130_fd_sc_hd__a221o_1
XFILLER_169_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13571_ _13571_/A _13571_/B vssd1 vssd1 vccd1 vccd1 _13572_/B sky130_fd_sc_hd__nor2_1
XFILLER_213_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _20920_/Q _15323_/A _15309_/X _14972_/A _15308_/X vssd1 vssd1 vccd1 vccd1
+ _15310_/X sky130_fd_sc_hd__a221o_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _20915_/Q _12982_/C vssd1 vssd1 vccd1 vccd1 _12522_/Y sky130_fd_sc_hd__nor2_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _18054_/A _16290_/B _16294_/C vssd1 vssd1 vccd1 vccd1 _19704_/D sky130_fd_sc_hd__nor3_1
XFILLER_197_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15241_ _19738_/Q _15453_/A2 _15231_/X _15021_/A _15240_/X vssd1 vssd1 vccd1 vccd1
+ _15241_/X sky130_fd_sc_hd__a221o_1
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12453_ _16028_/A _16028_/B _12451_/Y _12449_/X vssd1 vssd1 vccd1 vccd1 _12454_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_184_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11404_ _11400_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11772_/B sky130_fd_sc_hd__and2b_2
X_12384_ _12383_/A _12370_/Y _09502_/A vssd1 vssd1 vccd1 vccd1 _12384_/Y sky130_fd_sc_hd__a21oi_1
X_15172_ _15357_/S _15172_/B vssd1 vssd1 vccd1 vccd1 _15172_/X sky130_fd_sc_hd__or2_1
XFILLER_126_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11335_ _19873_/Q _19774_/Q _11342_/S vssd1 vssd1 vccd1 vccd1 _11335_/X sky130_fd_sc_hd__mux2_1
X_14123_ _19494_/Q _14123_/B vssd1 vssd1 vccd1 vccd1 _14131_/A sky130_fd_sc_hd__nand2_1
X_19980_ _20816_/CLK _19980_/D vssd1 vssd1 vccd1 vccd1 _19980_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18931_ _18538_/X _18971_/B _18929_/X _18930_/Y vssd1 vssd1 vccd1 vccd1 _18932_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_268_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14054_ _19186_/Q _14108_/A2 _14053_/X _16097_/B1 vssd1 vssd1 vccd1 vccd1 _19186_/D
+ sky130_fd_sc_hd__o211a_1
X_11266_ _11266_/A1 _20657_/Q _11270_/A2 _11256_/S vssd1 vssd1 vccd1 vccd1 _11266_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10217_ _19413_/Q _20572_/Q _10217_/S vssd1 vssd1 vccd1 vccd1 _10217_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13005_ _20976_/Q _20910_/Q vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__nand2_1
XFILLER_239_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18862_ _18508_/X _18861_/B _18860_/X _18861_/Y vssd1 vssd1 vccd1 vccd1 _18863_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_267_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11197_ _19367_/Q _12412_/A2 _11195_/X _09738_/A _11196_/X vssd1 vssd1 vccd1 vccd1
+ _11197_/X sky130_fd_sc_hd__o221a_1
XFILLER_279_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17813_ _17851_/A _17851_/B _17813_/C vssd1 vssd1 vccd1 vccd1 _17813_/X sky130_fd_sc_hd__and3_4
XFILLER_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10148_ _20638_/Q _20602_/Q _10924_/S vssd1 vssd1 vccd1 vccd1 _10148_/X sky130_fd_sc_hd__mux2_1
XFILLER_282_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18793_ _20984_/Q _18840_/B vssd1 vssd1 vccd1 vccd1 _18793_/Y sky130_fd_sc_hd__nand2_1
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17744_ _17744_/A _17850_/B vssd1 vssd1 vccd1 vccd1 _17745_/C sky130_fd_sc_hd__nor2_1
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14956_ _14957_/B vssd1 vssd1 vccd1 vccd1 _14956_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10079_ _19877_/Q _10400_/S vssd1 vssd1 vccd1 vccd1 _10079_/X sky130_fd_sc_hd__or2_1
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13907_ _13907_/A _13921_/B vssd1 vssd1 vccd1 vccd1 _13907_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17675_ _17850_/A _17675_/B vssd1 vssd1 vccd1 vccd1 _17676_/C sky130_fd_sc_hd__nor2_1
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _14885_/B _14886_/X _15170_/A vssd1 vssd1 vccd1 vccd1 _14887_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19414_ _20573_/CLK _19414_/D vssd1 vssd1 vccd1 vccd1 _19414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16626_ _19885_/Q _17940_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19885_/D sky130_fd_sc_hd__mux2_1
X_13838_ _20258_/Q _20257_/Q vssd1 vssd1 vccd1 vccd1 _13839_/D sky130_fd_sc_hd__nand2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19345_ _20711_/CLK _19345_/D vssd1 vssd1 vccd1 vccd1 _19345_/Q sky130_fd_sc_hd__dfxtp_1
X_16557_ _16557_/A _16557_/B vssd1 vssd1 vccd1 vccd1 _19844_/D sky130_fd_sc_hd__or2_1
XFILLER_241_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13769_ _13769_/A _13769_/B vssd1 vssd1 vccd1 vccd1 _13770_/B sky130_fd_sc_hd__nor2_8
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15508_ _21024_/Q _20992_/Q _15508_/S vssd1 vssd1 vccd1 vccd1 _15508_/X sky130_fd_sc_hd__mux2_1
X_19276_ _20706_/CLK _19276_/D vssd1 vssd1 vccd1 vccd1 _19276_/Q sky130_fd_sc_hd__dfxtp_1
X_16488_ _19797_/Q _17708_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19797_/D sky130_fd_sc_hd__mux2_1
X_18227_ _18418_/A _18227_/B vssd1 vssd1 vccd1 vccd1 _20799_/D sky130_fd_sc_hd__and2_1
XFILLER_176_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15439_ _10540_/X _15500_/A0 _12470_/Y _13611_/A _12579_/D vssd1 vssd1 vccd1 vccd1
+ _15439_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_191_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18158_ _11235_/A _18198_/B vssd1 vssd1 vccd1 vccd1 _18158_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_191_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17109_ _20079_/Q _17945_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20079_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18089_ _20770_/Q _18087_/B _18088_/Y vssd1 vssd1 vccd1 vccd1 _20770_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20120_ _20563_/CLK _20120_/D vssd1 vssd1 vccd1 vccd1 _20120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09931_ _19419_/Q _20578_/Q _09931_/S vssd1 vssd1 vccd1 vccd1 _09931_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout805 _17461_/X vssd1 vssd1 vccd1 vccd1 _17495_/A1 sky130_fd_sc_hd__buf_8
Xfanout816 _13740_/B vssd1 vssd1 vccd1 vccd1 _13659_/A sky130_fd_sc_hd__buf_4
X_20051_ _20662_/CLK _20051_/D vssd1 vssd1 vccd1 vccd1 _20051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _09862_/A vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__inv_2
Xfanout827 _13685_/A vssd1 vssd1 vccd1 vccd1 _13718_/A sky130_fd_sc_hd__buf_6
XFILLER_97_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout838 _18491_/B2 vssd1 vssd1 vccd1 vccd1 _18557_/B2 sky130_fd_sc_hd__buf_4
Xfanout849 _18324_/Y vssd1 vssd1 vccd1 vccd1 _18343_/B sky130_fd_sc_hd__buf_6
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _19887_/Q _19788_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _09793_/X sky130_fd_sc_hd__mux2_1
XFILLER_274_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20953_ _21019_/CLK _20953_/D vssd1 vssd1 vccd1 vccd1 _20953_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _21015_/CLK _20884_/D vssd1 vssd1 vccd1 vccd1 _20884_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11120_ _12427_/A1 _19464_/Q _19432_/Q _11126_/B _12347_/C1 vssd1 vssd1 vccd1 vccd1
+ _11120_/X sky130_fd_sc_hd__a221o_1
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20318_ _20645_/CLK _20318_/D vssd1 vssd1 vccd1 vccd1 _20318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11051_ _11054_/B vssd1 vssd1 vccd1 vccd1 _11051_/Y sky130_fd_sc_hd__inv_2
X_20249_ _20300_/CLK _20249_/D vssd1 vssd1 vccd1 vccd1 _20249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10002_ _09999_/X _10001_/X _11949_/S vssd1 vssd1 vccd1 vccd1 _10002_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _12583_/B _14809_/Y _16133_/B _16133_/A vssd1 vssd1 vccd1 vccd1 _14810_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _13414_/Y _15981_/B _15219_/Y vssd1 vssd1 vccd1 vccd1 _15790_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14741_ _19495_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14741_/X sky130_fd_sc_hd__or2_1
XFILLER_83_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _19519_/Q _15870_/A _15895_/S vssd1 vssd1 vccd1 vccd1 _12115_/B sky130_fd_sc_hd__mux2_8
XFILLER_218_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10904_ _19933_/Q _09623_/B _11169_/B _11170_/B1 vssd1 vssd1 vccd1 vccd1 _10904_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _20265_/Q _17460_/A2 _16191_/A _17459_/X vssd1 vssd1 vccd1 vccd1 _20265_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14672_ _19431_/Q _17678_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19431_/D sky130_fd_sc_hd__mux2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ _19552_/Q _12155_/A2 _12155_/B1 _19616_/Q vssd1 vssd1 vccd1 vccd1 _11884_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16411_ _18094_/A _16411_/B _16412_/B vssd1 vssd1 vccd1 vccd1 _19749_/D sky130_fd_sc_hd__nor3_1
XFILLER_72_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13623_ _13626_/A1 _13388_/C _13428_/B _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13623_/X
+ sky130_fd_sc_hd__a22o_2
X_10835_ _12324_/S _10834_/X _10833_/X _12398_/C1 vssd1 vssd1 vccd1 vccd1 _10835_/X
+ sky130_fd_sc_hd__a211o_1
X_17391_ _20244_/Q _17401_/A2 _17390_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _20244_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19130_ _20930_/CLK _19130_/D vssd1 vssd1 vccd1 vccd1 _19130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16342_ _16346_/C _16342_/B vssd1 vssd1 vccd1 vccd1 _19723_/D sky130_fd_sc_hd__nor2_1
XFILLER_198_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13554_ _16241_/A _13915_/A vssd1 vssd1 vccd1 vccd1 _13554_/Y sky130_fd_sc_hd__nor2_2
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10766_ _19500_/Q _11189_/B vssd1 vssd1 vccd1 vccd1 _10766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12505_ _12513_/A _12513_/B _12514_/C _19168_/Q vssd1 vssd1 vccd1 vccd1 _12506_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19061_ _20406_/Q vssd1 vssd1 vccd1 vccd1 _20406_/D sky130_fd_sc_hd__clkbuf_2
X_16273_ _19689_/Q _17704_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19689_/D sky130_fd_sc_hd__mux2_1
X_10697_ _20372_/Q _20436_/Q _12268_/S vssd1 vssd1 vccd1 vccd1 _10697_/X sky130_fd_sc_hd__mux2_1
X_13485_ _19217_/Q _14110_/C _13575_/C vssd1 vssd1 vccd1 vccd1 _13485_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18012_ _18096_/A _18012_/B _18013_/B vssd1 vssd1 vccd1 vccd1 _20742_/D sky130_fd_sc_hd__nor3_1
XFILLER_139_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15224_ _15610_/A1 _15223_/X _15610_/B1 vssd1 vssd1 vccd1 vccd1 _15224_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_157_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12436_ _12436_/A _12443_/B vssd1 vssd1 vccd1 vccd1 _16026_/S sky130_fd_sc_hd__and2_4
XFILLER_154_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15155_ _15051_/X _15054_/X _15155_/S vssd1 vssd1 vccd1 vccd1 _15155_/X sky130_fd_sc_hd__mux2_1
Xoutput408 _13852_/X vssd1 vssd1 vccd1 vccd1 jtag_tdo sky130_fd_sc_hd__buf_4
XFILLER_5_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput419 _19979_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[18] sky130_fd_sc_hd__buf_4
X_12367_ _10385_/A _12366_/X _12365_/X vssd1 vssd1 vccd1 vccd1 _12367_/X sky130_fd_sc_hd__a21o_2
XFILLER_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ _19212_/Q _14106_/A2 _14105_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1 _19212_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_181_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11318_ _13495_/A _11780_/B _11052_/Y vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__a21o_2
X_15086_ _20851_/Q _15085_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15086_/X sky130_fd_sc_hd__mux2_1
X_12298_ _12306_/A1 _12296_/X _12297_/X vssd1 vssd1 vccd1 vccd1 _12298_/X sky130_fd_sc_hd__o21a_1
X_19963_ _20624_/CLK _19963_/D vssd1 vssd1 vccd1 vccd1 _19963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14037_ _19179_/Q _14043_/A2 _14040_/B1 _14036_/X _14104_/C1 vssd1 vssd1 vccd1 vccd1
+ _19179_/D sky130_fd_sc_hd__o221a_1
X_11249_ _19662_/Q _20150_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _11249_/X sky130_fd_sc_hd__mux2_1
X_18914_ _09491_/Y _18913_/X _18955_/A vssd1 vssd1 vccd1 vccd1 _18914_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19894_ _20179_/CLK _19894_/D vssd1 vssd1 vccd1 vccd1 _19894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18845_ _19129_/Q _12533_/B _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18845_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18776_ _18463_/X _09478_/Y _18840_/B vssd1 vssd1 vccd1 vccd1 _18776_/X sky130_fd_sc_hd__mux2_1
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15988_ _15988_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15988_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17727_ _20508_/Q _17901_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20508_/D sky130_fd_sc_hd__mux2_1
X_14939_ _14945_/A _14983_/A vssd1 vssd1 vccd1 vccd1 _14939_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17658_ _20444_/Q _17935_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20444_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16609_ _19868_/Q _17189_/A1 _16620_/S vssd1 vssd1 vccd1 vccd1 _19868_/D sky130_fd_sc_hd__mux2_1
XFILLER_211_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17589_ _20347_/Q _17866_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20347_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19328_ _20683_/CLK _19328_/D vssd1 vssd1 vccd1 vccd1 _19328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19259_ _21016_/CLK _19259_/D vssd1 vssd1 vccd1 vccd1 _19259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20103_ _20641_/CLK _20103_/D vssd1 vssd1 vccd1 vccd1 _20103_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout602 _14635_/X vssd1 vssd1 vccd1 vccd1 _14650_/S sky130_fd_sc_hd__buf_12
X_09914_ _11851_/A _20678_/Q _11851_/C vssd1 vssd1 vccd1 vccd1 _09914_/X sky130_fd_sc_hd__or3_1
XFILLER_104_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout613 _14531_/X vssd1 vssd1 vccd1 vccd1 _14563_/S sky130_fd_sc_hd__buf_12
XFILLER_99_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout624 _13903_/Y vssd1 vssd1 vccd1 vccd1 _13932_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout635 _16887_/A vssd1 vssd1 vccd1 vccd1 _16849_/A sky130_fd_sc_hd__buf_4
XFILLER_259_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout646 _16067_/X vssd1 vssd1 vccd1 vccd1 _16081_/B sky130_fd_sc_hd__buf_6
X_20034_ _20479_/CLK _20034_/D vssd1 vssd1 vccd1 vccd1 _20034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09845_ _12103_/A1 _09843_/X _09844_/X vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__o21ai_1
Xfanout657 _14810_/X vssd1 vssd1 vccd1 vccd1 _15591_/A sky130_fd_sc_hd__buf_8
XFILLER_274_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout668 _14082_/A2 vssd1 vssd1 vccd1 vccd1 _14108_/A2 sky130_fd_sc_hd__buf_6
XFILLER_219_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout679 _14004_/A2 vssd1 vssd1 vccd1 vccd1 _17919_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09776_ _09772_/X _09775_/X _09776_/S vssd1 vssd1 vccd1 vccd1 _09776_/X sky130_fd_sc_hd__mux2_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _21008_/CLK _20936_/D vssd1 vssd1 vccd1 vccd1 _20936_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _21029_/CLK _20867_/D vssd1 vssd1 vccd1 vccd1 _20867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ _10618_/X _10619_/X _12023_/S vssd1 vssd1 vccd1 vccd1 _10620_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20798_ _20861_/CLK _20798_/D vssd1 vssd1 vccd1 vccd1 _20798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10551_ _11228_/A1 _09672_/B _10550_/X _11228_/B1 _19848_/Q vssd1 vssd1 vccd1 vccd1
+ _10551_/X sky130_fd_sc_hd__o32a_1
XFILLER_167_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10482_ _20471_/Q _20311_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _10482_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13270_ _13270_/A _13270_/B _13270_/C vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__and3_1
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ _12396_/A1 _19491_/Q _19459_/Q _12381_/S _12371_/C1 vssd1 vssd1 vccd1 vccd1
+ _12221_/X sky130_fd_sc_hd__a221o_1
XFILLER_135_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ _12152_/A1 _12144_/X _12151_/X _12137_/X vssd1 vssd1 vccd1 vccd1 _12152_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_269_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11103_ _19496_/Q _11189_/B vssd1 vssd1 vccd1 vccd1 _11103_/Y sky130_fd_sc_hd__nor2_1
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_169_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21040_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16960_ _16950_/Y _16959_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16960_/Y sky130_fd_sc_hd__o21bai_4
X_12083_ _12084_/A _20519_/Q _10628_/S _20551_/Q vssd1 vssd1 vccd1 vccd1 _12083_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11034_ _12430_/S _11034_/B vssd1 vssd1 vccd1 vccd1 _11034_/Y sky130_fd_sc_hd__nor2_1
X_15911_ _20940_/Q _16044_/A2 _15910_/X vssd1 vssd1 vccd1 vccd1 _15911_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16891_ _16981_/A1 _15671_/X _16879_/X _16890_/X vssd1 vssd1 vccd1 vccd1 _16891_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_238_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18630_ _18877_/A _18630_/B vssd1 vssd1 vccd1 vccd1 _20930_/D sky130_fd_sc_hd__nor2_1
XFILLER_134_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _19550_/Q _15980_/A2 _15841_/X _17432_/A vssd1 vssd1 vccd1 vccd1 _19550_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _18559_/B _18560_/X _18559_/Y _19048_/A2 vssd1 vssd1 vccd1 vccd1 _18562_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_246_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _21033_/Q _21001_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _15773_/X sky130_fd_sc_hd__mux2_1
XFILLER_264_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12985_ _19221_/Q _13545_/B vssd1 vssd1 vccd1 vccd1 _13559_/B sky130_fd_sc_hd__nand2_1
XFILLER_252_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17512_ _20291_/Q _17522_/B vssd1 vssd1 vccd1 vccd1 _17512_/Y sky130_fd_sc_hd__nand2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _19481_/Q _17939_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19481_/D sky130_fd_sc_hd__mux2_1
XFILLER_261_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18492_ _18598_/A _18492_/B vssd1 vssd1 vccd1 vccd1 _20890_/D sky130_fd_sc_hd__nor2_1
XFILLER_18_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11936_ _19890_/Q _19791_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _11936_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_540 _11204_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_551 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_562 _16815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17443_ _17443_/A _17443_/B _17443_/C _17443_/D vssd1 vssd1 vccd1 vccd1 _17443_/X
+ sky130_fd_sc_hd__or4_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_573 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14655_ _19417_/Q _17871_/A1 _14662_/S vssd1 vssd1 vccd1 vccd1 _19417_/D sky130_fd_sc_hd__mux2_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _20485_/Q _11944_/S _11946_/C1 vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__o21a_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_584 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_595 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ _13605_/A _13605_/B _13605_/Y _13519_/S vssd1 vssd1 vccd1 vccd1 _13606_/X
+ sky130_fd_sc_hd__a211o_1
X_10818_ _20562_/Q _12295_/B vssd1 vssd1 vccd1 vccd1 _10818_/X sky130_fd_sc_hd__or2_1
XFILLER_158_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17374_ _20235_/Q _17378_/A2 _17382_/B1 _20284_/Q _17380_/C1 vssd1 vssd1 vccd1 vccd1
+ _17374_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14586_ _19352_/Q _17938_/A1 _14594_/S vssd1 vssd1 vccd1 vccd1 _19352_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11798_ _15789_/A _15789_/B _11793_/X _11797_/X vssd1 vssd1 vccd1 vccd1 _11798_/X
+ sky130_fd_sc_hd__a211o_1
X_19113_ _20273_/CLK _19113_/D vssd1 vssd1 vccd1 vccd1 _19113_/Q sky130_fd_sc_hd__dfxtp_4
X_16325_ _19717_/Q _16324_/B _18708_/A vssd1 vssd1 vccd1 vccd1 _16326_/B sky130_fd_sc_hd__o21ai_1
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13537_ _16241_/A _13913_/A vssd1 vssd1 vccd1 vccd1 _13537_/Y sky130_fd_sc_hd__nor2_2
X_10749_ _12324_/S _10748_/X _10747_/X _12314_/C1 vssd1 vssd1 vccd1 vccd1 _10749_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19044_ _18305_/Y _19046_/A2 _19017_/X _12553_/B _19048_/C1 vssd1 vssd1 vccd1 vccd1
+ _19044_/X sky130_fd_sc_hd__a221o_1
X_16256_ _19672_/Q _17687_/A1 _16275_/S vssd1 vssd1 vccd1 vccd1 _19672_/D sky130_fd_sc_hd__mux2_1
X_13468_ _13468_/A _13468_/B _13468_/C vssd1 vssd1 vccd1 vccd1 _13468_/Y sky130_fd_sc_hd__nor3_4
XFILLER_185_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15207_ _15348_/B2 _12656_/X _15185_/A _12578_/A _10935_/B vssd1 vssd1 vccd1 vccd1
+ _15208_/C sky130_fd_sc_hd__o221a_1
X_12419_ _10692_/A _20395_/Q _20459_/Q _12268_/S _12419_/C1 vssd1 vssd1 vccd1 vccd1
+ _12419_/X sky130_fd_sc_hd__a221o_1
X_16187_ _16187_/A _16187_/B vssd1 vssd1 vccd1 vccd1 _19617_/D sky130_fd_sc_hd__and2_1
X_13399_ _13393_/Y _13398_/X _13205_/A vssd1 vssd1 vccd1 vccd1 _13399_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ _09480_/Y _15568_/A2 _15322_/B vssd1 vssd1 vccd1 vccd1 _15138_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15069_ _14841_/S _15068_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _15069_/X sky130_fd_sc_hd__o21a_1
X_19946_ _20075_/CLK _19946_/D vssd1 vssd1 vccd1 vccd1 _19946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19877_ _20451_/CLK _19877_/D vssd1 vssd1 vccd1 vccd1 _19877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_268_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09630_ _09630_/A _09630_/B _09630_/C _09630_/D vssd1 vssd1 vccd1 vccd1 _09630_/X
+ sky130_fd_sc_hd__or4_1
X_18828_ _18842_/A _18828_/B vssd1 vssd1 vccd1 vccd1 _20989_/D sky130_fd_sc_hd__nor2_1
XFILLER_95_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09561_ _12708_/A _09734_/B _09561_/C _09561_/D vssd1 vssd1 vccd1 vccd1 _14881_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_270_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18759_ _20979_/Q _18763_/A1 _12982_/C _18758_/X _18476_/A vssd1 vssd1 vccd1 vccd1
+ _20978_/D sky130_fd_sc_hd__o311a_1
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09492_ _19501_/Q vssd1 vssd1 vccd1 vccd1 _12634_/A sky130_fd_sc_hd__clkinv_2
XFILLER_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20721_ _20721_/CLK _20721_/D vssd1 vssd1 vccd1 vccd1 _20721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20652_ _20706_/CLK _20652_/D vssd1 vssd1 vccd1 vccd1 _20652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20583_ _20583_/CLK _20583_/D vssd1 vssd1 vccd1 vccd1 _20583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1408 _11303_/S vssd1 vssd1 vccd1 vccd1 _11042_/B sky130_fd_sc_hd__clkbuf_8
Xfanout1419 _12272_/B2 vssd1 vssd1 vccd1 vccd1 _12268_/S sky130_fd_sc_hd__buf_6
XFILLER_63_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20017_ _20017_/CLK _20017_/D vssd1 vssd1 vccd1 vccd1 _20017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09828_ _09829_/A _19919_/Q _10092_/S _20044_/Q vssd1 vssd1 vccd1 vccd1 _09828_/X
+ sky130_fd_sc_hd__o22a_1
Xfanout498 _17851_/X vssd1 vssd1 vccd1 vccd1 _17883_/S sky130_fd_sc_hd__buf_12
XFILLER_150_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ _20420_/Q _20356_/Q _20648_/Q _20612_/Q _11848_/S0 _12008_/C vssd1 vssd1
+ vccd1 vccd1 _09759_/X sky130_fd_sc_hd__mux4_1
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12771_/C _12771_/D vssd1 vssd1 vccd1 vccd1 _13600_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _12105_/A _12023_/S _11718_/X _11720_/X vssd1 vssd1 vccd1 vccd1 _11721_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_230_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20919_ _21017_/CLK _20919_/D vssd1 vssd1 vccd1 vccd1 _20919_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14440_ _14443_/B vssd1 vssd1 vccd1 vccd1 _14440_/Y sky130_fd_sc_hd__inv_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _13167_/A _13166_/A vssd1 vssd1 vccd1 vccd1 _13418_/A sky130_fd_sc_hd__and2b_4
XFILLER_230_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ _19632_/Q _10603_/B vssd1 vssd1 vccd1 vccd1 _10603_/X sky130_fd_sc_hd__or2_1
X_14371_ _20291_/Q _14431_/A2 _14431_/B1 input232/X vssd1 vssd1 vccd1 vccd1 _14373_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_211_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11583_ _11977_/A1 _20708_/Q _11979_/S _11582_/X vssd1 vssd1 vccd1 vccd1 _11583_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ _09944_/X _16132_/A2 _16109_/X vssd1 vssd1 vccd1 vccd1 _19579_/D sky130_fd_sc_hd__o21a_1
X_13322_ _19224_/Q _13587_/B _12991_/D _19233_/Q vssd1 vssd1 vccd1 vccd1 _13323_/B
+ sky130_fd_sc_hd__a31o_1
X_17090_ _20060_/Q _17649_/A1 _17114_/S vssd1 vssd1 vccd1 vccd1 _20060_/D sky130_fd_sc_hd__mux2_1
X_10534_ _20407_/Q _20343_/Q _20635_/Q _20599_/Q _11203_/S _11290_/C vssd1 vssd1 vccd1
+ vccd1 _10534_/X sky130_fd_sc_hd__mux4_1
XFILLER_183_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16041_ _20753_/Q _16041_/A2 _16041_/B1 _20785_/Q vssd1 vssd1 vccd1 vccd1 _16041_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_109_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10465_ _10465_/A _10465_/B vssd1 vssd1 vccd1 vccd1 _10465_/Y sky130_fd_sc_hd__nand2_1
X_13253_ _13253_/A _13253_/B _13253_/C vssd1 vssd1 vccd1 vccd1 _13253_/X sky130_fd_sc_hd__and3_1
XFILLER_182_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12204_ _11804_/A _11804_/B _12112_/A vssd1 vssd1 vccd1 vccd1 _12206_/C sky130_fd_sc_hd__a21oi_1
X_13184_ _13653_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13184_/X sky130_fd_sc_hd__and2_1
X_10396_ _09829_/A _19345_/Q _20700_/Q _10397_/S _12100_/B1 vssd1 vssd1 vccd1 vccd1
+ _10396_/X sky130_fd_sc_hd__a221o_1
X_19800_ _20061_/CLK _19800_/D vssd1 vssd1 vccd1 vccd1 _19800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12135_ _12135_/A _12135_/B vssd1 vssd1 vccd1 vccd1 _12135_/X sky130_fd_sc_hd__or2_1
X_17992_ _18080_/A _17997_/C vssd1 vssd1 vccd1 vccd1 _17992_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1920 _16179_/A vssd1 vssd1 vccd1 vccd1 _16159_/C1 sky130_fd_sc_hd__buf_4
X_16943_ _16940_/Y _16942_/Y _16822_/A vssd1 vssd1 vccd1 vccd1 _16943_/Y sky130_fd_sc_hd__a21oi_4
X_19731_ _20990_/CLK _19731_/D vssd1 vssd1 vccd1 vccd1 _19731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1931 _14185_/C1 vssd1 vssd1 vccd1 vccd1 _18476_/A sky130_fd_sc_hd__clkbuf_8
X_12066_ _19649_/Q _12070_/S _12043_/X _12071_/S vssd1 vssd1 vccd1 vccd1 _12066_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout1942 _14458_/A vssd1 vssd1 vccd1 vccd1 _16097_/B1 sky130_fd_sc_hd__buf_4
XFILLER_277_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1953 _18418_/A vssd1 vssd1 vccd1 vccd1 _18692_/A sky130_fd_sc_hd__buf_4
XFILLER_265_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ _11015_/Y _11016_/Y _11313_/B vssd1 vssd1 vccd1 vccd1 _11017_/X sky130_fd_sc_hd__a21o_1
Xfanout1964 _18905_/A vssd1 vssd1 vccd1 vccd1 _18960_/A sky130_fd_sc_hd__buf_4
XFILLER_77_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19662_ _20557_/CLK _19662_/D vssd1 vssd1 vccd1 vccd1 _19662_/Q sky130_fd_sc_hd__dfxtp_1
X_16874_ _16884_/S _09528_/Y _16809_/X _16873_/Y vssd1 vssd1 vccd1 vccd1 _16874_/X
+ sky130_fd_sc_hd__o211a_4
Xfanout1975 _18842_/A vssd1 vssd1 vccd1 vccd1 _18856_/A sky130_fd_sc_hd__buf_6
Xfanout1986 _18808_/A vssd1 vssd1 vccd1 vccd1 _16896_/C1 sky130_fd_sc_hd__buf_4
XFILLER_226_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1997 _18086_/A vssd1 vssd1 vccd1 vccd1 _18080_/A sky130_fd_sc_hd__buf_4
XFILLER_253_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15825_ _20745_/Q _15934_/A2 _15934_/B1 _20777_/Q vssd1 vssd1 vccd1 vccd1 _15825_/X
+ sky130_fd_sc_hd__a22o_1
X_18613_ _18502_/X _18621_/A2 _18611_/Y _18612_/Y vssd1 vssd1 vccd1 vccd1 _18614_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_231_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19593_ _19606_/CLK _19593_/D vssd1 vssd1 vccd1 vccd1 _19593_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ _18560_/A _18544_/B vssd1 vssd1 vccd1 vccd1 _18544_/X sky130_fd_sc_hd__or2_1
X_15756_ _15246_/A _15754_/Y _15755_/X _13417_/A _12578_/A vssd1 vssd1 vccd1 vccd1
+ _15756_/X sky130_fd_sc_hd__o32a_1
X_12968_ _19093_/Q _19092_/Q _19091_/Q _12968_/D vssd1 vssd1 vccd1 vccd1 _12975_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_66_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20662_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14707_ _19464_/Q _16608_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19464_/D sky130_fd_sc_hd__mux2_1
XFILLER_261_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18475_ _18589_/B _12557_/Y _13192_/Y _18474_/X vssd1 vssd1 vccd1 vccd1 _18476_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11919_ _12144_/C1 _11908_/X _11911_/X _11918_/X _12152_/A1 vssd1 vssd1 vccd1 vccd1
+ _11919_/X sky130_fd_sc_hd__a311o_1
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15687_ _19720_/Q _15961_/A2 _15961_/B1 _19752_/Q vssd1 vssd1 vccd1 vccd1 _15687_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _12883_/B _12893_/B _12911_/A vssd1 vssd1 vccd1 vccd1 _12900_/B sky130_fd_sc_hd__o21a_1
XANTENNA_370 _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_381 ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_392 _16878_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17426_ _17432_/A _17426_/B vssd1 vssd1 vccd1 vccd1 _20257_/D sky130_fd_sc_hd__and2_1
X_14638_ _19400_/Q _17782_/A1 _14650_/S vssd1 vssd1 vccd1 vccd1 _19400_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17357_ _20227_/Q _17371_/A2 _17356_/X _18418_/A vssd1 vssd1 vccd1 vccd1 _20227_/D
+ sky130_fd_sc_hd__o211a_1
X_14569_ _19335_/Q _17921_/A1 _14599_/S vssd1 vssd1 vccd1 vccd1 _19335_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16308_ _19711_/Q _16308_/B vssd1 vssd1 vccd1 vccd1 _16314_/C sky130_fd_sc_hd__and2_2
XFILLER_147_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17288_ _20201_/Q _17327_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17288_/X sky130_fd_sc_hd__a21o_1
X_19027_ _21032_/Q _19015_/B _19026_/X _18748_/A vssd1 vssd1 vccd1 vccd1 _21032_/D
+ sky130_fd_sc_hd__o211a_1
X_16239_ _13441_/X _16239_/B vssd1 vssd1 vccd1 vccd1 _16239_/X sky130_fd_sc_hd__and2b_1
XFILLER_115_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19929_ _20315_/CLK _19929_/D vssd1 vssd1 vccd1 vccd1 _19929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09613_ _09613_/A _09613_/B _09643_/A vssd1 vssd1 vccd1 vccd1 _09632_/B sky130_fd_sc_hd__or3b_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _19156_/Q _19155_/Q vssd1 vssd1 vccd1 vccd1 _12579_/C sky130_fd_sc_hd__nor2_2
XFILLER_37_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20704_ _20704_/CLK _20704_/D vssd1 vssd1 vccd1 vccd1 _20704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_197_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20635_ _20635_/CLK _20635_/D vssd1 vssd1 vccd1 vccd1 _20635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20566_ _20698_/CLK _20566_/D vssd1 vssd1 vccd1 vccd1 _20566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20497_ _20690_/CLK _20497_/D vssd1 vssd1 vccd1 vccd1 _20497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10250_ _10248_/X _10249_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _10250_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10181_ _10172_/X _10180_/X _10260_/S vssd1 vssd1 vccd1 vccd1 _10181_/X sky130_fd_sc_hd__mux2_2
XFILLER_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1205 _17232_/X vssd1 vssd1 vccd1 vccd1 _17331_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_278_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1216 _14477_/S vssd1 vssd1 vccd1 vccd1 _14469_/S sky130_fd_sc_hd__buf_6
Xfanout1227 _12738_/B vssd1 vssd1 vccd1 vccd1 _15527_/A sky130_fd_sc_hd__buf_4
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1238 _12365_/A2 vssd1 vssd1 vccd1 vccd1 _12155_/A2 sky130_fd_sc_hd__buf_6
Xfanout1249 _17336_/Y vssd1 vssd1 vccd1 vccd1 _17370_/C1 sky130_fd_sc_hd__buf_6
X_13940_ _19144_/Q _13946_/B1 _13906_/X _13220_/Y vssd1 vssd1 vccd1 vccd1 _19144_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13871_ _19089_/Q _13863_/B _13896_/B1 _19155_/Q _16193_/A vssd1 vssd1 vccd1 vccd1
+ _19089_/D sky130_fd_sc_hd__o221a_1
XFILLER_247_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15610_ _15610_/A1 _14841_/X _15610_/B1 vssd1 vssd1 vccd1 vccd1 _15610_/Y sky130_fd_sc_hd__o21ai_2
X_12822_ _13389_/A _12822_/B vssd1 vssd1 vccd1 vccd1 _12822_/Y sky130_fd_sc_hd__nand2_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16590_ _19861_/Q _16592_/A2 _16592_/B1 input33/X vssd1 vssd1 vccd1 vccd1 _16591_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_216_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15541_ _15606_/A1 _15530_/X _15540_/X vssd1 vssd1 vccd1 vccd1 _16851_/B sky130_fd_sc_hd__a21oi_4
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12753_ _19504_/Q _12782_/A _19505_/Q vssd1 vssd1 vccd1 vccd1 _12754_/B sky130_fd_sc_hd__a21oi_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18526_/B vssd1 vssd1 vccd1 vccd1 _18260_/Y sky130_fd_sc_hd__inv_2
X_11704_ _20415_/Q _20351_/Q _20643_/Q _20607_/Q _10622_/S _09834_/C vssd1 vssd1 vccd1
+ vccd1 _11704_/X sky130_fd_sc_hd__mux4_1
XFILLER_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15472_ _15470_/X _15471_/X _15326_/A vssd1 vssd1 vccd1 vccd1 _15472_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_231_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12684_ _19498_/Q _12758_/B vssd1 vssd1 vccd1 vccd1 _12686_/C sky130_fd_sc_hd__nand2_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _20175_/Q _17805_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20175_/D sky130_fd_sc_hd__mux2_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _19524_/Q _14423_/B vssd1 vssd1 vccd1 vccd1 _14426_/C sky130_fd_sc_hd__nor2_1
X_18191_ _20792_/Q _18190_/Y _18236_/S vssd1 vssd1 vccd1 vccd1 _18192_/B sky130_fd_sc_hd__mux2_1
X_11635_ _12102_/A1 _19481_/Q _19449_/Q _12025_/S vssd1 vssd1 vccd1 vccd1 _11635_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17142_ _20110_/Q _17804_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20110_/D sky130_fd_sc_hd__mux2_1
X_14354_ _14354_/A _14354_/B _14354_/C vssd1 vssd1 vccd1 vccd1 _14356_/A sky130_fd_sc_hd__and3_1
XFILLER_195_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11566_ _12191_/C1 _11945_/S _11563_/X _11565_/X vssd1 vssd1 vccd1 vccd1 _11566_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_184_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20685_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13305_ _20965_/Q _13305_/B vssd1 vssd1 vccd1 vccd1 _13305_/Y sky130_fd_sc_hd__nand2_1
X_10517_ _10356_/A _19472_/Q _19440_/Q _10518_/S vssd1 vssd1 vccd1 vccd1 _10517_/X
+ sky130_fd_sc_hd__a22o_1
X_17073_ _20045_/Q _17107_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20045_/D sky130_fd_sc_hd__mux2_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14285_ _14306_/A1 _14284_/X _13357_/X vssd1 vssd1 vccd1 vccd1 _14286_/C sky130_fd_sc_hd__o21ba_1
X_11497_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _13420_/A sky130_fd_sc_hd__and2_4
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_113_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20014_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_170_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16024_ _16024_/A1 _16022_/X _16023_/Y _13181_/A _16052_/B2 vssd1 vssd1 vccd1 vccd1
+ _16024_/X sky130_fd_sc_hd__a32o_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13236_ _13015_/X _13016_/Y _13084_/Y vssd1 vssd1 vccd1 vccd1 _13236_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10448_ _12073_/C1 _10431_/X _10447_/X _12074_/B1 vssd1 vssd1 vccd1 vccd1 _10448_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13167_ _13167_/A _13167_/B vssd1 vssd1 vccd1 vccd1 _13416_/B sky130_fd_sc_hd__or2_4
XFILLER_123_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10379_ input126/X input161/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10379_/X sky130_fd_sc_hd__mux2_8
XFILLER_112_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12118_ _12288_/B _12117_/Y _13431_/A vssd1 vssd1 vccd1 vccd1 _12118_/X sky130_fd_sc_hd__a21o_1
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17975_ _17975_/A _17975_/B vssd1 vssd1 vccd1 vccd1 _20729_/D sky130_fd_sc_hd__nor2_1
X_13098_ _13004_/X _13097_/X _09488_/A vssd1 vssd1 vccd1 vccd1 _13100_/A sky130_fd_sc_hd__o21ai_4
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19714_ _20856_/CLK _19714_/D vssd1 vssd1 vccd1 vccd1 _19714_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1750 _12302_/S vssd1 vssd1 vccd1 vccd1 _12377_/S sky130_fd_sc_hd__buf_6
X_16926_ _16885_/A _16925_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16926_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12049_ _20391_/Q _20455_/Q _12053_/S vssd1 vssd1 vccd1 vccd1 _12049_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1761 _09488_/Y vssd1 vssd1 vccd1 vccd1 _14295_/C1 sky130_fd_sc_hd__buf_2
XFILLER_272_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1772 _13609_/A vssd1 vssd1 vccd1 vccd1 _14244_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1783 _18313_/B vssd1 vssd1 vccd1 vccd1 _18308_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_265_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1794 _18199_/A1 vssd1 vssd1 vccd1 vccd1 _18149_/S sky130_fd_sc_hd__buf_4
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19645_ _20647_/CLK _19645_/D vssd1 vssd1 vccd1 vccd1 _19645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16857_ _17008_/B1 _16854_/X _16856_/X _16875_/B2 vssd1 vssd1 vccd1 vccd1 _16858_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15808_ _15973_/A1 _15807_/X _15795_/Y vssd1 vssd1 vccd1 vccd1 _15808_/Y sky130_fd_sc_hd__a21boi_1
X_19576_ _19590_/CLK _19576_/D vssd1 vssd1 vccd1 vccd1 _19576_/Q sky130_fd_sc_hd__dfxtp_1
X_16788_ _16718_/X _16787_/X _17008_/B1 vssd1 vssd1 vccd1 vccd1 _16788_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18527_ _20902_/Q fanout750/X _18526_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18528_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15739_ _15983_/A _15468_/B _15736_/Y _15738_/X vssd1 vssd1 vccd1 vccd1 _15739_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_179_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18458_ _18767_/A _18458_/B vssd1 vssd1 vccd1 vccd1 _18458_/X sky130_fd_sc_hd__and2_4
XFILLER_21_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17409_ _17460_/A2 _17446_/A _17457_/B _20252_/Q vssd1 vssd1 vccd1 vccd1 _17409_/X
+ sky130_fd_sc_hd__a31o_1
X_18389_ _18389_/A _18389_/B _18389_/C vssd1 vssd1 vccd1 vccd1 _18755_/B sky130_fd_sc_hd__or3_4
X_20420_ _20421_/CLK _20420_/D vssd1 vssd1 vccd1 vccd1 _20420_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_267_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20351_ _20675_/CLK _20351_/D vssd1 vssd1 vccd1 vccd1 _20351_/Q sky130_fd_sc_hd__dfxtp_1
X_20282_ _21026_/CLK _20282_/D vssd1 vssd1 vccd1 vccd1 _20282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_283_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09527_ input48/X vssd1 vssd1 vccd1 vccd1 _09527_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11420_ _19882_/Q _19783_/Q _12124_/S vssd1 vssd1 vccd1 vccd1 _11420_/X sky130_fd_sc_hd__mux2_1
X_20618_ _20686_/CLK _20618_/D vssd1 vssd1 vccd1 vccd1 _20618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11351_ _12230_/A1 _20501_/Q _11359_/S _11350_/X vssd1 vssd1 vccd1 vccd1 _11351_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20549_ _20678_/CLK _20549_/D vssd1 vssd1 vccd1 vccd1 _20549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10302_ _19676_/Q _20164_/Q _10303_/S vssd1 vssd1 vccd1 vccd1 _10302_/X sky130_fd_sc_hd__mux2_1
X_14070_ _19194_/Q _14082_/A2 _14069_/X _14070_/C1 vssd1 vssd1 vccd1 vccd1 _19194_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11282_ _11280_/Y _11281_/Y _11313_/B vssd1 vssd1 vccd1 vccd1 _11282_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ _20968_/Q _20902_/Q vssd1 vssd1 vccd1 vccd1 _13021_/Y sky130_fd_sc_hd__nor2_2
X_10233_ _19638_/Q _19944_/Q _10986_/B vssd1 vssd1 vccd1 vccd1 _10233_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1002 _15021_/A vssd1 vssd1 vccd1 vccd1 _15396_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10164_ _12403_/A1 _13688_/A _12403_/B1 vssd1 vssd1 vccd1 vccd1 _10164_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_117_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1013 _15185_/B vssd1 vssd1 vccd1 vccd1 _16028_/C sky130_fd_sc_hd__buf_4
Xfanout1024 _16720_/X vssd1 vssd1 vccd1 vccd1 _16963_/B1 sky130_fd_sc_hd__buf_6
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1035 _17886_/A1 vssd1 vssd1 vccd1 vccd1 _17780_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 _17782_/A1 vssd1 vssd1 vccd1 vccd1 _16608_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1057 _17891_/A1 vssd1 vssd1 vccd1 vccd1 _17751_/A1 sky130_fd_sc_hd__clkbuf_4
X_14972_ _14972_/A _14972_/B _14972_/C vssd1 vssd1 vccd1 vccd1 _14972_/X sky130_fd_sc_hd__or3_1
X_17760_ _20539_/Q _17900_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20539_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10095_ _10260_/S _10094_/X _12342_/A vssd1 vssd1 vccd1 vccd1 _10095_/X sky130_fd_sc_hd__o21a_1
Xfanout1068 _12107_/A1 vssd1 vssd1 vccd1 vccd1 _12194_/A1 sky130_fd_sc_hd__buf_4
XFILLER_254_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1079 _12577_/X vssd1 vssd1 vccd1 vccd1 _15526_/B sky130_fd_sc_hd__buf_6
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16711_ _16711_/A _16714_/D vssd1 vssd1 vccd1 vccd1 _16711_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13923_ _19127_/Q _13921_/B _13932_/B1 _13610_/X vssd1 vssd1 vccd1 vccd1 _19127_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_263_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17691_ _20475_/Q _17691_/A1 _17706_/S vssd1 vssd1 vccd1 vccd1 _20475_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16642_ _19899_/Q _17679_/A1 _16670_/S vssd1 vssd1 vccd1 vccd1 _19899_/D sky130_fd_sc_hd__mux2_1
XFILLER_274_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19430_ _20704_/CLK _19430_/D vssd1 vssd1 vccd1 vccd1 _19430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13854_ _16598_/A _16594_/B _13853_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_267_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ _12483_/Y _12804_/Y _15795_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12805_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16573_ _16591_/A _16573_/B vssd1 vssd1 vccd1 vccd1 _19852_/D sky130_fd_sc_hd__or2_1
XFILLER_204_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19361_ _20583_/CLK _19361_/D vssd1 vssd1 vccd1 vccd1 _19361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ split3/X _13542_/X _13554_/Y _16240_/A1 vssd1 vssd1 vccd1 vccd1 _13785_/X
+ sky130_fd_sc_hd__a22o_4
X_10997_ _20628_/Q _11169_/B _09688_/A vssd1 vssd1 vccd1 vccd1 _10997_/X sky130_fd_sc_hd__a21o_1
XFILLER_250_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18312_ _18700_/A _18312_/B vssd1 vssd1 vccd1 vccd1 _20816_/D sky130_fd_sc_hd__and2_1
XFILLER_37_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15524_ _15591_/A _15524_/B vssd1 vssd1 vccd1 vccd1 _15524_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ _20047_/CLK _19292_/D vssd1 vssd1 vccd1 vccd1 _19292_/Q sky130_fd_sc_hd__dfxtp_1
X_12736_ _12736_/A _12736_/B _12736_/C vssd1 vssd1 vccd1 vccd1 _12749_/B sky130_fd_sc_hd__and3_1
XFILLER_231_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _19544_/Q _18248_/B vssd1 vssd1 vccd1 vccd1 _18243_/Y sky130_fd_sc_hd__nand2b_2
X_15455_ _15021_/A _15444_/X _15454_/X vssd1 vssd1 vccd1 vccd1 _16824_/B sky130_fd_sc_hd__a21oi_4
X_12667_ _14803_/A1 _12582_/C _12682_/B _12666_/Y vssd1 vssd1 vccd1 vccd1 _12667_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14406_ _14417_/S _14406_/B vssd1 vssd1 vccd1 vccd1 _14406_/X sky130_fd_sc_hd__or2_1
X_18174_ _18199_/A1 _14148_/B _18173_/Y vssd1 vssd1 vccd1 vccd1 _18471_/B sky130_fd_sc_hd__o21ai_4
XFILLER_175_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ _20320_/Q _11641_/S _12013_/S _11945_/S vssd1 vssd1 vccd1 vccd1 _11618_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15386_ _20890_/Q _14971_/A _15566_/B1 _15385_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15386_/X sky130_fd_sc_hd__a221o_1
X_12598_ _19499_/Q _19498_/Q _12680_/B vssd1 vssd1 vccd1 vccd1 _12647_/A sky130_fd_sc_hd__and3_1
X_17125_ _20093_/Q _17927_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20093_/D sky130_fd_sc_hd__mux2_1
XFILLER_117_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14337_ _09488_/A _14336_/X _13274_/Y vssd1 vssd1 vccd1 vccd1 _14338_/C sky130_fd_sc_hd__o21a_1
X_11549_ _20413_/Q _20349_/Q _20641_/Q _20605_/Q _12174_/S _09986_/C vssd1 vssd1 vccd1
+ vccd1 _11549_/X sky130_fd_sc_hd__mux4_1
XFILLER_274_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17056_ _20028_/Q _17683_/A1 _17080_/S vssd1 vssd1 vccd1 vccd1 _20028_/D sky130_fd_sc_hd__mux2_1
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14268_ _19509_/Q _14269_/B vssd1 vssd1 vccd1 vccd1 _14278_/A sky130_fd_sc_hd__and2_1
XFILLER_109_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16007_ _16007_/A _16007_/B _16007_/C vssd1 vssd1 vccd1 vccd1 _16007_/Y sky130_fd_sc_hd__nand3_1
X_13219_ _13139_/A _19242_/Q _13218_/Y vssd1 vssd1 vccd1 vccd1 _13220_/A sky130_fd_sc_hd__a21boi_2
XFILLER_124_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14199_ _14197_/Y _14199_/B vssd1 vssd1 vccd1 vccd1 _14201_/A sky130_fd_sc_hd__and2b_1
XFILLER_152_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17958_ _20723_/Q _17959_/C _17957_/Y vssd1 vssd1 vccd1 vccd1 _20723_/D sky130_fd_sc_hd__o21a_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_81_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _19620_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1580 _11009_/B2 vssd1 vssd1 vccd1 vccd1 _09688_/A sky130_fd_sc_hd__buf_6
X_16909_ input53/X input89/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16909_/X sky130_fd_sc_hd__mux2_8
Xfanout1591 _11008_/A3 vssd1 vssd1 vccd1 vccd1 _09623_/B sky130_fd_sc_hd__buf_8
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17889_ _20660_/Q _17889_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20660_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20583_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19628_ _20085_/CLK _19628_/D vssd1 vssd1 vccd1 vccd1 _19628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19559_ _19560_/CLK _19559_/D vssd1 vssd1 vccd1 vccd1 _19559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20403_ _20759_/CLK _20403_/D vssd1 vssd1 vccd1 vccd1 _20403_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20334_ _20659_/CLK _20334_/D vssd1 vssd1 vccd1 vccd1 _20334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20265_ _20421_/CLK _20265_/D vssd1 vssd1 vccd1 vccd1 _20265_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_115_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20196_ _20688_/CLK _20196_/D vssd1 vssd1 vccd1 vccd1 _20196_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput105 dout0[8] vssd1 vssd1 vccd1 vccd1 _09521_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput116 dout1[18] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput127 dout1[28] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_hd__clkbuf_2
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput138 dout1[38] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__clkbuf_2
XFILLER_248_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput149 dout1[48] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__clkbuf_2
XFILLER_236_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10920_ _11268_/A _20305_/Q _10979_/C vssd1 vssd1 vccd1 vccd1 _10920_/X sky130_fd_sc_hd__and3_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _19499_/Q _10935_/B vssd1 vssd1 vccd1 vccd1 _10851_/Y sky130_fd_sc_hd__nor2_1
XFILLER_112_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13570_ _13570_/A _13570_/B vssd1 vssd1 vccd1 vccd1 _15369_/A sky130_fd_sc_hd__xnor2_4
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _19871_/Q _19772_/Q _11116_/S vssd1 vssd1 vccd1 vccd1 _10782_/X sky130_fd_sc_hd__mux2_1
XFILLER_241_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12521_ _19216_/Q _13334_/A _12533_/A _13602_/A1 vssd1 vssd1 vccd1 vccd1 _12521_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _17251_/A _15239_/X _15452_/S vssd1 vssd1 vccd1 vccd1 _15240_/X sky130_fd_sc_hd__mux2_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap1805 _19694_/Q vssd1 vssd1 vccd1 vccd1 _11241_/S sky130_fd_sc_hd__buf_12
X_12452_ _12286_/A _13182_/A _13178_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _16028_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11403_ _10804_/Y _11319_/X _11323_/Y _13570_/A _10805_/Y vssd1 vssd1 vccd1 vccd1
+ _11772_/A sky130_fd_sc_hd__o311a_4
XFILLER_138_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15171_ _15167_/S _15035_/X _15170_/X vssd1 vssd1 vccd1 vccd1 _15172_/B sky130_fd_sc_hd__o21ai_1
X_12383_ _12383_/A _12383_/B vssd1 vssd1 vccd1 vccd1 _12383_/X sky130_fd_sc_hd__or2_1
XFILLER_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14122_ _19494_/Q _14202_/S _14123_/B vssd1 vssd1 vccd1 vccd1 _14122_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11334_ _11332_/X _11333_/X _12376_/S vssd1 vssd1 vccd1 vccd1 _11334_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14053_ _14107_/A _14107_/B _14053_/C vssd1 vssd1 vccd1 vccd1 _14053_/X sky130_fd_sc_hd__or3_1
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18930_ _21004_/Q _18971_/B vssd1 vssd1 vccd1 vccd1 _18930_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11265_ _11266_/A1 _20493_/Q _10324_/S _20525_/Q vssd1 vssd1 vccd1 vccd1 _11265_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13004_ _13363_/B _12920_/X _13002_/Y _13003_/Y vssd1 vssd1 vccd1 vccd1 _13004_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_234_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10216_ _20133_/Q _20101_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _10216_/X sky130_fd_sc_hd__mux2_1
X_18861_ _20994_/Q _18861_/B vssd1 vssd1 vccd1 vccd1 _18861_/Y sky130_fd_sc_hd__nand2_1
X_11196_ _12332_/A _20658_/Q _12337_/C vssd1 vssd1 vccd1 vccd1 _11196_/X sky130_fd_sc_hd__or3_1
XFILLER_122_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17812_ _17812_/A _17850_/B vssd1 vssd1 vccd1 vccd1 _17813_/C sky130_fd_sc_hd__nor2_1
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _18765_/A _20506_/Q _10152_/S _10146_/X vssd1 vssd1 vccd1 vccd1 _10147_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_267_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18792_ _18581_/Y _18867_/A2 _18791_/X _18901_/S vssd1 vssd1 vccd1 vccd1 _18792_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17743_ _20524_/Q _17917_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20524_/D sky130_fd_sc_hd__mux2_1
X_14955_ _15019_/B _14955_/B _15133_/B vssd1 vssd1 vccd1 vccd1 _14957_/B sky130_fd_sc_hd__and3_2
XFILLER_130_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10078_ _12403_/B1 _10077_/Y _12468_/B _11398_/S vssd1 vssd1 vccd1 vccd1 _10112_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13906_ _16189_/A _13906_/B vssd1 vssd1 vccd1 vccd1 _13906_/X sky130_fd_sc_hd__and2_4
X_17674_ _20460_/Q _17674_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20460_/D sky130_fd_sc_hd__mux2_1
X_14886_ _15035_/S _15494_/B _14836_/X vssd1 vssd1 vccd1 vccd1 _14886_/X sky130_fd_sc_hd__o21a_1
XFILLER_263_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19413_ _20702_/CLK _19413_/D vssd1 vssd1 vccd1 vccd1 _19413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13837_ _17441_/A _17457_/B vssd1 vssd1 vccd1 vccd1 _17438_/B sky130_fd_sc_hd__and2_2
XFILLER_63_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16625_ _19884_/Q _17939_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19884_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16556_ _19844_/Q _16576_/A2 _16576_/B1 input14/X vssd1 vssd1 vccd1 vccd1 _16557_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19344_ _20701_/CLK _19344_/D vssd1 vssd1 vccd1 vccd1 _19344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13768_ _13688_/X _13741_/B _13741_/Y _13689_/X _13767_/X vssd1 vssd1 vccd1 vccd1
+ _13769_/B sky130_fd_sc_hd__o221a_4
X_15507_ _20734_/Q _16041_/A2 _16041_/B1 _20766_/Q vssd1 vssd1 vccd1 vccd1 _15507_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12719_ _12479_/A _12730_/A2 _12731_/B _12718_/X vssd1 vssd1 vccd1 vccd1 _12719_/X
+ sky130_fd_sc_hd__a211o_1
X_19275_ _20181_/CLK _19275_/D vssd1 vssd1 vccd1 vccd1 _19275_/Q sky130_fd_sc_hd__dfxtp_1
X_16487_ _19796_/Q _17707_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19796_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13699_ _13735_/A _13735_/B vssd1 vssd1 vccd1 vccd1 _13699_/Y sky130_fd_sc_hd__nor2_1
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18226_ _20799_/Q _18225_/Y _18236_/S vssd1 vssd1 vccd1 vccd1 _18227_/B sky130_fd_sc_hd__mux2_1
X_15438_ _15066_/S _15255_/X _15610_/B1 vssd1 vssd1 vccd1 vccd1 _15438_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_129_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18157_ _18157_/A _18157_/B _18690_/A _18157_/D vssd1 vssd1 vccd1 vccd1 _18157_/Y
+ sky130_fd_sc_hd__nor4_4
X_15369_ _15369_/A _15494_/B vssd1 vssd1 vccd1 vccd1 _15369_/X sky130_fd_sc_hd__or2_1
XFILLER_157_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17108_ _20078_/Q _17876_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20078_/D sky130_fd_sc_hd__mux2_1
X_18088_ _18094_/A _18093_/C vssd1 vssd1 vccd1 vccd1 _18088_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17039_ _20017_/Q _12928_/C _17040_/S vssd1 vssd1 vccd1 vccd1 _20017_/D sky130_fd_sc_hd__mux2_1
X_09930_ _11946_/A1 _19355_/Q _20710_/Q _09931_/S _11946_/C1 vssd1 vssd1 vccd1 vccd1
+ _09930_/X sky130_fd_sc_hd__a221o_1
XFILLER_132_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20050_ _20681_/CLK _20050_/D vssd1 vssd1 vccd1 vccd1 _20050_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout806 _14525_/B vssd1 vssd1 vccd1 vccd1 _13612_/A sky130_fd_sc_hd__clkbuf_8
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _09861_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09862_/A sky130_fd_sc_hd__and2_2
Xfanout817 _12562_/A vssd1 vssd1 vccd1 vccd1 _13740_/B sky130_fd_sc_hd__buf_8
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout828 _13735_/A vssd1 vssd1 vccd1 vccd1 _13685_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_258_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout839 _18491_/B2 vssd1 vssd1 vccd1 vccd1 _18458_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_274_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _20387_/Q _20451_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _09792_/X sky130_fd_sc_hd__mux2_1
XFILLER_218_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _21018_/CLK _20952_/D vssd1 vssd1 vccd1 vccd1 _20952_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_242_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20883_ _20980_/CLK _20883_/D vssd1 vssd1 vccd1 vccd1 _20883_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_216_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20714_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20317_ _20573_/CLK _20317_/D vssd1 vssd1 vccd1 vccd1 _20317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11050_ _11313_/B _12658_/A _11019_/Y vssd1 vssd1 vccd1 vccd1 _11054_/B sky130_fd_sc_hd__o21bai_4
X_20248_ _20296_/CLK _20248_/D vssd1 vssd1 vccd1 vccd1 _20248_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10001_ _20321_/Q _11944_/S _10000_/X vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__a21o_1
XFILLER_277_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20179_ _20179_/CLK _20179_/D vssd1 vssd1 vccd1 vccd1 _20179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _19117_/Q _14802_/A2 _14739_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _19494_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _12194_/A1 _17877_/A1 _11951_/X _12194_/B2 vssd1 vssd1 vccd1 vccd1 _15870_/A
+ sky130_fd_sc_hd__a22o_2
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10903_ _19271_/Q _11169_/B _09688_/A vssd1 vssd1 vccd1 vccd1 _10903_/X sky130_fd_sc_hd__a21o_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14671_ _19430_/Q _17920_/A1 _14685_/S vssd1 vssd1 vccd1 vccd1 _19430_/D sky130_fd_sc_hd__mux2_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _11882_/Y _11798_/X _11883_/C _11883_/D vssd1 vssd1 vccd1 vccd1 _11883_/X
+ sky130_fd_sc_hd__and4bb_2
XFILLER_260_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16410_ _19748_/Q _19749_/Q _16410_/C vssd1 vssd1 vccd1 vccd1 _16412_/B sky130_fd_sc_hd__and3_4
XFILLER_205_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13622_ _13481_/A _13361_/A _13428_/C _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13622_/X
+ sky130_fd_sc_hd__a22o_2
X_10834_ _20630_/Q _20594_/Q _12389_/S vssd1 vssd1 vccd1 vccd1 _10834_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17390_ _20243_/Q _17390_/A2 _17530_/A2 _20292_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17390_/X sky130_fd_sc_hd__a221o_1
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16341_ _19723_/Q _16340_/B _18720_/A vssd1 vssd1 vccd1 vccd1 _16342_/B sky130_fd_sc_hd__o21ai_1
X_13553_ _13582_/A _19221_/Q _14184_/A vssd1 vssd1 vccd1 vccd1 _13915_/A sky130_fd_sc_hd__a21oi_4
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10765_ _19176_/Q _11367_/B _10764_/Y _11189_/B vssd1 vssd1 vccd1 vccd1 _10799_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19060_ _20405_/Q vssd1 vssd1 vccd1 vccd1 _20405_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_197_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ _12504_/A _12504_/B _19165_/Q vssd1 vssd1 vccd1 vccd1 _12511_/B sky130_fd_sc_hd__or3_1
XFILLER_13_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16272_ _19688_/Q _17946_/A1 _16272_/S vssd1 vssd1 vccd1 vccd1 _19688_/D sky130_fd_sc_hd__mux2_1
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _12676_/B _13483_/Y _12664_/C vssd1 vssd1 vccd1 vccd1 _13484_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10696_ _10690_/X _10695_/X _12415_/S vssd1 vssd1 vccd1 vccd1 _10696_/X sky130_fd_sc_hd__mux2_2
XFILLER_139_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18011_ _20742_/Q _20741_/Q _18011_/C vssd1 vssd1 vccd1 vccd1 _18013_/B sky130_fd_sc_hd__and3_1
X_15223_ _14841_/S _15157_/A _14885_/X vssd1 vssd1 vccd1 vccd1 _15223_/X sky130_fd_sc_hd__o21a_2
X_12435_ _12436_/A _12443_/B vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__nor2_2
XFILLER_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15154_ _19529_/Q _15492_/A _15153_/Y _16159_/C1 vssd1 vssd1 vccd1 vccd1 _19529_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12366_ _12366_/A1 _10290_/B _10037_/B vssd1 vssd1 vccd1 vccd1 _12366_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput409 _19993_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_ack_o sky130_fd_sc_hd__buf_4
X_14105_ _14105_/A _14107_/B _14105_/C vssd1 vssd1 vccd1 vccd1 _14105_/X sky130_fd_sc_hd__or3_1
XFILLER_5_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11317_ _13482_/A _11781_/B _11136_/X vssd1 vssd1 vccd1 vccd1 _11780_/B sky130_fd_sc_hd__a21o_1
X_15085_ _20947_/Q _15568_/A2 _15568_/B1 _20819_/Q _15084_/X vssd1 vssd1 vccd1 vccd1
+ _15085_/X sky130_fd_sc_hd__a221o_2
X_19962_ _20624_/CLK _19962_/D vssd1 vssd1 vccd1 vccd1 _19962_/Q sky130_fd_sc_hd__dfxtp_1
X_12297_ _12371_/A1 _19365_/Q _20720_/Q _12296_/S _12304_/C1 vssd1 vssd1 vccd1 vccd1
+ _12297_/X sky130_fd_sc_hd__a221o_1
X_14036_ _19211_/Q _14103_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _14036_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18913_ _19106_/Q _18974_/A2 _12591_/X _13414_/Y vssd1 vssd1 vccd1 vccd1 _18913_/X
+ sky130_fd_sc_hd__o2bb2a_2
X_11248_ _20118_/Q _20086_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _11248_/X sky130_fd_sc_hd__mux2_1
X_19893_ _20677_/CLK _19893_/D vssd1 vssd1 vccd1 vccd1 _19893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_267_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18844_ _18968_/A _18844_/B vssd1 vssd1 vccd1 vccd1 _18844_/Y sky130_fd_sc_hd__nand2_1
X_11179_ _18765_/A _19335_/Q _20690_/Q _10924_/S _12519_/C vssd1 vssd1 vccd1 vccd1
+ _11179_/X sky130_fd_sc_hd__a221o_1
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18775_ _19118_/Q _18774_/Y _18867_/A2 _18570_/Y vssd1 vssd1 vccd1 vccd1 _18775_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_83_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _15219_/Y _15981_/X _15982_/X _15986_/X vssd1 vssd1 vccd1 vccd1 _15987_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17726_ _20507_/Q _17900_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20507_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14938_ _15019_/B _14967_/A vssd1 vssd1 vccd1 vccd1 _14938_/Y sky130_fd_sc_hd__nand2_2
XFILLER_224_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17657_ _20443_/Q _17657_/A1 _17657_/S vssd1 vssd1 vccd1 vccd1 _20443_/D sky130_fd_sc_hd__mux2_1
X_14869_ _11138_/B _12279_/Y _14870_/S vssd1 vssd1 vccd1 vccd1 _14869_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _19867_/Q _16608_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19867_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17588_ _20346_/Q _17899_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20346_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19327_ _20047_/CLK _19327_/D vssd1 vssd1 vccd1 vccd1 _19327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16539_ _16593_/A _16539_/B vssd1 vssd1 vccd1 vccd1 _19835_/D sky130_fd_sc_hd__or2_1
XFILLER_149_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19258_ _21016_/CLK _19258_/D vssd1 vssd1 vccd1 vccd1 _19258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18209_ _18209_/A1 _14218_/B _18208_/Y vssd1 vssd1 vccd1 vccd1 _18496_/B sky130_fd_sc_hd__o21ai_4
X_19189_ _20341_/CLK _19189_/D vssd1 vssd1 vccd1 vccd1 _19189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20102_ _20573_/CLK _20102_/D vssd1 vssd1 vccd1 vccd1 _20102_/Q sky130_fd_sc_hd__dfxtp_1
X_09913_ _11851_/A _20514_/Q _12182_/S _20546_/Q vssd1 vssd1 vccd1 vccd1 _09913_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_160_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout603 _14601_/X vssd1 vssd1 vccd1 vccd1 _14630_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_59_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout614 _14531_/X vssd1 vssd1 vccd1 vccd1 _14562_/S sky130_fd_sc_hd__buf_8
XFILLER_259_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout625 _14043_/B1 vssd1 vssd1 vccd1 vccd1 _14040_/B1 sky130_fd_sc_hd__buf_4
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout636 _17011_/B1 vssd1 vssd1 vccd1 vccd1 _16887_/A sky130_fd_sc_hd__buf_4
X_20033_ _20539_/CLK _20033_/D vssd1 vssd1 vccd1 vccd1 _20033_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout647 _16077_/B vssd1 vssd1 vccd1 vccd1 _16079_/B sky130_fd_sc_hd__buf_4
XFILLER_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09844_ _09829_/A _19356_/Q _20711_/Q _10397_/S _12100_/B1 vssd1 vssd1 vccd1 vccd1
+ _09844_/X sky130_fd_sc_hd__a221o_1
XFILLER_259_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout658 _14737_/X vssd1 vssd1 vccd1 vccd1 _14801_/B sky130_fd_sc_hd__buf_4
XFILLER_101_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout669 _14044_/Y vssd1 vssd1 vccd1 vccd1 _14082_/A2 sky130_fd_sc_hd__buf_8
XFILLER_246_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09775_ _12015_/A1 _09774_/X _09773_/X vssd1 vssd1 vccd1 vccd1 _09775_/X sky130_fd_sc_hd__o21a_1
XFILLER_274_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ _21000_/CLK _20935_/D vssd1 vssd1 vccd1 vccd1 _20935_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20866_ _20962_/CLK _20866_/D vssd1 vssd1 vccd1 vccd1 _20866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20797_ _20861_/CLK _20797_/D vssd1 vssd1 vccd1 vccd1 _20797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10550_ input115/X input150/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10550_/X sky130_fd_sc_hd__mux2_8
XFILLER_128_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10481_ _11259_/S _10479_/X _10480_/X vssd1 vssd1 vccd1 vccd1 _10481_/X sky130_fd_sc_hd__o21a_1
XFILLER_185_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12220_ _19894_/Q _19795_/Q _12381_/S vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ _12151_/A1 _12150_/X _12147_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _12151_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11102_ _11100_/X _11101_/Y _11313_/B vssd1 vssd1 vccd1 vccd1 _11102_/X sky130_fd_sc_hd__a21o_1
XFILLER_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12082_ _12080_/X _12081_/X _12082_/S vssd1 vssd1 vccd1 vccd1 _12082_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11033_ _11031_/X _11032_/X _11033_/S vssd1 vssd1 vccd1 vccd1 _11034_/B sky130_fd_sc_hd__mux2_1
X_15910_ _20908_/Q _15937_/A2 _16043_/B1 _15909_/X _15937_/C1 vssd1 vssd1 vccd1 vccd1
+ _15910_/X sky130_fd_sc_hd__a221o_1
XFILLER_238_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16890_ _19232_/Q _16980_/A2 _16980_/B1 _19101_/Q _16889_/X vssd1 vssd1 vccd1 vccd1
+ _16890_/X sky130_fd_sc_hd__o221a_1
XFILLER_277_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _15841_/A _15841_/B _15814_/A vssd1 vssd1 vccd1 vccd1 _15841_/X sky130_fd_sc_hd__or3b_2
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_138_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _19698_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _18560_/A _18560_/B vssd1 vssd1 vccd1 vccd1 _18560_/X sky130_fd_sc_hd__or2_1
XFILLER_252_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _19220_/Q _19219_/Q _19218_/Q _13498_/B vssd1 vssd1 vccd1 vccd1 _13545_/B
+ sky130_fd_sc_hd__and4_2
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _20871_/Q _16018_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15772_/X sky130_fd_sc_hd__o21ba_1
XFILLER_264_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17511_ _17525_/A1 _17510_/Y _17430_/A vssd1 vssd1 vccd1 vccd1 _20290_/D sky130_fd_sc_hd__a21oi_1
X_11935_ _09752_/A _19487_/Q _19455_/Q _11936_/S _12016_/C1 vssd1 vssd1 vccd1 vccd1
+ _11935_/X sky130_fd_sc_hd__a221o_1
X_14723_ _19480_/Q _17938_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19480_/D sky130_fd_sc_hd__mux2_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ _20890_/Q fanout753/X _18490_/X _18491_/B2 vssd1 vssd1 vccd1 vccd1 _18492_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_530 _14563_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_541 _12426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17442_ _17442_/A _17446_/B vssd1 vssd1 vccd1 vccd1 _17443_/D sky130_fd_sc_hd__nor2_1
X_14654_ _19416_/Q _17938_/A1 _14662_/S vssd1 vssd1 vccd1 vccd1 _19416_/D sky130_fd_sc_hd__mux2_1
XANTENNA_552 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _11948_/A1 _11865_/X _11864_/X vssd1 vssd1 vccd1 vccd1 _11866_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_563 _16860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_574 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_585 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_596 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13605_ _13605_/A _13605_/B vssd1 vssd1 vccd1 vccd1 _13605_/Y sky130_fd_sc_hd__nor2_1
X_10817_ _12230_/A1 _19467_/Q _19435_/Q _12389_/S _09695_/A vssd1 vssd1 vccd1 vccd1
+ _10817_/X sky130_fd_sc_hd__a221o_1
XFILLER_232_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14585_ _19351_/Q _17937_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19351_/D sky130_fd_sc_hd__mux2_1
X_17373_ _20235_/Q _17381_/A2 _17372_/X _14482_/A vssd1 vssd1 vccd1 vccd1 _20235_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11797_ _15652_/A _15652_/B _15734_/B _15734_/A _15582_/A vssd1 vssd1 vccd1 vccd1
+ _11797_/X sky130_fd_sc_hd__a221o_1
XFILLER_41_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19112_ _20273_/CLK _19112_/D vssd1 vssd1 vccd1 vccd1 _19112_/Q sky130_fd_sc_hd__dfxtp_4
X_16324_ _19717_/Q _16324_/B vssd1 vssd1 vccd1 vccd1 _16330_/C sky130_fd_sc_hd__and2_4
XFILLER_201_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13536_ _18763_/A1 _19220_/Q _14173_/A vssd1 vssd1 vccd1 vccd1 _13913_/A sky130_fd_sc_hd__a21oi_4
X_10748_ _20631_/Q _20595_/Q _12313_/S vssd1 vssd1 vccd1 vccd1 _10748_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19043_ _21040_/Q _19049_/A2 _19042_/X _18736_/A vssd1 vssd1 vccd1 vccd1 _21040_/D
+ sky130_fd_sc_hd__o211a_1
X_16255_ _19671_/Q _17861_/A1 _16272_/S vssd1 vssd1 vccd1 vccd1 _19671_/D sky130_fd_sc_hd__mux2_1
X_13467_ _20015_/Q _20016_/Q _20017_/Q _20018_/Q vssd1 vssd1 vccd1 vccd1 _13468_/C
+ sky130_fd_sc_hd__or4_4
X_10679_ _10664_/X _10678_/X _12401_/A1 vssd1 vssd1 vccd1 vccd1 _10679_/X sky130_fd_sc_hd__a21o_2
XFILLER_174_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15206_ _15246_/A _15206_/B _15206_/C vssd1 vssd1 vccd1 vccd1 _15208_/B sky130_fd_sc_hd__or3_1
X_12418_ _12420_/B1 _12417_/X _12416_/X vssd1 vssd1 vccd1 vccd1 _12418_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_173_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16186_ _19617_/Q _15916_/X _16190_/S vssd1 vssd1 vccd1 vccd1 _16187_/B sky130_fd_sc_hd__mux2_1
X_13398_ _13395_/Y _13396_/X _13397_/Y _18651_/B vssd1 vssd1 vccd1 vccd1 _13398_/X
+ sky130_fd_sc_hd__o211a_2
X_15137_ _20820_/Q _15388_/S _15135_/X _15136_/X _15568_/A2 vssd1 vssd1 vccd1 vccd1
+ _15137_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12349_ _11118_/A _12345_/X _11384_/S vssd1 vssd1 vccd1 vccd1 _12349_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15068_ _14885_/B _15067_/X _15254_/S vssd1 vssd1 vccd1 vccd1 _15068_/X sky130_fd_sc_hd__mux2_1
X_19945_ _20673_/CLK _19945_/D vssd1 vssd1 vccd1 vccd1 _19945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14019_ _12513_/D _14043_/A2 _14034_/B1 _14018_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1
+ _19173_/D sky130_fd_sc_hd__o221a_1
XFILLER_141_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19876_ _20472_/CLK _19876_/D vssd1 vssd1 vccd1 vccd1 _19876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18827_ _18493_/X _18861_/B _18825_/X _18826_/Y vssd1 vssd1 vccd1 vccd1 _18828_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09560_ _12708_/A _09734_/B _09561_/C _09561_/D vssd1 vssd1 vccd1 vccd1 _09560_/X
+ sky130_fd_sc_hd__or4_1
X_18758_ _20978_/Q _18756_/Y _18757_/X vssd1 vssd1 vccd1 vccd1 _18758_/X sky130_fd_sc_hd__a21o_1
XFILLER_209_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17709_ _19095_/Q _19094_/Q _17709_/C vssd1 vssd1 vccd1 vccd1 _17850_/B sky130_fd_sc_hd__or3_2
XFILLER_247_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09491_ _19139_/Q vssd1 vssd1 vccd1 vccd1 _09491_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18689_ _18980_/A _18689_/B vssd1 vssd1 vccd1 vccd1 _20945_/D sky130_fd_sc_hd__nor2_1
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20720_ _20720_/CLK _20720_/D vssd1 vssd1 vccd1 vccd1 _20720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20651_ _20683_/CLK _20651_/D vssd1 vssd1 vccd1 vccd1 _20651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20582_ _20714_/CLK _20582_/D vssd1 vssd1 vccd1 vccd1 _20582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1409 _10174_/S vssd1 vssd1 vccd1 vccd1 _11303_/S sky130_fd_sc_hd__buf_6
XFILLER_120_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20016_ _20017_/CLK _20016_/D vssd1 vssd1 vccd1 vccd1 _20016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09827_ _11981_/C1 _16063_/B2 _09826_/X vssd1 vssd1 vccd1 vccd1 _09861_/A sky130_fd_sc_hd__a21oi_2
XFILLER_59_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout488 _17946_/S vssd1 vssd1 vccd1 vccd1 _17948_/S sky130_fd_sc_hd__buf_12
XFILLER_86_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout499 _17851_/X vssd1 vssd1 vccd1 vccd1 _17882_/S sky130_fd_sc_hd__buf_6
XFILLER_86_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09758_ _19389_/Q _12085_/A2 _09756_/X _12190_/C1 _09757_/X vssd1 vssd1 vccd1 vccd1
+ _09758_/X sky130_fd_sc_hd__o221a_1
XFILLER_234_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _09689_/A _10152_/S _09689_/C _09689_/D vssd1 vssd1 vccd1 vccd1 _09689_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _12105_/A _12091_/S _11719_/X _12088_/S vssd1 vssd1 vccd1 vccd1 _11720_/X
+ sky130_fd_sc_hd__a31o_1
X_20918_ _20949_/CLK _20918_/D vssd1 vssd1 vccd1 vccd1 _20918_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11651_ _11651_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__or2_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20849_ _21043_/CLK _20849_/D vssd1 vssd1 vccd1 vccd1 _20849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10602_ _20063_/Q _10628_/S _10601_/X vssd1 vssd1 vccd1 vccd1 _10602_/X sky130_fd_sc_hd__a21o_1
X_14370_ _19239_/Q _14438_/A2 _14369_/X _18752_/A vssd1 vssd1 vccd1 vccd1 _19239_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11582_ _11977_/A1 _11983_/A1 _19353_/Q _12129_/S vssd1 vssd1 vccd1 vccd1 _11582_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_70_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ _13321_/A _13321_/B _13321_/C vssd1 vssd1 vccd1 vccd1 _13321_/Y sky130_fd_sc_hd__nand3_1
XFILLER_195_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10533_ _19376_/Q _11291_/A2 _10531_/X _11291_/B2 _10532_/X vssd1 vssd1 vccd1 vccd1
+ _10533_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16040_ _21043_/Q _21011_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _16040_/X sky130_fd_sc_hd__mux2_1
X_13252_ _13389_/B _13389_/C _13389_/A vssd1 vssd1 vccd1 vccd1 _13253_/C sky130_fd_sc_hd__o21ai_4
XFILLER_108_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10464_ _19577_/Q _10463_/X _11240_/S vssd1 vssd1 vccd1 vccd1 _10465_/B sky130_fd_sc_hd__mux2_1
XFILLER_89_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12203_ _12286_/A _12203_/B vssd1 vssd1 vccd1 vccd1 _15955_/A sky130_fd_sc_hd__and2_1
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13183_ _13183_/A _13183_/B vssd1 vssd1 vccd1 vccd1 _13183_/Y sky130_fd_sc_hd__xnor2_4
X_10395_ _10390_/X _10394_/X _12850_/A1 vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__a21o_1
X_12134_ _12132_/X _12133_/X _12134_/S vssd1 vssd1 vccd1 vccd1 _12135_/B sky130_fd_sc_hd__mux2_1
XFILLER_269_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17991_ _20735_/Q _20734_/Q _17991_/C vssd1 vssd1 vccd1 vccd1 _17997_/C sky130_fd_sc_hd__and3_2
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19730_ _20990_/CLK _19730_/D vssd1 vssd1 vccd1 vccd1 _19730_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16942_ _16885_/A _16941_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16942_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_145_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1910 _18726_/A vssd1 vssd1 vccd1 vccd1 _14772_/C1 sky130_fd_sc_hd__clkbuf_4
X_12065_ _09806_/S _12064_/X _12063_/X _12068_/C1 vssd1 vssd1 vccd1 vccd1 _12065_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout1921 _15288_/C1 vssd1 vssd1 vccd1 vccd1 _16179_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1932 _18702_/A vssd1 vssd1 vccd1 vccd1 _18985_/A sky130_fd_sc_hd__buf_4
XFILLER_278_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1943 _13890_/C1 vssd1 vssd1 vccd1 vccd1 _14458_/A sky130_fd_sc_hd__buf_4
Xfanout1954 _18422_/A vssd1 vssd1 vccd1 vccd1 _18418_/A sky130_fd_sc_hd__clkbuf_4
X_11016_ _19173_/Q _11281_/B vssd1 vssd1 vccd1 vccd1 _11016_/Y sky130_fd_sc_hd__nand2_1
XFILLER_238_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19661_ _19697_/CLK _19661_/D vssd1 vssd1 vccd1 vccd1 _19661_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_237_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16873_ _16884_/S input84/X vssd1 vssd1 vccd1 vccd1 _16873_/Y sky130_fd_sc_hd__nand2_1
Xfanout1965 _18112_/A vssd1 vssd1 vccd1 vccd1 _18966_/A sky130_fd_sc_hd__buf_4
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1976 _18842_/A vssd1 vssd1 vccd1 vccd1 _18863_/A sky130_fd_sc_hd__buf_4
Xfanout1987 _18808_/A vssd1 vssd1 vccd1 vccd1 _18795_/A sky130_fd_sc_hd__buf_2
Xfanout1998 fanout2002/X vssd1 vssd1 vccd1 vccd1 _18086_/A sky130_fd_sc_hd__buf_4
XFILLER_237_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18612_ _19506_/Q _18612_/B vssd1 vssd1 vccd1 vccd1 _18612_/Y sky130_fd_sc_hd__nand2_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15824_ _19725_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15824_/X sky130_fd_sc_hd__or2_1
XFILLER_253_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19592_ _19606_/CLK _19592_/D vssd1 vssd1 vccd1 vccd1 _19592_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _18966_/A _18543_/B vssd1 vssd1 vccd1 vccd1 _20907_/D sky130_fd_sc_hd__nor2_1
X_12967_ _19099_/Q _12967_/B _19095_/Q _19094_/Q vssd1 vssd1 vccd1 vccd1 _12968_/D
+ sky130_fd_sc_hd__or4_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15755_ _16051_/A1 _15741_/X _16051_/B1 vssd1 vssd1 vccd1 vccd1 _15755_/X sky130_fd_sc_hd__o21a_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14706_ _19463_/Q _17678_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19463_/D sky130_fd_sc_hd__mux2_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _12151_/A1 _11917_/X _11914_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _11918_/X
+ sky130_fd_sc_hd__o211a_1
X_18474_ _18473_/Y _20885_/Q _18474_/S vssd1 vssd1 vccd1 vccd1 _18474_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_360 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12898_ _12877_/B _12887_/B _12911_/A vssd1 vssd1 vccd1 vccd1 _13221_/B sky130_fd_sc_hd__o21a_1
X_15686_ _15686_/A _16037_/B vssd1 vssd1 vccd1 vccd1 _15686_/Y sky130_fd_sc_hd__nor2_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_371 _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_382 _15218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17425_ _20257_/Q _20250_/Q _17433_/S vssd1 vssd1 vccd1 vccd1 _17426_/B sky130_fd_sc_hd__mux2_1
X_14637_ _19399_/Q _17921_/A1 _14650_/S vssd1 vssd1 vccd1 vccd1 _19399_/D sky130_fd_sc_hd__mux2_1
XANTENNA_393 _15662_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11849_ _11847_/X _11848_/X _11849_/S vssd1 vssd1 vccd1 vccd1 _11849_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17356_ _20226_/Q _17356_/A2 _17362_/B1 _20275_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17356_/X sky130_fd_sc_hd__a221o_1
XFILLER_193_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14568_ _19334_/Q _17780_/A1 _14599_/S vssd1 vssd1 vccd1 vccd1 _19334_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20539_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_174_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16307_ _18054_/A _16307_/B _16308_/B vssd1 vssd1 vccd1 vccd1 _19710_/D sky130_fd_sc_hd__nor3_1
XFILLER_174_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13519_ _13518_/X _20950_/Q _13519_/S vssd1 vssd1 vccd1 vccd1 _13519_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17287_ _17287_/A _17290_/B _17290_/C vssd1 vssd1 vccd1 vccd1 _17287_/X sky130_fd_sc_hd__and3_1
XFILLER_173_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14499_ _19277_/Q _17896_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19277_/D sky130_fd_sc_hd__mux2_1
XFILLER_256_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19026_ _18260_/Y _19046_/A2 _19048_/B1 _12550_/A _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19026_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16238_ _16240_/A1 _16237_/X _19695_/D vssd1 vssd1 vccd1 vccd1 _19657_/D sky130_fd_sc_hd__o21a_2
XFILLER_173_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16169_ _16189_/A _16169_/B vssd1 vssd1 vccd1 vccd1 _19608_/D sky130_fd_sc_hd__and2_1
XFILLER_173_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19928_ _20085_/CLK _19928_/D vssd1 vssd1 vccd1 vccd1 _19928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19859_ _20017_/CLK _19859_/D vssd1 vssd1 vccd1 vccd1 _19859_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09612_ _09686_/A _12976_/B _09686_/C vssd1 vssd1 vccd1 vccd1 _09612_/X sky130_fd_sc_hd__or3_4
XFILLER_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09543_ _12480_/B _13867_/A vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__nand2_4
XFILLER_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20703_ _20703_/CLK _20703_/D vssd1 vssd1 vccd1 vccd1 _20703_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20634_ _20698_/CLK _20634_/D vssd1 vssd1 vccd1 vccd1 _20634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20565_ _20565_/CLK _20565_/D vssd1 vssd1 vccd1 vccd1 _20565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20496_ _20667_/CLK _20496_/D vssd1 vssd1 vccd1 vccd1 _20496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10180_ _11375_/S _10175_/X _10179_/X vssd1 vssd1 vccd1 vccd1 _10180_/X sky130_fd_sc_hd__o21a_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1206 _17232_/X vssd1 vssd1 vccd1 vccd1 _17328_/A2 sky130_fd_sc_hd__buf_4
XFILLER_182_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1217 _14483_/S vssd1 vssd1 vccd1 vccd1 _14477_/S sky130_fd_sc_hd__buf_8
Xfanout1228 _12482_/Y vssd1 vssd1 vccd1 vccd1 _12738_/B sky130_fd_sc_hd__buf_4
Xfanout1239 _12365_/A2 vssd1 vssd1 vccd1 vccd1 _09613_/A sky130_fd_sc_hd__buf_6
XFILLER_275_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13870_ _19088_/Q _13902_/B _13869_/Y _16167_/C1 vssd1 vssd1 vccd1 vccd1 _19088_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12821_ _13264_/A _13362_/A _13253_/B vssd1 vssd1 vccd1 vccd1 _12822_/B sky130_fd_sc_hd__nor3_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15540_ _19715_/Q _15395_/S _15539_/X vssd1 vssd1 vccd1 vccd1 _15540_/X sky130_fd_sc_hd__o21a_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _12752_/A _12752_/B vssd1 vssd1 vccd1 vccd1 _12752_/Y sky130_fd_sc_hd__nand2_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11703_ _11701_/X _11702_/X _11718_/S vssd1 vssd1 vccd1 vccd1 _11703_/X sky130_fd_sc_hd__mux2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15471_ _10456_/B _12466_/Y _12468_/X _10453_/A _15465_/Y vssd1 vssd1 vccd1 vccd1
+ _15471_/X sky130_fd_sc_hd__o221a_1
XFILLER_242_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12683_ _12681_/X _12682_/Y _12708_/B vssd1 vssd1 vccd1 vccd1 _12686_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _19524_/Q _14423_/B vssd1 vssd1 vccd1 vccd1 _14432_/A sky130_fd_sc_hd__and2_1
X_17210_ _20174_/Q _17804_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20174_/D sky130_fd_sc_hd__mux2_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _19884_/Q _11641_/S _11708_/B _11632_/X _11633_/X vssd1 vssd1 vccd1 vccd1
+ _11634_/X sky130_fd_sc_hd__a311o_1
X_18190_ _18483_/B vssd1 vssd1 vccd1 vccd1 _18190_/Y sky130_fd_sc_hd__inv_2
XFILLER_230_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14353_ _14361_/A _14353_/B vssd1 vssd1 vccd1 vccd1 _14354_/C sky130_fd_sc_hd__or2_1
X_17141_ _20109_/Q _17666_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20109_/D sky130_fd_sc_hd__mux2_1
X_11565_ _11872_/A _12006_/S _11564_/X _12012_/S vssd1 vssd1 vccd1 vccd1 _11565_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_155_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _13303_/A _13303_/B _13303_/C vssd1 vssd1 vccd1 vccd1 _13304_/Y sky130_fd_sc_hd__a21oi_1
X_10516_ _10512_/X _10515_/X _10516_/S vssd1 vssd1 vccd1 vccd1 _10516_/X sky130_fd_sc_hd__mux2_1
X_17072_ _20044_/Q _17874_/A1 _17076_/S vssd1 vssd1 vccd1 vccd1 _20044_/D sky130_fd_sc_hd__mux2_1
X_14284_ _14281_/B _14283_/Y _14417_/S vssd1 vssd1 vccd1 vccd1 _14284_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11496_ _11497_/B vssd1 vssd1 vccd1 vccd1 _11496_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13235_ _13002_/A _13233_/X _13234_/Y _13232_/X vssd1 vssd1 vccd1 vccd1 _13239_/B
+ sky130_fd_sc_hd__a31o_1
X_16023_ _16051_/A1 _16009_/X _16051_/B1 vssd1 vssd1 vccd1 vccd1 _16023_/Y sky130_fd_sc_hd__o21ai_1
X_10447_ _12072_/C1 _10435_/X _10438_/X _10446_/X vssd1 vssd1 vccd1 vccd1 _10447_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_226_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13166_ _13166_/A _13166_/B _13166_/C vssd1 vssd1 vccd1 vccd1 _13167_/B sky130_fd_sc_hd__and3_2
X_10378_ _10032_/Y _10377_/Y _09638_/Y vssd1 vssd1 vccd1 vccd1 _10378_/X sky130_fd_sc_hd__a21o_1
XFILLER_258_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_153_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20990_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12117_ _13432_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12117_/Y sky130_fd_sc_hd__nand2_1
XFILLER_285_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17974_ _20729_/Q _17976_/C _17974_/B1 vssd1 vssd1 vccd1 vccd1 _17975_/B sky130_fd_sc_hd__o21ai_1
X_13097_ _18667_/B _13097_/B vssd1 vssd1 vccd1 vccd1 _13097_/X sky130_fd_sc_hd__and2_1
XFILLER_78_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19713_ _20795_/CLK _19713_/D vssd1 vssd1 vccd1 vccd1 _19713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1740 _12304_/C1 vssd1 vssd1 vccd1 vccd1 _12371_/C1 sky130_fd_sc_hd__buf_6
X_16925_ input56/X input91/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16925_/X sky130_fd_sc_hd__mux2_8
X_12048_ _20487_/Q _20327_/Q _12053_/S vssd1 vssd1 vccd1 vccd1 _12048_/X sky130_fd_sc_hd__mux2_1
Xfanout1751 _10308_/S vssd1 vssd1 vccd1 vccd1 _12302_/S sky130_fd_sc_hd__buf_8
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1762 _12584_/A vssd1 vssd1 vccd1 vccd1 _18763_/A1 sky130_fd_sc_hd__buf_6
Xfanout1773 output482/A vssd1 vssd1 vccd1 vccd1 _13609_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19644_ _20075_/CLK _19644_/D vssd1 vssd1 vccd1 vccd1 _19644_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1784 _18313_/B vssd1 vssd1 vccd1 vccd1 _18299_/A1 sky130_fd_sc_hd__buf_12
Xfanout1795 _18209_/A1 vssd1 vssd1 vccd1 vccd1 _18199_/A1 sky130_fd_sc_hd__buf_6
X_16856_ _16884_/S _09526_/Y _16809_/X _16855_/Y vssd1 vssd1 vccd1 vccd1 _16856_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_281_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15807_ _15941_/B2 _15796_/X _15797_/X _15806_/X vssd1 vssd1 vccd1 vccd1 _15807_/X
+ sky130_fd_sc_hd__a22o_4
X_19575_ _20665_/CLK _19575_/D vssd1 vssd1 vccd1 vccd1 _19575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16787_ _19221_/Q _16996_/A2 _16713_/X _16784_/Y _16786_/X vssd1 vssd1 vccd1 vccd1
+ _16787_/X sky130_fd_sc_hd__o2111a_1
XFILLER_1_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13999_ _14035_/A1 _14011_/A2 _10550_/X _14038_/B1 _19848_/Q vssd1 vssd1 vccd1 vccd1
+ _14079_/C sky130_fd_sc_hd__o32a_2
XFILLER_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18526_ _18683_/B _18526_/B vssd1 vssd1 vccd1 vccd1 _18526_/X sky130_fd_sc_hd__or2_1
XFILLER_280_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15738_ _13416_/A _12565_/B _15737_/X vssd1 vssd1 vccd1 vccd1 _15738_/X sky130_fd_sc_hd__a21o_1
XFILLER_206_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _18320_/A _18457_/B _18457_/C vssd1 vssd1 vccd1 vccd1 _18457_/Y sky130_fd_sc_hd__nand3b_2
XFILLER_179_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15669_ _20803_/Q _15998_/A2 _15662_/X _14904_/X _15668_/X vssd1 vssd1 vccd1 vccd1
+ _15669_/X sky130_fd_sc_hd__a221o_1
XANTENNA_190 _19179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17408_ _17402_/Y _17407_/X _17406_/X _17432_/A vssd1 vssd1 vccd1 vccd1 _20251_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18388_ _20849_/Q _18387_/B _18387_/Y _18730_/A vssd1 vssd1 vccd1 vccd1 _20849_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17339_ _20218_/Q _17371_/A2 _17338_/X _18985_/A vssd1 vssd1 vccd1 vccd1 _20218_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20350_ _20685_/CLK _20350_/D vssd1 vssd1 vccd1 vccd1 _20350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19009_ _21024_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _19009_/X sky130_fd_sc_hd__or2_1
XFILLER_146_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20281_ _21024_/CLK _20281_/D vssd1 vssd1 vccd1 vccd1 _20281_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09526_ input47/X vssd1 vssd1 vccd1 vccd1 _09526_/Y sky130_fd_sc_hd__inv_2
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20617_ _20685_/CLK _20617_/D vssd1 vssd1 vccd1 vccd1 _20617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11350_ _20533_/Q _12300_/S vssd1 vssd1 vccd1 vccd1 _11350_/X sky130_fd_sc_hd__or2_1
XFILLER_165_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20548_ _20717_/CLK _20548_/D vssd1 vssd1 vccd1 vccd1 _20548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _12519_/C _10298_/X _10300_/X vssd1 vssd1 vccd1 vccd1 _10301_/X sky130_fd_sc_hd__a21o_1
XFILLER_192_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11281_ _11281_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11281_/Y sky130_fd_sc_hd__nand2_1
XFILLER_180_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20479_ _20479_/CLK _20479_/D vssd1 vssd1 vccd1 vccd1 _20479_/Q sky130_fd_sc_hd__dfxtp_1
X_13020_ _20969_/Q _20903_/Q vssd1 vssd1 vccd1 vccd1 _13258_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10232_ _11008_/A3 _10231_/X _10228_/X _11275_/A vssd1 vssd1 vccd1 vccd1 _10232_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_279_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1003 _15019_/A vssd1 vssd1 vccd1 vccd1 _15021_/A sky130_fd_sc_hd__clkbuf_16
X_10163_ _12245_/A1 _17899_/A1 _10162_/X vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1014 _15185_/B vssd1 vssd1 vccd1 vccd1 _15494_/B sky130_fd_sc_hd__buf_6
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1025 _16963_/A2 vssd1 vssd1 vccd1 vccd1 _16979_/A2 sky130_fd_sc_hd__buf_4
Xfanout1036 _17886_/A1 vssd1 vssd1 vccd1 vccd1 _17920_/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout1047 _11063_/X vssd1 vssd1 vccd1 vccd1 _17782_/A1 sky130_fd_sc_hd__buf_8
XFILLER_0_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14971_ _14971_/A _14971_/B _14971_/C vssd1 vssd1 vccd1 vccd1 _14972_/C sky130_fd_sc_hd__or3_1
XFILLER_121_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10094_ _10090_/X _10093_/X _10516_/S vssd1 vssd1 vccd1 vccd1 _10094_/X sky130_fd_sc_hd__mux2_1
Xfanout1058 _17891_/A1 vssd1 vssd1 vccd1 vccd1 _17857_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1069 _09748_/Y vssd1 vssd1 vccd1 vccd1 _12107_/A1 sky130_fd_sc_hd__buf_4
X_16710_ _16710_/A _16710_/B vssd1 vssd1 vccd1 vccd1 _16714_/D sky130_fd_sc_hd__or2_1
XFILLER_275_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13922_ _19126_/Q _13921_/B _13921_/Y _14758_/C1 vssd1 vssd1 vccd1 vccd1 _19126_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_248_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17690_ _20474_/Q _17933_/A1 _17706_/S vssd1 vssd1 vccd1 vccd1 _20474_/D sky130_fd_sc_hd__mux2_1
XFILLER_19_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16641_ _19898_/Q _17051_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19898_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13853_ _19661_/Q _13853_/B vssd1 vssd1 vccd1 vccd1 _13853_/Y sky130_fd_sc_hd__nand2_8
XFILLER_263_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12804_ _19516_/Q _12804_/B vssd1 vssd1 vccd1 vccd1 _12804_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19360_ _20715_/CLK _19360_/D vssd1 vssd1 vccd1 vccd1 _19360_/Q sky130_fd_sc_hd__dfxtp_1
X_16572_ _19852_/Q _16576_/A2 _16576_/B1 input23/X vssd1 vssd1 vccd1 vccd1 _16573_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10996_ _11268_/A _20592_/Q _11261_/C vssd1 vssd1 vccd1 vccd1 _10996_/X sky130_fd_sc_hd__and3_1
XFILLER_16_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13784_ _16240_/A1 _13537_/Y _13539_/Y split3/X vssd1 vssd1 vccd1 vccd1 _13784_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_215_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18311_ _20816_/Q _18310_/Y _18311_/S vssd1 vssd1 vccd1 vccd1 _18312_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _12468_/B _16063_/A2 _15522_/X vssd1 vssd1 vccd1 vccd1 _15524_/B sky130_fd_sc_hd__a21oi_1
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19291_ _20681_/CLK _19291_/D vssd1 vssd1 vccd1 vccd1 _19291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12735_ _12736_/B _12736_/C _12736_/A vssd1 vssd1 vccd1 vccd1 _13281_/A sky130_fd_sc_hd__a21o_2
XFILLER_204_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18242_ _18718_/A _18242_/B vssd1 vssd1 vccd1 vccd1 _20802_/D sky130_fd_sc_hd__and2_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15454_ _19712_/Q _15453_/X _15454_/S vssd1 vssd1 vccd1 vccd1 _15454_/X sky130_fd_sc_hd__mux2_2
XFILLER_188_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12666_ _12666_/A vssd1 vssd1 vccd1 vccd1 _12666_/Y sky130_fd_sc_hd__inv_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14405_ _14405_/A _14405_/B vssd1 vssd1 vccd1 vccd1 _14405_/X sky130_fd_sc_hd__xor2_1
X_11617_ _19681_/Q _12013_/S _11616_/X _12003_/C vssd1 vssd1 vccd1 vccd1 _11617_/X
+ sky130_fd_sc_hd__o211a_1
X_18173_ _19530_/Q _18198_/B vssd1 vssd1 vccd1 vccd1 _18173_/Y sky130_fd_sc_hd__nand2b_2
X_15385_ _21020_/Q _20988_/Q _15508_/S vssd1 vssd1 vccd1 vccd1 _15385_/X sky130_fd_sc_hd__mux2_1
X_12597_ _19497_/Q _12665_/A vssd1 vssd1 vccd1 vccd1 _12680_/B sky130_fd_sc_hd__and2_2
XFILLER_156_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17124_ _20092_/Q _17926_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20092_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11548_ _11546_/X _11547_/X _11563_/S vssd1 vssd1 vccd1 vccd1 _11548_/X sky130_fd_sc_hd__mux2_1
X_14336_ _14427_/A _14332_/B _14335_/X vssd1 vssd1 vccd1 vccd1 _14336_/X sky130_fd_sc_hd__a21bo_1
XFILLER_237_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17055_ _20027_/Q _17751_/A1 _17080_/S vssd1 vssd1 vccd1 vccd1 _20027_/D sky130_fd_sc_hd__mux2_1
XFILLER_274_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14267_ _20281_/Q _14267_/A2 _14267_/B1 input221/X vssd1 vssd1 vccd1 vccd1 _14269_/B
+ sky130_fd_sc_hd__a22o_4
X_11479_ _20642_/Q _20606_/Q _12182_/S vssd1 vssd1 vccd1 vccd1 _11479_/X sky130_fd_sc_hd__mux2_1
X_13218_ _13373_/A _13218_/B _13218_/C vssd1 vssd1 vccd1 vccd1 _13218_/Y sky130_fd_sc_hd__nand3_1
X_16006_ _19179_/Q _16063_/A2 _15981_/A _16034_/S vssd1 vssd1 vccd1 vccd1 _16007_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_171_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14198_ _19502_/Q _14198_/B vssd1 vssd1 vccd1 vccd1 _14199_/B sky130_fd_sc_hd__nand2_2
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13149_ _15264_/A _13538_/B _10798_/X _10885_/A vssd1 vssd1 vccd1 vccd1 _13150_/B
+ sky130_fd_sc_hd__a211o_2
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _18054_/A _17962_/C vssd1 vssd1 vccd1 vccd1 _17957_/Y sky130_fd_sc_hd__nor2_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1570 _09625_/Y vssd1 vssd1 vccd1 vccd1 _12392_/C1 sky130_fd_sc_hd__buf_4
XFILLER_226_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16908_ _16932_/A1 _16907_/X _16932_/B1 vssd1 vssd1 vccd1 vccd1 _16908_/Y sky130_fd_sc_hd__o21ai_2
Xfanout1581 _11353_/C1 vssd1 vssd1 vccd1 vccd1 _12398_/C1 sky130_fd_sc_hd__buf_6
XFILLER_238_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17888_ _20659_/Q _17888_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20659_/D sky130_fd_sc_hd__mux2_1
Xfanout1592 _11363_/A1 vssd1 vssd1 vccd1 vccd1 _12399_/A1 sky130_fd_sc_hd__buf_6
XFILLER_266_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19627_ _20667_/CLK _19627_/D vssd1 vssd1 vccd1 vccd1 _19627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16839_ _16932_/B1 _16836_/X _16838_/X _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16840_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_254_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19558_ _19617_/CLK _19558_/D vssd1 vssd1 vccd1 vccd1 _19558_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20719_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18509_ _20896_/Q _18474_/S _18508_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18510_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_202_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19489_ _20580_/CLK _19489_/D vssd1 vssd1 vccd1 vccd1 _19489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20402_ _20759_/CLK _20402_/D vssd1 vssd1 vccd1 vccd1 _20402_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20333_ _20667_/CLK _20333_/D vssd1 vssd1 vccd1 vccd1 _20333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20264_ _20421_/CLK _20264_/D vssd1 vssd1 vccd1 vccd1 _20264_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20195_ _20688_/CLK _20195_/D vssd1 vssd1 vccd1 vccd1 _20195_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput106 dout0[9] vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput117 dout1[19] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput128 dout1[29] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput139 dout1[39] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__clkbuf_2
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _11368_/A1 _13653_/B _10849_/X _11189_/B vssd1 vssd1 vccd1 vccd1 _10884_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _12510_/A vssd1 vssd1 vccd1 vccd1 _14894_/A sky130_fd_sc_hd__inv_8
X_10781_ _12265_/A _10781_/B vssd1 vssd1 vccd1 vccd1 _10781_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ _18765_/C _12588_/C _12520_/C _12520_/D vssd1 vssd1 vccd1 vccd1 _12982_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_213_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12450_/A _12445_/B _16054_/A vssd1 vssd1 vccd1 vccd1 _12451_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11402_ _11774_/B vssd1 vssd1 vccd1 vccd1 _13570_/A sky130_fd_sc_hd__inv_2
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15170_ _15170_/A _15170_/B vssd1 vssd1 vccd1 vccd1 _15170_/X sky130_fd_sc_hd__or2_1
X_12382_ _12380_/X _12381_/X _12391_/S vssd1 vssd1 vccd1 vccd1 _12383_/B sky130_fd_sc_hd__mux2_1
XFILLER_193_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_90 _11806_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ _14121_/A _16710_/B vssd1 vssd1 vccd1 vccd1 _14121_/X sky130_fd_sc_hd__or2_4
XFILLER_165_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11333_ _20373_/Q _20437_/Q _12375_/S vssd1 vssd1 vccd1 vccd1 _11333_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14052_ _19185_/Q _14082_/A2 _14051_/X _16097_/B1 vssd1 vssd1 vccd1 vccd1 _19185_/D
+ sky130_fd_sc_hd__o211a_1
X_11264_ _20397_/Q _09689_/D _11262_/X _11263_/X vssd1 vssd1 vccd1 vccd1 _11264_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13003_ _20945_/Q _13363_/B _18667_/B vssd1 vssd1 vccd1 vccd1 _13003_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_234_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10215_ _19677_/Q _20165_/Q _10217_/S vssd1 vssd1 vccd1 vccd1 _10215_/X sky130_fd_sc_hd__mux2_1
XFILLER_268_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18860_ _18620_/Y _18867_/A2 _18858_/Y _18859_/Y vssd1 vssd1 vccd1 vccd1 _18860_/X
+ sky130_fd_sc_hd__a22o_1
X_11195_ _12332_/A _20494_/Q _12339_/S0 _20526_/Q vssd1 vssd1 vccd1 vccd1 _11195_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17811_ _20588_/Q _17951_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20588_/D sky130_fd_sc_hd__mux2_1
XFILLER_267_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10146_ _20538_/Q _10924_/S vssd1 vssd1 vccd1 vccd1 _10146_/X sky130_fd_sc_hd__or2_1
XFILLER_79_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ _09494_/Y _18790_/X _18830_/A vssd1 vssd1 vccd1 vccd1 _18791_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17742_ _20523_/Q _17916_/A1 _17742_/S vssd1 vssd1 vccd1 vccd1 _20523_/D sky130_fd_sc_hd__mux2_1
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14954_ _15308_/B _15308_/C vssd1 vssd1 vccd1 vccd1 _14954_/X sky130_fd_sc_hd__and2_1
X_10077_ _11367_/B _13684_/A vssd1 vssd1 vccd1 vccd1 _10077_/Y sky130_fd_sc_hd__nand2_1
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _19118_/Q _13906_/B _13932_/B1 _13479_/A vssd1 vssd1 vccd1 vccd1 _19118_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_130_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17673_ _20459_/Q _17707_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20459_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14885_ _15577_/S _14885_/B vssd1 vssd1 vccd1 vccd1 _14885_/X sky130_fd_sc_hd__or2_4
XFILLER_223_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19412_ _20701_/CLK _19412_/D vssd1 vssd1 vccd1 vccd1 _19412_/Q sky130_fd_sc_hd__dfxtp_1
X_16624_ _19883_/Q _17938_/A1 _16632_/S vssd1 vssd1 vccd1 vccd1 _19883_/D sky130_fd_sc_hd__mux2_1
X_13836_ _20264_/Q _20265_/Q vssd1 vssd1 vccd1 vccd1 _17457_/B sky130_fd_sc_hd__and2b_4
XFILLER_189_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _20698_/CLK _19343_/D vssd1 vssd1 vccd1 vccd1 _19343_/Q sky130_fd_sc_hd__dfxtp_1
X_16555_ _16557_/A _16555_/B vssd1 vssd1 vccd1 vccd1 _19843_/D sky130_fd_sc_hd__or2_1
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10979_ _11268_/A _20304_/Q _10979_/C vssd1 vssd1 vccd1 vccd1 _10979_/X sky130_fd_sc_hd__and3_1
XFILLER_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13767_ _13777_/A _13767_/B vssd1 vssd1 vccd1 vccd1 _13767_/X sky130_fd_sc_hd__or2_1
XFILLER_204_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15506_ _19714_/Q _15595_/A2 _15595_/B1 _19746_/Q vssd1 vssd1 vccd1 vccd1 _15506_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19274_ _20467_/CLK _19274_/D vssd1 vssd1 vccd1 vccd1 _19274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12718_ _12718_/A _12718_/B vssd1 vssd1 vccd1 vccd1 _12718_/X sky130_fd_sc_hd__or2_1
X_16486_ _19795_/Q _17706_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19795_/D sky130_fd_sc_hd__mux2_1
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13698_ _13698_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13698_/X sky130_fd_sc_hd__or2_4
X_18225_ _18505_/B vssd1 vssd1 vccd1 vccd1 _18225_/Y sky130_fd_sc_hd__inv_4
XFILLER_248_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15437_ _15468_/A _15437_/B vssd1 vssd1 vccd1 vccd1 _15437_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12649_ _15267_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _12649_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18156_ _18389_/A _18156_/B _18156_/C _18318_/A vssd1 vssd1 vccd1 vccd1 _18157_/D
+ sky130_fd_sc_hd__or4b_2
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15368_ _19534_/Q _15492_/A _15367_/Y _16179_/A vssd1 vssd1 vccd1 vccd1 _19534_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17107_ _20077_/Q _17107_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20077_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ _19234_/Q _14398_/A2 _14318_/X _14776_/C1 vssd1 vssd1 vccd1 vccd1 _19234_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18087_ _20770_/Q _18087_/B vssd1 vssd1 vccd1 vccd1 _18093_/C sky130_fd_sc_hd__and2_2
XFILLER_172_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15299_ _15468_/A _15294_/X _15297_/Y _14870_/S _15298_/X vssd1 vssd1 vccd1 vccd1
+ _15299_/X sky130_fd_sc_hd__a221o_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17038_ _20016_/Q _12928_/A _17038_/S vssd1 vssd1 vccd1 vccd1 _20016_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09860_ _09861_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__or2_2
Xfanout807 _13184_/X vssd1 vssd1 vccd1 vccd1 _14525_/B sky130_fd_sc_hd__buf_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout818 _15633_/Y vssd1 vssd1 vccd1 vccd1 fanout818/X sky130_fd_sc_hd__buf_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout829 _13740_/A vssd1 vssd1 vccd1 vccd1 _13735_/A sky130_fd_sc_hd__buf_2
XFILLER_140_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09791_ _20483_/Q _20323_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _09791_/X sky130_fd_sc_hd__mux2_1
XFILLER_274_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18989_ _21014_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _18989_/X sky130_fd_sc_hd__or2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20951_ _21017_/CLK _20951_/D vssd1 vssd1 vccd1 vccd1 _20951_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20882_ _20980_/CLK _20882_/D vssd1 vssd1 vccd1 vccd1 _20882_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20316_ _20702_/CLK _20316_/D vssd1 vssd1 vccd1 vccd1 _20316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20247_ _20296_/CLK _20247_/D vssd1 vssd1 vccd1 vccd1 _20247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ _20481_/Q _11616_/B _11948_/A1 vssd1 vssd1 vccd1 vccd1 _10000_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20178_ _20641_/CLK _20178_/D vssd1 vssd1 vccd1 vccd1 _20178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09989_ _09987_/X _09988_/X _12006_/S vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _11942_/X _11950_/Y _12192_/A1 _11934_/X vssd1 vssd1 vccd1 vccd1 _11951_/X
+ sky130_fd_sc_hd__o2bb2a_2
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10902_ _11268_/A _20058_/Q _11261_/C vssd1 vssd1 vccd1 vccd1 _10902_/X sky130_fd_sc_hd__and3_1
XFILLER_45_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14670_ _16605_/A _17574_/B _14670_/C vssd1 vssd1 vccd1 vccd1 _14670_/X sky130_fd_sc_hd__and3_4
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11882_ _13418_/A _11882_/B vssd1 vssd1 vccd1 vccd1 _11882_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_232_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10833_ _12230_/A1 _20498_/Q _12309_/S _10823_/X vssd1 vssd1 vccd1 vccd1 _10833_/X
+ sky130_fd_sc_hd__o211a_1
X_13621_ _13626_/A1 _13361_/C _13427_/A _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13621_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16340_ _19723_/Q _16340_/B vssd1 vssd1 vccd1 vccd1 _16346_/C sky130_fd_sc_hd__and2_2
X_10764_ _11367_/B _13657_/B vssd1 vssd1 vccd1 vccd1 _10764_/Y sky130_fd_sc_hd__nand2_1
X_13552_ _13552_/A _13552_/B _13552_/C vssd1 vssd1 vccd1 vccd1 _14184_/A sky130_fd_sc_hd__and3_2
XFILLER_34_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ _12510_/A _14808_/A _12510_/C _15095_/B vssd1 vssd1 vccd1 vccd1 _18765_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13483_ _12675_/A _12675_/C _12675_/B vssd1 vssd1 vccd1 vccd1 _13483_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16271_ _19687_/Q _17805_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19687_/D sky130_fd_sc_hd__mux2_1
X_10695_ _10693_/X _10694_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _10695_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18010_ _20741_/Q _18011_/C _20742_/Q vssd1 vssd1 vccd1 vccd1 _18012_/B sky130_fd_sc_hd__a21oi_1
XFILLER_201_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15222_ _13524_/A _15259_/B _15220_/X _15221_/Y vssd1 vssd1 vccd1 vccd1 _15222_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12434_ _19524_/Q _16009_/A _15895_/S vssd1 vssd1 vccd1 vccd1 _12443_/B sky130_fd_sc_hd__mux2_8
XFILLER_201_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12365_ _19557_/Q _12365_/A2 _11225_/B _19621_/Q vssd1 vssd1 vccd1 vccd1 _12365_/X
+ sky130_fd_sc_hd__a22o_1
X_15153_ _11103_/Y _15152_/X _15492_/A vssd1 vssd1 vccd1 vccd1 _15153_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14104_ _19211_/Q _14104_/A2 _14103_/X _14104_/C1 vssd1 vssd1 vccd1 vccd1 _19211_/D
+ sky130_fd_sc_hd__o211a_1
X_11316_ _15075_/A _15075_/B _11223_/A _11223_/B vssd1 vssd1 vccd1 vccd1 _11781_/B
+ sky130_fd_sc_hd__a2bb2o_4
X_15084_ _20915_/Q _15337_/A2 _15083_/X vssd1 vssd1 vccd1 vccd1 _15084_/X sky130_fd_sc_hd__o21a_1
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19961_ _20621_/CLK _19961_/D vssd1 vssd1 vccd1 vccd1 _19961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12296_ _19429_/Q _20588_/Q _12296_/S vssd1 vssd1 vccd1 vccd1 _12296_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14035_ _14035_/A1 _14041_/A2 _10121_/X _14035_/B1 _19860_/Q vssd1 vssd1 vccd1 vccd1
+ _14103_/C sky130_fd_sc_hd__o32a_1
X_18912_ _18973_/A _18912_/B vssd1 vssd1 vccd1 vccd1 _21001_/D sky130_fd_sc_hd__nor2_1
X_11247_ _09595_/Y _11237_/X _11246_/Y _11235_/A vssd1 vssd1 vccd1 vccd1 _11247_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_141_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19892_ _20580_/CLK _19892_/D vssd1 vssd1 vccd1 vccd1 _19892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18843_ _19096_/Q _18864_/A2 _18864_/B1 _15494_/A vssd1 vssd1 vccd1 vccd1 _18844_/B
+ sky130_fd_sc_hd__a22o_1
X_11178_ _20558_/Q _10924_/S _11177_/X vssd1 vssd1 vccd1 vccd1 _11178_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10129_ _19411_/Q _20570_/Q _10217_/S vssd1 vssd1 vccd1 vccd1 _10129_/X sky130_fd_sc_hd__mux2_1
X_18774_ _19117_/Q _18773_/X _18901_/S vssd1 vssd1 vccd1 vccd1 _18774_/Y sky130_fd_sc_hd__o21ai_1
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ _16053_/A _15123_/X _15983_/Y _15985_/Y vssd1 vssd1 vccd1 vccd1 _15986_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17725_ _20506_/Q _17899_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20506_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14937_ _15019_/A _15014_/B _15133_/B vssd1 vssd1 vccd1 vccd1 _14967_/A sky130_fd_sc_hd__and3_1
XFILLER_270_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ _20442_/Q _17933_/A1 _17657_/S vssd1 vssd1 vccd1 vccd1 _20442_/D sky130_fd_sc_hd__mux2_1
X_14868_ _15039_/B _14867_/X _15062_/S vssd1 vssd1 vccd1 vccd1 _14868_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16607_ _19866_/Q _17921_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19866_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13819_ _13822_/A1 _13765_/B split9/X input235/X vssd1 vssd1 vccd1 vccd1 _13819_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17587_ _20345_/Q _17898_/A1 _17601_/S vssd1 vssd1 vccd1 vccd1 _20345_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14799_ _19524_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14799_/X sky130_fd_sc_hd__or2_1
XFILLER_259_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19326_ _20649_/CLK _19326_/D vssd1 vssd1 vccd1 vccd1 _19326_/Q sky130_fd_sc_hd__dfxtp_1
X_16538_ _19835_/Q _16592_/A2 _16592_/B1 input36/X vssd1 vssd1 vccd1 vccd1 _16539_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19257_ _21013_/CLK _19257_/D vssd1 vssd1 vccd1 vccd1 _19257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16469_ _19778_/Q _17689_/A1 _16483_/S vssd1 vssd1 vccd1 vccd1 _19778_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18208_ _19537_/Q _18213_/B vssd1 vssd1 vccd1 vccd1 _18208_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_148_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19188_ _20273_/CLK _19188_/D vssd1 vssd1 vccd1 vccd1 _19188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18139_ _18323_/B _18139_/B vssd1 vssd1 vccd1 vccd1 _18981_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20101_ _20557_/CLK _20101_/D vssd1 vssd1 vccd1 vccd1 _20101_/Q sky130_fd_sc_hd__dfxtp_1
X_09912_ _09910_/X _09911_/X _11849_/S vssd1 vssd1 vccd1 vccd1 _09912_/X sky130_fd_sc_hd__mux2_1
XFILLER_259_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout604 _14601_/X vssd1 vssd1 vccd1 vccd1 _14628_/S sky130_fd_sc_hd__buf_6
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout615 _14488_/X vssd1 vssd1 vccd1 vccd1 _14517_/S sky130_fd_sc_hd__buf_12
Xfanout626 _14043_/B1 vssd1 vssd1 vccd1 vccd1 _14034_/B1 sky130_fd_sc_hd__buf_2
XFILLER_98_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20032_ _20657_/CLK _20032_/D vssd1 vssd1 vccd1 vccd1 _20032_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout637 _16707_/X vssd1 vssd1 vccd1 vccd1 _17011_/B1 sky130_fd_sc_hd__buf_12
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09843_ _19420_/Q _20579_/Q _10397_/S vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__mux2_1
Xfanout648 _16077_/B vssd1 vssd1 vccd1 vccd1 _16127_/A2 sky130_fd_sc_hd__buf_4
XFILLER_58_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout659 _14737_/X vssd1 vssd1 vccd1 vccd1 _14797_/B sky130_fd_sc_hd__buf_2
XFILLER_258_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09774_ _19421_/Q _20580_/Q _12013_/S vssd1 vssd1 vccd1 vccd1 _09774_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20934_ _21008_/CLK _20934_/D vssd1 vssd1 vccd1 vccd1 _20934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20865_ _21020_/CLK _20865_/D vssd1 vssd1 vccd1 vccd1 _20865_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20796_ _20796_/CLK _20796_/D vssd1 vssd1 vccd1 vccd1 _20796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10480_ _11273_/A1 _19344_/Q _20699_/Q _10485_/S _12519_/C vssd1 vssd1 vccd1 vccd1
+ _10480_/X sky130_fd_sc_hd__a221o_1
XFILLER_194_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12150_ _12148_/X _12149_/X _12150_/S vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11101_ _11101_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11101_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ _19649_/Q _19955_/Q _19293_/Q _20080_/Q _12081_/S0 _12084_/C vssd1 vssd1
+ vccd1 vccd1 _12081_/X sky130_fd_sc_hd__mux4_1
XFILLER_118_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ _20464_/Q _20304_/Q _11039_/S vssd1 vssd1 vccd1 vccd1 _11032_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _12513_/D _15978_/A2 _15816_/A _16063_/B2 vssd1 vssd1 vccd1 vccd1 _15841_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _20743_/Q _15934_/A2 _15934_/B1 _20775_/Q vssd1 vssd1 vccd1 vccd1 _15771_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_252_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12983_ _19218_/Q _13498_/B vssd1 vssd1 vccd1 vccd1 _13499_/A sky130_fd_sc_hd__and2_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _20290_/Q _17524_/B vssd1 vssd1 vccd1 vccd1 _17510_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14722_ _19479_/Q _17937_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19479_/D sky130_fd_sc_hd__mux2_1
XFILLER_245_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18490_ _18490_/A _18490_/B vssd1 vssd1 vccd1 vccd1 _18490_/X sky130_fd_sc_hd__or2_4
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _11928_/X _11933_/X _12012_/S vssd1 vssd1 vccd1 vccd1 _11934_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_520 _13828_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_531 _14069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17441_ _17441_/A _17451_/A _17441_/C vssd1 vssd1 vccd1 vccd1 _17443_/C sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_178_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19246_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_542 _11897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14653_ _19415_/Q _17937_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19415_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_553 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_564 _11199_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11865_ _19889_/Q _19790_/Q _11947_/S vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__mux2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_575 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_107_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20766_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_260_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_586 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13604_ _13043_/Y _13604_/B vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__nand2b_1
X_10816_ _19870_/Q _19771_/Q _12389_/S vssd1 vssd1 vccd1 vccd1 _10816_/X sky130_fd_sc_hd__mux2_1
XFILLER_214_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_597 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17372_ _20234_/Q _17378_/A2 _17382_/B1 _20283_/Q _17380_/C1 vssd1 vssd1 vccd1 vccd1
+ _17372_/X sky130_fd_sc_hd__a221o_1
X_14584_ _19350_/Q _17936_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19350_/D sky130_fd_sc_hd__mux2_1
X_11796_ _13423_/A _11796_/B vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__xnor2_2
XFILLER_41_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19111_ _20273_/CLK _19111_/D vssd1 vssd1 vccd1 vccd1 _19111_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_213_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16323_ _18086_/A _16323_/B _16324_/B vssd1 vssd1 vccd1 vccd1 _19716_/D sky130_fd_sc_hd__nor3_1
X_13535_ _18462_/A _13534_/X _13531_/X _13552_/A vssd1 vssd1 vccd1 vccd1 _14173_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ _12312_/A1 _20499_/Q _12309_/S _10739_/X vssd1 vssd1 vccd1 vccd1 _10747_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19042_ _18300_/Y _19046_/A2 _19048_/B1 _12550_/B _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19042_/X sky130_fd_sc_hd__a221o_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16254_ _19670_/Q _17788_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19670_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ _12392_/C1 _10667_/X _10670_/X _10677_/X _12400_/A1 vssd1 vssd1 vccd1 vccd1
+ _10678_/X sky130_fd_sc_hd__a311o_1
XFILLER_199_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13466_ _13466_/A _13466_/B vssd1 vssd1 vccd1 vccd1 _13466_/X sky130_fd_sc_hd__or2_2
XFILLER_173_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15205_ _15026_/Y _15188_/X _15673_/B1 vssd1 vssd1 vccd1 vccd1 _15206_/C sky130_fd_sc_hd__o21a_1
X_12417_ _19895_/Q _19796_/Q _12417_/S vssd1 vssd1 vccd1 vccd1 _12417_/X sky130_fd_sc_hd__mux2_1
X_16185_ _16185_/A _16185_/B vssd1 vssd1 vccd1 vccd1 _19616_/D sky130_fd_sc_hd__and2_1
X_13397_ _20968_/Q _13397_/B vssd1 vssd1 vccd1 vccd1 _13397_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15136_ _20916_/Q _15567_/A2 _15388_/S vssd1 vssd1 vccd1 vccd1 _15136_/X sky130_fd_sc_hd__o21ba_1
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12348_ _12357_/A1 _12346_/X _12347_/X vssd1 vssd1 vccd1 vccd1 _12348_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19944_ _20660_/CLK _19944_/D vssd1 vssd1 vccd1 vccd1 _19944_/Q sky130_fd_sc_hd__dfxtp_1
X_15067_ _14838_/X _14885_/B _15067_/S vssd1 vssd1 vccd1 vccd1 _15067_/X sky130_fd_sc_hd__mux2_1
X_12279_ _12282_/B vssd1 vssd1 vccd1 vccd1 _12279_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _19205_/Q _14091_/C _14039_/S vssd1 vssd1 vccd1 vccd1 _14018_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19875_ _21047_/A _19875_/D vssd1 vssd1 vccd1 vccd1 _19875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18826_ _20989_/Q _18861_/B vssd1 vssd1 vccd1 vccd1 _18826_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18757_ _13552_/A _13107_/B _18470_/Y _18756_/B vssd1 vssd1 vccd1 vccd1 _18757_/X
+ sky130_fd_sc_hd__a22o_1
X_15969_ _16017_/C1 _15968_/X _15964_/X vssd1 vssd1 vccd1 vccd1 _15969_/X sky130_fd_sc_hd__o21a_4
XFILLER_64_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17708_ _20492_/Q _17708_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20492_/D sky130_fd_sc_hd__mux2_1
XFILLER_237_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09490_ _19146_/Q vssd1 vssd1 vccd1 vccd1 _09490_/Y sky130_fd_sc_hd__inv_2
X_18688_ _18560_/X _18688_/A2 _18686_/Y _18687_/Y vssd1 vssd1 vccd1 vccd1 _18689_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17639_ _20395_/Q _17707_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20395_/D sky130_fd_sc_hd__mux2_1
XFILLER_252_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20650_ _20682_/CLK _20650_/D vssd1 vssd1 vccd1 vccd1 _20650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19309_ _20467_/CLK _19309_/D vssd1 vssd1 vccd1 vccd1 _19309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20581_ _20713_/CLK _20581_/D vssd1 vssd1 vccd1 vccd1 _20581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20015_ _20017_/CLK _20015_/D vssd1 vssd1 vccd1 vccd1 _20015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09826_ _11922_/A1 _13730_/A _12158_/B1 vssd1 vssd1 vccd1 vccd1 _09826_/X sky130_fd_sc_hd__o21a_1
XFILLER_247_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout489 _17919_/X vssd1 vssd1 vccd1 vccd1 _17946_/S sky130_fd_sc_hd__buf_6
XFILLER_274_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09757_ _12003_/A _20680_/Q _12008_/C vssd1 vssd1 vccd1 vccd1 _09757_/X sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20480_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_261_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09688_/A _09688_/B vssd1 vssd1 vccd1 vccd1 _09688_/Y sky130_fd_sc_hd__nand2_2
XFILLER_243_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20917_ _21015_/CLK _20917_/D vssd1 vssd1 vccd1 vccd1 _20917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_200_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20678_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_270_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11651_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _13167_/A sky130_fd_sc_hd__and2_2
XFILLER_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20848_ _21000_/CLK _20848_/D vssd1 vssd1 vccd1 vccd1 _20848_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10601_ _19276_/Q _11693_/B _12190_/C1 vssd1 vssd1 vccd1 vccd1 _10601_/X sky130_fd_sc_hd__a21o_1
XFILLER_168_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11581_ _20576_/Q _12044_/B _11580_/X _12123_/C1 vssd1 vssd1 vccd1 vccd1 _11581_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20779_ _20812_/CLK _20779_/D vssd1 vssd1 vccd1 vccd1 _20779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ _11290_/A _20667_/Q _11026_/C vssd1 vssd1 vccd1 vccd1 _10532_/X sky130_fd_sc_hd__or3_1
X_13320_ _14275_/A1 _19227_/Q _18352_/C1 _13319_/Y vssd1 vssd1 vccd1 vccd1 _13361_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10463_ _11239_/A1 _09670_/Y _10462_/X _11239_/B1 _19849_/Q vssd1 vssd1 vccd1 vccd1
+ _10463_/X sky130_fd_sc_hd__o32a_1
X_13251_ _13264_/A _13264_/C vssd1 vssd1 vccd1 vccd1 _13389_/C sky130_fd_sc_hd__nor2_2
XFILLER_171_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12202_ _12202_/A _12202_/B _13183_/A vssd1 vssd1 vccd1 vccd1 _12203_/B sky130_fd_sc_hd__nand3_1
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13182_ _13182_/A _13182_/B vssd1 vssd1 vccd1 vccd1 _15981_/A sky130_fd_sc_hd__xnor2_4
X_10394_ _10391_/X _10393_/X _18765_/B vssd1 vssd1 vccd1 vccd1 _10394_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12133_ _20393_/Q _20457_/Q _12133_/S vssd1 vssd1 vccd1 vccd1 _12133_/X sky130_fd_sc_hd__mux2_1
X_17990_ _20734_/Q _17991_/C _17989_/Y vssd1 vssd1 vccd1 vccd1 _20734_/D sky130_fd_sc_hd__o21a_1
XFILLER_151_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16941_ input58/X input93/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16941_/X sky130_fd_sc_hd__mux2_8
XFILLER_150_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1900 fanout1905/X vssd1 vssd1 vccd1 vccd1 _14780_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12064_ _19392_/Q _20683_/Q _12064_/S vssd1 vssd1 vccd1 vccd1 _12064_/X sky130_fd_sc_hd__mux2_1
Xfanout1911 _18724_/A vssd1 vssd1 vccd1 vccd1 _18728_/A sky130_fd_sc_hd__buf_4
Xfanout1922 _14070_/C1 vssd1 vssd1 vccd1 vccd1 _15288_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1933 _14185_/C1 vssd1 vssd1 vccd1 vccd1 _18702_/A sky130_fd_sc_hd__clkbuf_4
X_11015_ _09569_/A _13648_/B _11014_/X vssd1 vssd1 vccd1 vccd1 _11015_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_78_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1944 _17963_/B1 vssd1 vssd1 vccd1 vccd1 _16129_/B1 sky130_fd_sc_hd__buf_4
X_19660_ _21044_/CLK _19660_/D vssd1 vssd1 vccd1 vccd1 _19660_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1955 _18422_/A vssd1 vssd1 vccd1 vccd1 _18708_/A sky130_fd_sc_hd__clkbuf_4
X_16872_ _16805_/X _16869_/Y _16871_/X _17008_/A1 vssd1 vssd1 vccd1 vccd1 _16872_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_277_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1966 _18112_/A vssd1 vssd1 vccd1 vccd1 _18980_/A sky130_fd_sc_hd__buf_4
XFILLER_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1977 _18842_/A vssd1 vssd1 vccd1 vccd1 _18835_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_238_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18611_ _20926_/Q _18619_/B vssd1 vssd1 vccd1 vccd1 _18611_/Y sky130_fd_sc_hd__nand2_1
Xfanout990 _10045_/X vssd1 vssd1 vccd1 vccd1 _17898_/A1 sky130_fd_sc_hd__buf_4
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1988 _17952_/A vssd1 vssd1 vccd1 vccd1 _18808_/A sky130_fd_sc_hd__buf_4
X_15823_ _19725_/Q _15961_/A2 _15961_/B1 _19757_/Q vssd1 vssd1 vccd1 vccd1 _15823_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_253_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1999 _17998_/A vssd1 vssd1 vccd1 vccd1 _18094_/A sky130_fd_sc_hd__buf_4
X_19591_ _19606_/CLK _19591_/D vssd1 vssd1 vccd1 vccd1 _19591_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ _20907_/Q fanout750/X _18541_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18543_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15973_/A1 _15753_/X _15741_/X vssd1 vssd1 vccd1 vccd1 _15754_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12966_ _18198_/B _19301_/Q _12965_/X vssd1 vssd1 vccd1 vccd1 _14112_/C sky130_fd_sc_hd__nor3b_2
XFILLER_205_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _19462_/Q _17920_/A1 _14719_/S vssd1 vssd1 vccd1 vccd1 _19462_/D sky130_fd_sc_hd__mux2_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18473_ _18473_/A _18985_/B vssd1 vssd1 vccd1 vccd1 _18473_/Y sky130_fd_sc_hd__nand2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _11915_/X _11916_/X _11917_/S vssd1 vssd1 vccd1 vccd1 _11917_/X sky130_fd_sc_hd__mux2_1
X_15685_ _15683_/Y _15684_/X _15681_/Y vssd1 vssd1 vccd1 vccd1 _15685_/Y sky130_fd_sc_hd__a21oi_2
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 _18949_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ _12871_/A _12871_/B _12896_/X vssd1 vssd1 vccd1 vccd1 _13116_/A sky130_fd_sc_hd__a21o_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_361 _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_372 _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17424_ _17421_/Y _17423_/X _17460_/A2 vssd1 vssd1 vccd1 vccd1 _17433_/S sky130_fd_sc_hd__o21a_4
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _19398_/Q _17920_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19398_/D sky130_fd_sc_hd__mux2_1
XANTENNA_383 _16774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _19647_/Q _19953_/Q _19291_/Q _20078_/Q _11848_/S0 _11846_/C vssd1 vssd1
+ vccd1 vccd1 _11848_/X sky130_fd_sc_hd__mux4_1
XFILLER_221_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_394 _15807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _20226_/Q _17363_/A2 _17354_/X _18692_/A vssd1 vssd1 vccd1 vccd1 _20226_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14567_ _17919_/A _17919_/B _14567_/C vssd1 vssd1 vccd1 vccd1 _14567_/X sky130_fd_sc_hd__and3_4
XFILLER_159_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11779_ _13523_/A _11779_/B vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__xor2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16306_ _19709_/Q _19710_/Q _16306_/C vssd1 vssd1 vccd1 vccd1 _16308_/B sky130_fd_sc_hd__and3_1
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13518_ _13518_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13518_/X sky130_fd_sc_hd__xor2_1
X_17286_ _20201_/Q _17331_/A2 _17285_/X _17331_/C1 vssd1 vssd1 vccd1 vccd1 _20201_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14498_ _19276_/Q _17929_/A1 _14516_/S vssd1 vssd1 vccd1 vccd1 _19276_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19025_ _21031_/Q _19015_/B _19024_/X _18730_/A vssd1 vssd1 vccd1 vccd1 _21031_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_256_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ _13441_/X _16237_/B vssd1 vssd1 vccd1 vccd1 _16237_/X sky130_fd_sc_hd__and2b_1
X_13449_ _19226_/Q _13449_/B vssd1 vssd1 vccd1 vccd1 _13450_/B sky130_fd_sc_hd__nor2_1
XFILLER_127_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_75_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20561_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16168_ _19608_/Q _15671_/X _16170_/S vssd1 vssd1 vccd1 vccd1 _16169_/B sky130_fd_sc_hd__mux2_1
XFILLER_182_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15119_ _15468_/A _15983_/B vssd1 vssd1 vccd1 vccd1 _15119_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16099_ _09664_/X _09665_/X _16079_/B vssd1 vssd1 vccd1 vccd1 _16099_/X sky130_fd_sc_hd__a21bo_1
XFILLER_173_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19927_ _20084_/CLK _19927_/D vssd1 vssd1 vccd1 vccd1 _19927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19858_ _20862_/CLK _19858_/D vssd1 vssd1 vccd1 vccd1 _19858_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09611_ _09686_/A _12976_/B _09686_/C vssd1 vssd1 vccd1 vccd1 _09643_/A sky130_fd_sc_hd__or3_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18809_ _19091_/Q _12589_/B _12592_/C _13568_/Y vssd1 vssd1 vccd1 vccd1 _18809_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19789_ _20712_/CLK _19789_/D vssd1 vssd1 vccd1 vccd1 _19789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09542_ _19153_/Q _14112_/B vssd1 vssd1 vccd1 vccd1 _13867_/A sky130_fd_sc_hd__nor2_4
XFILLER_225_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20702_ _20702_/CLK _20702_/D vssd1 vssd1 vccd1 vccd1 _20702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20633_ _20633_/CLK _20633_/D vssd1 vssd1 vccd1 vccd1 _20633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20564_ _20586_/CLK _20564_/D vssd1 vssd1 vccd1 vccd1 _20564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20495_ _20662_/CLK _20495_/D vssd1 vssd1 vccd1 vccd1 _20495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1207 _15220_/X vssd1 vssd1 vccd1 vccd1 _16056_/B1 sky130_fd_sc_hd__buf_6
Xfanout1218 _14444_/X vssd1 vssd1 vccd1 vccd1 _14483_/S sky130_fd_sc_hd__buf_8
Xfanout1229 _12493_/A vssd1 vssd1 vccd1 vccd1 _15526_/A sky130_fd_sc_hd__buf_6
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21047_ _21047_/A vssd1 vssd1 vccd1 vccd1 _21047_/X sky130_fd_sc_hd__buf_2
XFILLER_87_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09809_ _12059_/A1 _09808_/X _09805_/X _12059_/C1 vssd1 vssd1 vccd1 vccd1 _09809_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_275_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12820_ _12906_/A _12820_/B vssd1 vssd1 vccd1 vccd1 _13253_/B sky130_fd_sc_hd__xnor2_2
XFILLER_264_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _19157_/Q _12479_/X _16005_/A1 _12710_/B vssd1 vssd1 vccd1 vccd1 _12751_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11702_ _09834_/A _19384_/Q _20675_/Q _10628_/S vssd1 vssd1 vccd1 vccd1 _11702_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15470_ _10456_/Y _12471_/X _14843_/S _15736_/B _15468_/Y vssd1 vssd1 vccd1 vccd1
+ _15470_/X sky130_fd_sc_hd__o221a_1
X_12682_ _12682_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _12682_/Y sky130_fd_sc_hd__nand2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _20296_/Q _14431_/A2 _14431_/B1 input238/X vssd1 vssd1 vccd1 vccd1 _14423_/B
+ sky130_fd_sc_hd__a22o_2
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _19785_/Q _11641_/S _10622_/S _12023_/S vssd1 vssd1 vccd1 vccd1 _11633_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_230_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _20108_/Q _17942_/A1 _17144_/S vssd1 vssd1 vccd1 vccd1 _20108_/D sky130_fd_sc_hd__mux2_1
X_14352_ _19517_/Q _14352_/B vssd1 vssd1 vccd1 vccd1 _14353_/B sky130_fd_sc_hd__nor2_1
X_11564_ _19639_/Q _19945_/Q _19283_/Q _20070_/Q _09931_/S _09986_/C vssd1 vssd1 vccd1
+ vccd1 _11564_/X sky130_fd_sc_hd__mux4_2
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ _13303_/A _13303_/B _13303_/C vssd1 vssd1 vccd1 vccd1 _13303_/X sky130_fd_sc_hd__and3_1
X_10515_ _10513_/X _10514_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__mux2_1
X_17071_ _20043_/Q _17835_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20043_/D sky130_fd_sc_hd__mux2_1
X_11495_ _11495_/A _11734_/B vssd1 vssd1 vccd1 vccd1 _11497_/B sky130_fd_sc_hd__nand2_1
X_14283_ _14283_/A _14283_/B vssd1 vssd1 vccd1 vccd1 _14283_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16022_ _16050_/A1 _16021_/X _16009_/X vssd1 vssd1 vccd1 vccd1 _16022_/X sky130_fd_sc_hd__a21o_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13234_ _13233_/A _13233_/C _13233_/B vssd1 vssd1 vccd1 vccd1 _13234_/Y sky130_fd_sc_hd__o21ai_1
X_10446_ _12073_/A1 _10442_/X _10445_/X _12059_/C1 vssd1 vssd1 vccd1 vccd1 _10446_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_171_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10377_ _10465_/A _10377_/B vssd1 vssd1 vccd1 vccd1 _10377_/Y sky130_fd_sc_hd__nand2_1
XFILLER_152_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _13166_/B _13166_/C vssd1 vssd1 vccd1 vccd1 _13418_/B sky130_fd_sc_hd__and2_2
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12116_ _13433_/A _11958_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _12206_/B sky130_fd_sc_hd__a21o_1
X_17973_ _20729_/Q _17976_/C vssd1 vssd1 vccd1 vccd1 _17975_/A sky130_fd_sc_hd__and2_1
XFILLER_3_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13096_ _20977_/Q _13096_/B vssd1 vssd1 vccd1 vccd1 _13097_/B sky130_fd_sc_hd__xnor2_2
XFILLER_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19712_ _20795_/CLK _19712_/D vssd1 vssd1 vccd1 vccd1 _19712_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1730 _09504_/Y vssd1 vssd1 vccd1 vccd1 _18765_/A sky130_fd_sc_hd__clkbuf_16
X_16924_ _16974_/A1 _16923_/X _16982_/B1 vssd1 vssd1 vccd1 vccd1 _16924_/Y sky130_fd_sc_hd__o21ai_2
X_12047_ _10430_/S _20715_/Q _12053_/S _12046_/X vssd1 vssd1 vccd1 vccd1 _12047_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout1741 _09695_/A vssd1 vssd1 vccd1 vccd1 _12304_/C1 sky130_fd_sc_hd__buf_6
XFILLER_242_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1752 _09501_/Y vssd1 vssd1 vccd1 vccd1 _10308_/S sky130_fd_sc_hd__buf_12
XFILLER_172_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1763 _13582_/A vssd1 vssd1 vccd1 vccd1 _12584_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1774 output482/A vssd1 vssd1 vccd1 vccd1 _13552_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_78_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_193_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19541_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_266_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16855_ _16884_/S input82/X vssd1 vssd1 vccd1 vccd1 _16855_/Y sky130_fd_sc_hd__nand2_1
X_19643_ _20717_/CLK _19643_/D vssd1 vssd1 vccd1 vccd1 _19643_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1785 _18223_/B vssd1 vssd1 vccd1 vccd1 _18313_/B sky130_fd_sc_hd__buf_12
XFILLER_253_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1796 _20184_/Q vssd1 vssd1 vccd1 vccd1 _18209_/A1 sky130_fd_sc_hd__buf_8
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_122_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20004_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15806_ _19756_/Q _15999_/A2 _15805_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15806_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_281_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19574_ _19574_/CLK _19574_/D vssd1 vssd1 vccd1 vccd1 _19574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16786_ _19090_/Q _16996_/B1 _16785_/X vssd1 vssd1 vccd1 vccd1 _16786_/X sky130_fd_sc_hd__o21a_1
X_13998_ _09731_/A _14031_/A2 _14040_/B1 _13997_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1
+ _19166_/D sky130_fd_sc_hd__o221a_1
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18525_ _18980_/A _18525_/B vssd1 vssd1 vccd1 vccd1 _20901_/D sky130_fd_sc_hd__nor2_1
XFILLER_234_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ _11743_/B _15984_/A2 _15984_/B1 _11741_/A _15890_/A vssd1 vssd1 vccd1 vccd1
+ _15737_/X sky130_fd_sc_hd__a221o_1
X_12949_ _19266_/Q _19265_/Q _19264_/Q vssd1 vssd1 vccd1 vccd1 _12949_/X sky130_fd_sc_hd__or3_4
XFILLER_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18456_ _18981_/B _18563_/C vssd1 vssd1 vccd1 vccd1 _18457_/C sky130_fd_sc_hd__nor2_2
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15668_ _16046_/A1 _15667_/X _15663_/X vssd1 vssd1 vccd1 vccd1 _15668_/X sky130_fd_sc_hd__o21a_2
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 _19228_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_191 _19158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17407_ _20258_/Q _20250_/Q _17442_/A vssd1 vssd1 vccd1 vccd1 _17407_/X sky130_fd_sc_hd__mux2_1
X_14619_ _19383_/Q _17903_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19383_/D sky130_fd_sc_hd__mux2_1
X_18387_ _18560_/B _18387_/B vssd1 vssd1 vccd1 vccd1 _18387_/Y sky130_fd_sc_hd__nand2_1
X_15599_ _20929_/Q _15995_/A2 _15598_/X vssd1 vssd1 vccd1 vccd1 _15599_/X sky130_fd_sc_hd__o21a_1
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17338_ _17236_/A _17364_/A2 _17362_/B1 _20266_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17338_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ _17269_/A _17275_/B _17269_/C vssd1 vssd1 vccd1 vccd1 _17269_/X sky130_fd_sc_hd__and3_1
XFILLER_119_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19008_ _18215_/Y _18982_/B _19016_/B1 _19007_/X vssd1 vssd1 vccd1 vccd1 _21023_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20280_ _20990_/CLK _20280_/D vssd1 vssd1 vccd1 vccd1 _20280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ input46/X vssd1 vssd1 vccd1 vccd1 _09525_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20616_ _20706_/CLK _20616_/D vssd1 vssd1 vccd1 vccd1 _20616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20547_ _20679_/CLK _20547_/D vssd1 vssd1 vccd1 vccd1 _20547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10300_ _19476_/Q _09695_/Y _10299_/X _10308_/S vssd1 vssd1 vccd1 vccd1 _10300_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_119_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11280_ _09569_/A _13641_/B _11279_/X vssd1 vssd1 vccd1 vccd1 _11280_/Y sky130_fd_sc_hd__o21ai_2
X_20478_ _20645_/CLK _20478_/D vssd1 vssd1 vccd1 vccd1 _20478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10231_ _10229_/X _10230_/X _10235_/S vssd1 vssd1 vccd1 vccd1 _10231_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10162_ _11012_/A _10161_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _10162_/X sky130_fd_sc_hd__o21a_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1004 _15606_/A1 vssd1 vssd1 vccd1 vccd1 _15019_/A sky130_fd_sc_hd__buf_8
Xfanout1015 _14880_/Y vssd1 vssd1 vccd1 vccd1 _15185_/B sky130_fd_sc_hd__buf_4
Xoutput390 _13813_/X vssd1 vssd1 vccd1 vccd1 din0[22] sky130_fd_sc_hd__buf_4
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1026 _17004_/A2 vssd1 vssd1 vccd1 vccd1 _16870_/A2 sky130_fd_sc_hd__buf_4
X_14970_ _15314_/B _15314_/C _15314_/D vssd1 vssd1 vccd1 vccd1 _14971_/C sky130_fd_sc_hd__nor3_1
Xfanout1037 _17852_/A1 vssd1 vssd1 vccd1 vccd1 _17886_/A1 sky130_fd_sc_hd__buf_4
XFILLER_120_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10093_ _10091_/X _10092_/X _12426_/S vssd1 vssd1 vccd1 vccd1 _10093_/X sky130_fd_sc_hd__mux2_1
Xfanout1048 _11049_/B1 vssd1 vssd1 vccd1 vccd1 _17855_/A1 sky130_fd_sc_hd__buf_4
Xfanout1059 _10813_/X vssd1 vssd1 vccd1 vccd1 _17925_/A1 sky130_fd_sc_hd__buf_6
XFILLER_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13921_ _13921_/A _13921_/B vssd1 vssd1 vccd1 vccd1 _13921_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ _19897_/Q _17886_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19897_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13852_ _17442_/A _20254_/Q _17438_/B _17231_/A _13851_/X vssd1 vssd1 vccd1 vccd1
+ _13852_/X sky130_fd_sc_hd__a32o_4
XFILLER_207_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12803_ _12906_/A _12803_/B vssd1 vssd1 vccd1 vccd1 _13264_/A sky130_fd_sc_hd__xnor2_4
X_16571_ _16593_/A _16571_/B vssd1 vssd1 vccd1 vccd1 _19851_/D sky130_fd_sc_hd__or2_1
XFILLER_62_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13783_ _13612_/A split3/A _13524_/Y _13522_/Y _16240_/A1 vssd1 vssd1 vccd1 vccd1
+ _13783_/X sky130_fd_sc_hd__a32o_4
X_10995_ _09502_/A _10982_/X _10985_/X _10994_/X _09689_/A vssd1 vssd1 vccd1 vccd1
+ _11012_/B sky130_fd_sc_hd__o311a_1
X_18310_ _18556_/B vssd1 vssd1 vccd1 vccd1 _18310_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_43_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _15589_/S _15494_/A _15520_/X _15521_/Y vssd1 vssd1 vccd1 vccd1 _15522_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19290_ _20077_/CLK _19290_/D vssd1 vssd1 vccd1 vccd1 _19290_/Q sky130_fd_sc_hd__dfxtp_1
X_12734_ _12736_/B _12736_/C _12736_/A vssd1 vssd1 vccd1 vccd1 _12749_/A sky130_fd_sc_hd__a21oi_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18241_ _20802_/Q _18240_/Y _18316_/S vssd1 vssd1 vccd1 vccd1 _18242_/B sky130_fd_sc_hd__mux2_1
X_15453_ _19744_/Q _15453_/A2 _15445_/X _15021_/A _15452_/X vssd1 vssd1 vccd1 vccd1
+ _15453_/X sky130_fd_sc_hd__a221o_1
XFILLER_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12666_/A sky130_fd_sc_hd__nor2_1
XFILLER_124_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _19521_/Q _14392_/B _14403_/X vssd1 vssd1 vccd1 vccd1 _14405_/B sky130_fd_sc_hd__o21ai_4
X_18172_ _18416_/A _18172_/B vssd1 vssd1 vccd1 vccd1 _20788_/D sky130_fd_sc_hd__and2_1
X_11616_ _20169_/Q _11616_/B vssd1 vssd1 vccd1 vccd1 _11616_/X sky130_fd_sc_hd__or2_1
X_15384_ _14983_/A _15314_/D _15016_/Y vssd1 vssd1 vccd1 vccd1 _15384_/Y sky130_fd_sc_hd__o21ai_2
X_12596_ _19495_/Q _12664_/C _19496_/Q vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__o21a_1
XFILLER_168_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17123_ _20091_/Q _17925_/A1 _17132_/S vssd1 vssd1 vccd1 vccd1 _20091_/D sky130_fd_sc_hd__mux2_1
X_14335_ _14427_/A _14335_/B _14343_/B vssd1 vssd1 vccd1 vccd1 _14335_/X sky130_fd_sc_hd__or3b_1
XFILLER_117_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11547_ _09986_/A _19382_/Q _20673_/Q _12174_/S vssd1 vssd1 vccd1 vccd1 _11547_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17054_ _20026_/Q _17750_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20026_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14266_ _19229_/Q _14398_/A2 _14265_/X _14772_/C1 vssd1 vssd1 vccd1 vccd1 _19229_/D
+ sky130_fd_sc_hd__o211a_1
X_11478_ _12011_/S _11475_/X _11477_/X _12183_/C1 vssd1 vssd1 vccd1 vccd1 _11478_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16005_ _16005_/A1 _12624_/X _16004_/X _12832_/B vssd1 vssd1 vccd1 vccd1 _16007_/B
+ sky130_fd_sc_hd__a22o_1
X_13217_ _20973_/Q _13272_/B _13215_/X _13216_/Y _18767_/A vssd1 vssd1 vccd1 vccd1
+ _13218_/C sky130_fd_sc_hd__a221o_2
X_10429_ _12060_/A1 _19473_/Q _19441_/Q _10428_/S vssd1 vssd1 vccd1 vccd1 _10429_/X
+ sky130_fd_sc_hd__a22o_1
X_14197_ _19502_/Q _14198_/B vssd1 vssd1 vccd1 vccd1 _14197_/Y sky130_fd_sc_hd__nor2_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13148_ _15264_/A _13538_/B _10885_/A vssd1 vssd1 vccd1 vccd1 _13541_/B sky130_fd_sc_hd__a21oi_4
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17956_ _20723_/Q _17959_/C vssd1 vssd1 vccd1 vccd1 _17962_/C sky130_fd_sc_hd__and2_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _13303_/A _13303_/C _13303_/B vssd1 vssd1 vccd1 vccd1 _13368_/A sky130_fd_sc_hd__a21boi_4
XFILLER_66_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1560 _10842_/S vssd1 vssd1 vccd1 vccd1 _12389_/S sky130_fd_sc_hd__buf_6
XFILLER_39_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16907_ _16981_/A1 _15725_/X _16879_/X _16906_/X vssd1 vssd1 vccd1 vccd1 _16907_/X
+ sky130_fd_sc_hd__o211a_2
X_17887_ _20658_/Q _17887_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20658_/D sky130_fd_sc_hd__mux2_1
Xfanout1571 _09624_/Y vssd1 vssd1 vccd1 vccd1 _12151_/C1 sky130_fd_sc_hd__buf_8
Xfanout1582 _11353_/C1 vssd1 vssd1 vccd1 vccd1 _12314_/C1 sky130_fd_sc_hd__buf_4
XFILLER_239_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1593 _11363_/A1 vssd1 vssd1 vccd1 vccd1 _12318_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19626_ _20657_/CLK _19626_/D vssd1 vssd1 vccd1 vccd1 _19626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16838_ _16846_/A _09524_/Y _16809_/X _16837_/Y vssd1 vssd1 vccd1 vccd1 _16838_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_66_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19557_ _19609_/CLK _19557_/D vssd1 vssd1 vccd1 vccd1 _19557_/Q sky130_fd_sc_hd__dfxtp_4
X_16769_ input87/X input72/X _16769_/S vssd1 vssd1 vccd1 vccd1 _16770_/A sky130_fd_sc_hd__mux2_2
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18508_ _18612_/B _18508_/B vssd1 vssd1 vccd1 vccd1 _18508_/X sky130_fd_sc_hd__or2_1
XFILLER_62_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19488_ _20583_/CLK _19488_/D vssd1 vssd1 vccd1 vccd1 _19488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18439_ _20874_/Q _18280_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18440_/B sky130_fd_sc_hd__mux2_1
XFILLER_210_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19590_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401_ _20667_/CLK _20401_/D vssd1 vssd1 vccd1 vccd1 _20401_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_174_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20332_ _20687_/CLK _20332_/D vssd1 vssd1 vccd1 vccd1 _20332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20263_ _20263_/CLK _20263_/D vssd1 vssd1 vccd1 vccd1 _20263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20194_ _20428_/CLK _20194_/D vssd1 vssd1 vccd1 vccd1 _20194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_249_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput107 dout1[0] vssd1 vssd1 vccd1 vccd1 input107/X sky130_fd_sc_hd__clkbuf_2
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput118 dout1[1] vssd1 vssd1 vccd1 vccd1 input118/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput129 dout1[2] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__clkbuf_2
XFILLER_131_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09508_ _19165_/Q vssd1 vssd1 vccd1 vccd1 _09508_/Y sky130_fd_sc_hd__inv_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10778_/X _10779_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _10781_/B sky130_fd_sc_hd__mux2_1
XFILLER_13_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12450_ _12450_/A _12450_/B vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__and2_1
XFILLER_184_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _15374_/S _11401_/B vssd1 vssd1 vccd1 vccd1 _11774_/B sky130_fd_sc_hd__nor2_2
XFILLER_21_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12381_ _20395_/Q _20459_/Q _12381_/S vssd1 vssd1 vccd1 vccd1 _12381_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_80 _09750_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_91 _11807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _14121_/A _16710_/B vssd1 vssd1 vccd1 vccd1 _14120_/Y sky130_fd_sc_hd__nor2_2
XFILLER_193_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11332_ _20469_/Q _20309_/Q _11342_/S vssd1 vssd1 vccd1 vccd1 _11332_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14051_ _14081_/A _14069_/B _14051_/C vssd1 vssd1 vccd1 vccd1 _14051_/X sky130_fd_sc_hd__or3_1
XFILLER_137_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11263_ _20333_/Q _11270_/A2 _09688_/B _11250_/S vssd1 vssd1 vccd1 vccd1 _11263_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ _13002_/A _13002_/B vssd1 vssd1 vccd1 vccd1 _13002_/Y sky130_fd_sc_hd__nor2_1
X_10214_ _11338_/A1 _10211_/X _10213_/X vssd1 vssd1 vccd1 vccd1 _10214_/X sky130_fd_sc_hd__a21o_1
XFILLER_180_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11194_ _11192_/X _11193_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _11194_/X sky130_fd_sc_hd__mux2_1
XFILLER_268_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17810_ _20587_/Q _17950_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20587_/D sky130_fd_sc_hd__mux2_1
X_10145_ _20035_/Q _12296_/S vssd1 vssd1 vccd1 vccd1 _10145_/X sky130_fd_sc_hd__or2_1
X_18790_ _19088_/Q _18785_/A2 _12591_/X _13524_/A vssd1 vssd1 vccd1 vccd1 _18790_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ _20522_/Q _17881_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20522_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14953_ _15314_/B _15020_/A vssd1 vssd1 vccd1 vccd1 _15308_/C sky130_fd_sc_hd__nor2_2
X_10076_ _13670_/A1 _17898_/A1 _10075_/X _12075_/C1 vssd1 vssd1 vccd1 vccd1 _13684_/A
+ sky130_fd_sc_hd__o211a_2
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _13478_/A _13943_/S _13903_/Y _19117_/Q vssd1 vssd1 vccd1 vccd1 _19117_/D
+ sky130_fd_sc_hd__a22o_1
X_17672_ _20458_/Q _17706_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20458_/D sky130_fd_sc_hd__mux2_1
X_14884_ _15578_/S _14885_/B vssd1 vssd1 vccd1 vccd1 _14884_/X sky130_fd_sc_hd__or2_2
XFILLER_236_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19411_ _20570_/CLK _19411_/D vssd1 vssd1 vccd1 vccd1 _19411_/Q sky130_fd_sc_hd__dfxtp_1
X_16623_ _19882_/Q _17937_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19882_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13835_ _20005_/Q split1/X _13789_/X split2/X vssd1 vssd1 vccd1 vccd1 _13835_/X sky130_fd_sc_hd__a22o_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19342_ _20559_/CLK _19342_/D vssd1 vssd1 vccd1 vccd1 _19342_/Q sky130_fd_sc_hd__dfxtp_1
X_16554_ _19843_/Q _16578_/A2 _16578_/B1 input13/X vssd1 vssd1 vccd1 vccd1 _16555_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ _12245_/Y _13730_/B _13776_/B1 vssd1 vssd1 vccd1 vccd1 _13769_/A sky130_fd_sc_hd__o21a_2
X_10978_ _10127_/A _10973_/Y _10977_/X _10971_/X vssd1 vssd1 vccd1 vccd1 _10978_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15505_ _15283_/A _15504_/Y _15096_/B vssd1 vssd1 vccd1 vccd1 _15505_/X sky130_fd_sc_hd__a21o_1
X_19273_ _20467_/CLK _19273_/D vssd1 vssd1 vccd1 vccd1 _19273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12717_ _19507_/Q _12740_/B _19508_/Q vssd1 vssd1 vccd1 vccd1 _12718_/B sky130_fd_sc_hd__a21oi_1
X_16485_ _19794_/Q _17112_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19794_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13697_ _16598_/C _13697_/B vssd1 vssd1 vccd1 vccd1 _13697_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18224_ _18223_/B _14249_/B _18223_/Y vssd1 vssd1 vccd1 vccd1 _18505_/B sky130_fd_sc_hd__o21ai_4
XFILLER_188_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15436_ _15261_/X _15435_/X _15578_/S vssd1 vssd1 vccd1 vccd1 _15437_/B sky130_fd_sc_hd__mux2_4
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _14803_/A1 _12657_/A2 _12682_/B _12647_/X vssd1 vssd1 vccd1 vccd1 _12648_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18155_ _18563_/A _18390_/A vssd1 vssd1 vccd1 vccd1 _18690_/A sky130_fd_sc_hd__or2_4
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15367_ _10685_/Y _15366_/X _15492_/A vssd1 vssd1 vccd1 vccd1 _15367_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_156_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12579_ _13869_/A _12579_/B _12579_/C _12579_/D vssd1 vssd1 vccd1 vccd1 _12978_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17106_ _20076_/Q _17874_/A1 _17111_/S vssd1 vssd1 vccd1 vccd1 _20076_/D sky130_fd_sc_hd__mux2_1
X_14318_ _14397_/A _14397_/B _14318_/C vssd1 vssd1 vccd1 vccd1 _14318_/X sky130_fd_sc_hd__or3_1
X_18086_ _18086_/A _18086_/B _18087_/B vssd1 vssd1 vccd1 vccd1 _20769_/D sky130_fd_sc_hd__nor3_1
X_15298_ _10798_/X _15500_/A0 _12470_/Y _13541_/A _12579_/D vssd1 vssd1 vccd1 vccd1
+ _15298_/X sky130_fd_sc_hd__a221o_1
XFILLER_172_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17037_ _20015_/Q _12928_/B _17038_/S vssd1 vssd1 vccd1 vccd1 _20015_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14249_ _19507_/Q _14249_/B vssd1 vssd1 vccd1 vccd1 _14250_/C sky130_fd_sc_hd__xnor2_1
XFILLER_171_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout808 _18974_/B1 vssd1 vssd1 vccd1 vccd1 _18967_/B1 sky130_fd_sc_hd__buf_4
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout819 _15633_/Y vssd1 vssd1 vccd1 vccd1 fanout819/X sky130_fd_sc_hd__buf_2
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09790_ _10561_/A _09789_/X _09785_/X vssd1 vssd1 vccd1 vccd1 _09790_/X sky130_fd_sc_hd__a21o_4
XFILLER_140_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18988_ _18165_/Y _18983_/B _19016_/B1 _18987_/X vssd1 vssd1 vccd1 vccd1 _21013_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _20708_/Q _17939_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20708_/D sky130_fd_sc_hd__mux2_1
XFILLER_273_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1390 _12165_/S vssd1 vssd1 vccd1 vccd1 _12182_/S sky130_fd_sc_hd__buf_6
X_20950_ _21013_/CLK _20950_/D vssd1 vssd1 vccd1 vccd1 _20950_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19609_ _19609_/CLK _19609_/D vssd1 vssd1 vccd1 vccd1 _19609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20881_ _21041_/CLK _20881_/D vssd1 vssd1 vccd1 vccd1 _20881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20315_ _20315_/CLK _20315_/D vssd1 vssd1 vccd1 vccd1 _20315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20246_ _20296_/CLK _20246_/D vssd1 vssd1 vccd1 vccd1 _20246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20177_ _20716_/CLK _20177_/D vssd1 vssd1 vccd1 vccd1 _20177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09988_ _19643_/Q _19949_/Q _19287_/Q _20074_/Q _11932_/S0 _12003_/C vssd1 vssd1
+ vccd1 vccd1 _09988_/X sky130_fd_sc_hd__mux4_1
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _12020_/C1 _11949_/X _11872_/A vssd1 vssd1 vccd1 vccd1 _11950_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_273_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _19370_/Q _11009_/A2 _10899_/X _09688_/A _10900_/X vssd1 vssd1 vccd1 vccd1
+ _10901_/X sky130_fd_sc_hd__o221a_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11881_ _13419_/A _11752_/B _11733_/Y vssd1 vssd1 vccd1 vccd1 _11882_/B sky130_fd_sc_hd__o21ai_1
XFILLER_264_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13620_ _13626_/A1 _13345_/X _13427_/B _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13620_/X
+ sky130_fd_sc_hd__a22o_2
X_10832_ _09621_/A _10831_/X _10828_/X _12385_/C1 vssd1 vssd1 vccd1 vccd1 _10832_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13551_ _20952_/Q _13564_/B _13550_/X vssd1 vssd1 vccd1 vccd1 _13552_/C sky130_fd_sc_hd__a21bo_1
XFILLER_73_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10763_ _11012_/A _10761_/X _10762_/X vssd1 vssd1 vccd1 vccd1 _13657_/B sky130_fd_sc_hd__o21ai_4
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ _19163_/Q _19161_/Q _12502_/C vssd1 vssd1 vccd1 vccd1 _14808_/A sky130_fd_sc_hd__or3_4
XFILLER_41_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16270_ _19686_/Q _17804_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19686_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13482_ _13482_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _15127_/A sky130_fd_sc_hd__xor2_4
X_10694_ _20404_/Q _20340_/Q _20632_/Q _20596_/Q _11116_/S _12406_/C vssd1 vssd1 vccd1
+ vccd1 _10694_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15221_ _15221_/A _15259_/B vssd1 vssd1 vccd1 vccd1 _15221_/Y sky130_fd_sc_hd__nor2_1
X_12433_ _12433_/A1 _17916_/A1 _12432_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _16009_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_201_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15152_ _15326_/A _15126_/X _15128_/X _15151_/Y vssd1 vssd1 vccd1 vccd1 _15152_/X
+ sky130_fd_sc_hd__o31a_1
X_12364_ _12449_/A vssd1 vssd1 vccd1 vccd1 _12447_/A sky130_fd_sc_hd__inv_2
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14103_ _14105_/A _14107_/B _14103_/C vssd1 vssd1 vccd1 vccd1 _14103_/X sky130_fd_sc_hd__or3_1
XFILLER_154_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11315_ _15062_/S _11783_/B vssd1 vssd1 vccd1 vccd1 _15075_/B sky130_fd_sc_hd__nor2_1
XFILLER_4_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19960_ _20664_/CLK _19960_/D vssd1 vssd1 vccd1 vccd1 _19960_/Q sky130_fd_sc_hd__dfxtp_1
X_15083_ _20883_/Q _14971_/A _15566_/B1 _15082_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15083_/X sky130_fd_sc_hd__a221o_1
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12295_ _19960_/Q _12295_/B vssd1 vssd1 vccd1 vccd1 _12295_/X sky130_fd_sc_hd__or2_1
XFILLER_268_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14034_ _19178_/Q _14043_/A2 _14034_/B1 _14033_/X _16129_/B1 vssd1 vssd1 vccd1 vccd1
+ _19178_/D sky130_fd_sc_hd__o221a_1
XFILLER_153_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18911_ _18529_/X _18971_/B _18909_/X _18910_/Y vssd1 vssd1 vccd1 vccd1 _18912_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11246_ _11246_/A1 _11245_/Y _09613_/A vssd1 vssd1 vccd1 vccd1 _11246_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19891_ _20583_/CLK _19891_/D vssd1 vssd1 vccd1 vccd1 _19891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18842_ _18842_/A _18842_/B vssd1 vssd1 vccd1 vccd1 _20991_/D sky130_fd_sc_hd__nor2_1
X_11177_ _19399_/Q _11169_/B _11259_/S vssd1 vssd1 vccd1 vccd1 _11177_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10128_ _19540_/Q _09596_/B _10114_/X _10127_/Y vssd1 vssd1 vccd1 vccd1 _10128_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_249_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18773_ _19085_/Q _12589_/B _12591_/X _15076_/A vssd1 vssd1 vccd1 vccd1 _18773_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_15985_ _13182_/A _12565_/B _15984_/X vssd1 vssd1 vccd1 vccd1 _15985_/Y sky130_fd_sc_hd__a21oi_1
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14936_ _19702_/Q _15475_/A2 _15475_/B1 _19734_/Q vssd1 vssd1 vccd1 vccd1 _14936_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_208_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17724_ _20505_/Q _17898_/A1 _17738_/S vssd1 vssd1 vccd1 vccd1 _20505_/D sky130_fd_sc_hd__mux2_1
X_10059_ _11281_/A _20601_/Q _11268_/C vssd1 vssd1 vccd1 vccd1 _10059_/X sky130_fd_sc_hd__and3_1
XFILLER_250_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20690_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14867_ _11783_/B _14882_/A _14870_/S vssd1 vssd1 vccd1 vccd1 _14867_/X sky130_fd_sc_hd__mux2_1
X_17655_ _20441_/Q _17932_/A1 _17669_/S vssd1 vssd1 vccd1 vccd1 _20441_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16606_ _19865_/Q _17920_/A1 _16620_/S vssd1 vssd1 vccd1 vccd1 _19865_/D sky130_fd_sc_hd__mux2_1
X_13818_ _13822_/A1 _13760_/B split9/X input234/X vssd1 vssd1 vccd1 vccd1 _13818_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17586_ _20344_/Q split4/X _17601_/S vssd1 vssd1 vccd1 vccd1 _20344_/D sky130_fd_sc_hd__mux2_1
X_14798_ _19146_/Q _14798_/A2 _14797_/X _16187_/A vssd1 vssd1 vccd1 vccd1 _19523_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16537_ _16557_/A _16537_/B vssd1 vssd1 vccd1 vccd1 _19834_/D sky130_fd_sc_hd__or2_1
X_19325_ _20047_/CLK _19325_/D vssd1 vssd1 vccd1 vccd1 _19325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13749_ _13749_/A _13749_/B vssd1 vssd1 vccd1 vccd1 _13750_/B sky130_fd_sc_hd__nor2_8
XFILLER_250_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19256_ _21013_/CLK _19256_/D vssd1 vssd1 vccd1 vccd1 _19256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16468_ _19777_/Q _17163_/A1 _16471_/S vssd1 vssd1 vccd1 vccd1 _19777_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18207_ _18414_/A _18207_/B vssd1 vssd1 vccd1 vccd1 _20795_/D sky130_fd_sc_hd__and2_1
XFILLER_176_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15419_ _20955_/Q _15568_/A2 _15568_/B1 _20827_/Q _15418_/X vssd1 vssd1 vccd1 vccd1
+ _15419_/X sky130_fd_sc_hd__a221o_4
X_19187_ _21044_/CLK _19187_/D vssd1 vssd1 vccd1 vccd1 _19187_/Q sky130_fd_sc_hd__dfxtp_1
X_16399_ _19745_/Q _16402_/C _18086_/A vssd1 vssd1 vccd1 vccd1 _16399_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_157_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18138_ _18138_/A _18138_/B vssd1 vssd1 vccd1 vccd1 _18139_/B sky130_fd_sc_hd__and2_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18069_ _20763_/Q _20762_/Q _18069_/C vssd1 vssd1 vccd1 vccd1 _18071_/B sky130_fd_sc_hd__and3_1
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20100_ _20703_/CLK _20100_/D vssd1 vssd1 vccd1 vccd1 _20100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09911_ _19644_/Q _19950_/Q _19288_/Q _20075_/Q _12174_/S _11851_/C vssd1 vssd1 vccd1
+ vccd1 _09911_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout605 _14601_/X vssd1 vssd1 vccd1 vccd1 _14633_/S sky130_fd_sc_hd__buf_12
XFILLER_259_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout616 _14488_/X vssd1 vssd1 vccd1 vccd1 _14516_/S sky130_fd_sc_hd__buf_6
X_20031_ _20438_/CLK _20031_/D vssd1 vssd1 vccd1 vccd1 _20031_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout627 _13902_/Y vssd1 vssd1 vccd1 vccd1 _14043_/B1 sky130_fd_sc_hd__clkbuf_8
X_09842_ _09840_/X _09841_/X _12082_/S vssd1 vssd1 vccd1 vccd1 _09842_/X sky130_fd_sc_hd__mux2_1
Xfanout638 _16876_/A vssd1 vssd1 vccd1 vccd1 _17012_/A2 sky130_fd_sc_hd__buf_4
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout649 _16077_/B vssd1 vssd1 vccd1 vccd1 _16131_/A2 sky130_fd_sc_hd__buf_2
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09773_ _12007_/A1 _19357_/Q _20712_/Q _12013_/S _12016_/C1 vssd1 vssd1 vccd1 vccd1
+ _09773_/X sky130_fd_sc_hd__a221o_1
XFILLER_112_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20933_ _20998_/CLK _20933_/D vssd1 vssd1 vccd1 vccd1 _20933_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20864_ _21020_/CLK _20864_/D vssd1 vssd1 vccd1 vccd1 _20864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20795_ _20795_/CLK _20795_/D vssd1 vssd1 vccd1 vccd1 _20795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11100_ _12569_/A _13646_/B _11099_/Y _11281_/B vssd1 vssd1 vccd1 vccd1 _11100_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_135_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12080_ _19824_/Q _10603_/B _12078_/X _12085_/B2 _12079_/X vssd1 vssd1 vccd1 vccd1
+ _12080_/X sky130_fd_sc_hd__o221a_1
XFILLER_249_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11031_ _20368_/Q _20432_/Q _11039_/S vssd1 vssd1 vccd1 vccd1 _11031_/X sky130_fd_sc_hd__mux2_1
X_20229_ _21016_/CLK _20229_/D vssd1 vssd1 vccd1 vccd1 _20229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15770_ _19723_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15770_/X sky130_fd_sc_hd__or2_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _19217_/Q _12982_/B _12982_/C _14110_/C vssd1 vssd1 vccd1 vccd1 _13498_/B
+ sky130_fd_sc_hd__and4_2
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _19478_/Q _17936_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19478_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _11931_/X _11932_/X _11933_/S vssd1 vssd1 vccd1 vccd1 _11933_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_510 input216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_521 _13626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_532 _13637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _17437_/X _17438_/X _17439_/X _17454_/A _17457_/A vssd1 vssd1 vccd1 vccd1
+ _17443_/B sky130_fd_sc_hd__o32a_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _19414_/Q _17936_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19414_/D sky130_fd_sc_hd__mux2_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_543 _12041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ _11946_/A1 _19486_/Q _19454_/Q _11947_/S _11946_/C1 vssd1 vssd1 vccd1 vccd1
+ _11864_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_554 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_565 _13472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_576 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13603_ _13603_/A _13603_/B vssd1 vssd1 vccd1 vccd1 _13603_/X sky130_fd_sc_hd__or2_2
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _20370_/Q _20434_/Q _12389_/S vssd1 vssd1 vccd1 vccd1 _10815_/X sky130_fd_sc_hd__mux2_1
XANTENNA_587 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17371_ _20234_/Q _17371_/A2 _17370_/X _18720_/A vssd1 vssd1 vccd1 vccd1 _20234_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _19349_/Q _17935_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19349_/D sky130_fd_sc_hd__mux2_1
XFILLER_260_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_598 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11795_ _11795_/A _11795_/B _13416_/A vssd1 vssd1 vccd1 vccd1 _15734_/B sky130_fd_sc_hd__nand3_1
XFILLER_186_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16322_ _19715_/Q _19716_/Q _16322_/C vssd1 vssd1 vccd1 vccd1 _16324_/B sky130_fd_sc_hd__and3_1
X_19110_ _20273_/CLK _19110_/D vssd1 vssd1 vccd1 vccd1 _19110_/Q sky130_fd_sc_hd__dfxtp_4
X_13534_ _13532_/Y _13533_/X _20951_/Q _13564_/B vssd1 vssd1 vccd1 vccd1 _13534_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10746_ _09502_/A _10738_/X _10744_/X _10745_/Y _12385_/C1 vssd1 vssd1 vccd1 vccd1
+ _10746_/X sky130_fd_sc_hd__a221o_4
X_19041_ _21039_/Q _19049_/A2 _19040_/X _18730_/A vssd1 vssd1 vccd1 vccd1 _21039_/D
+ sky130_fd_sc_hd__o211a_1
X_16253_ _19669_/Q _17927_/A1 _16275_/S vssd1 vssd1 vccd1 vccd1 _19669_/D sky130_fd_sc_hd__mux2_1
XFILLER_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_147_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20930_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13465_ _20007_/Q _12948_/X _13464_/X _17015_/B vssd1 vssd1 vccd1 vccd1 _13468_/A
+ sky130_fd_sc_hd__o31a_1
X_10677_ _12399_/A1 _10673_/X _10676_/X _12399_/C1 vssd1 vssd1 vccd1 vccd1 _10677_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15204_ _15282_/A _16754_/B _15188_/X vssd1 vssd1 vccd1 vccd1 _15206_/B sky130_fd_sc_hd__o21ba_1
X_12416_ _12427_/A1 _19492_/Q _19460_/Q _12417_/S _12419_/C1 vssd1 vssd1 vccd1 vccd1
+ _12416_/X sky130_fd_sc_hd__a221o_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16184_ _19616_/Q _15882_/X _16190_/S vssd1 vssd1 vccd1 vccd1 _16185_/B sky130_fd_sc_hd__mux2_1
X_13396_ _13395_/A _13395_/B _13397_/B vssd1 vssd1 vccd1 vccd1 _13396_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15135_ _20884_/Q _14971_/A _15566_/B1 _15132_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15135_/X sky130_fd_sc_hd__a221o_1
XFILLER_154_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12347_ _12347_/A1 _19365_/Q _20720_/Q _12346_/S _12347_/C1 vssd1 vssd1 vccd1 vccd1
+ _12347_/X sky130_fd_sc_hd__a221o_1
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19943_ _20539_/CLK _19943_/D vssd1 vssd1 vccd1 vccd1 _19943_/Q sky130_fd_sc_hd__dfxtp_1
X_15066_ _15050_/X _15065_/X _15066_/S vssd1 vssd1 vccd1 vccd1 _15066_/X sky130_fd_sc_hd__mux2_4
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ _19523_/Q _15988_/A _15949_/A vssd1 vssd1 vccd1 vccd1 _12282_/B sky130_fd_sc_hd__mux2_8
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _14041_/A1 _09672_/B _09672_/C _14041_/B1 _19854_/Q vssd1 vssd1 vccd1 vccd1
+ _14091_/C sky130_fd_sc_hd__o32a_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11229_ _19583_/Q _11228_/X _11229_/S vssd1 vssd1 vccd1 vccd1 _11236_/C sky130_fd_sc_hd__mux2_4
X_19874_ _20706_/CLK _19874_/D vssd1 vssd1 vccd1 vccd1 _19874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18825_ _18600_/Y _18867_/A2 _18823_/Y _18824_/Y vssd1 vssd1 vccd1 vccd1 _18825_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_283_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18756_ _18760_/B _18756_/B vssd1 vssd1 vccd1 vccd1 _18756_/Y sky130_fd_sc_hd__nor2_1
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15968_ _20974_/Q _16045_/A2 _16016_/S _20846_/Q _15967_/X vssd1 vssd1 vccd1 vccd1
+ _15968_/X sky130_fd_sc_hd__a221o_1
XFILLER_271_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17707_ _20491_/Q _17707_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20491_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14919_ _14981_/A _15022_/B vssd1 vssd1 vccd1 vccd1 _14951_/C sky130_fd_sc_hd__nand2b_1
XFILLER_64_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18687_ _19525_/Q _18687_/B vssd1 vssd1 vccd1 vccd1 _18687_/Y sky130_fd_sc_hd__nand2_1
X_15899_ _12207_/Y _15925_/B _15219_/Y _15898_/Y vssd1 vssd1 vccd1 vccd1 _15903_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_224_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17638_ _20394_/Q _17706_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20394_/D sky130_fd_sc_hd__mux2_1
XFILLER_247_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17569_ _20329_/Q _17914_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20329_/D sky130_fd_sc_hd__mux2_1
X_19308_ _20061_/CLK _19308_/D vssd1 vssd1 vccd1 vccd1 _19308_/Q sky130_fd_sc_hd__dfxtp_1
X_20580_ _20580_/CLK _20580_/D vssd1 vssd1 vccd1 vccd1 _20580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19239_ _19246_/CLK _19239_/D vssd1 vssd1 vccd1 vccd1 _19239_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20014_ _20014_/CLK _20014_/D vssd1 vssd1 vccd1 vccd1 _20014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09825_ _13670_/A1 _09790_/X _09824_/X _12075_/C1 vssd1 vssd1 vccd1 vccd1 _13730_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_171_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09756_ _12003_/A _20516_/Q _12185_/S _20548_/Q vssd1 vssd1 vccd1 vccd1 _09756_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _12156_/A1 _09685_/X _09633_/X vssd1 vssd1 vccd1 vccd1 _09687_/X sky130_fd_sc_hd__a21o_1
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20916_ _21015_/CLK _20916_/D vssd1 vssd1 vccd1 vccd1 _20916_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20847_ _21006_/CLK _20847_/D vssd1 vssd1 vccd1 vccd1 _20847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10600_ _19503_/Q _15589_/S vssd1 vssd1 vccd1 vccd1 _10600_/Y sky130_fd_sc_hd__nor2_2
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11580_ _19417_/Q _11978_/S vssd1 vssd1 vccd1 vccd1 _11580_/X sky130_fd_sc_hd__or2_1
X_20778_ _20812_/CLK _20778_/D vssd1 vssd1 vccd1 vccd1 _20778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ _10937_/A _20503_/Q _11203_/S _20535_/Q vssd1 vssd1 vccd1 vccd1 _10531_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _13362_/B _13362_/C _13362_/A vssd1 vssd1 vccd1 vccd1 _13264_/C sky130_fd_sc_hd__a21o_2
X_10462_ input116/X input152/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10462_/X sky130_fd_sc_hd__mux2_8
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12201_ _12202_/A _12202_/B _13183_/A vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__a21o_2
XFILLER_136_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13181_ _13181_/A _13181_/B vssd1 vssd1 vccd1 vccd1 _13188_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10393_ _20312_/Q _10400_/S _10392_/X vssd1 vssd1 vccd1 vccd1 _10393_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12132_ _20489_/Q _20329_/Q _12133_/S vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16940_ _16974_/A1 _16939_/X _13468_/B vssd1 vssd1 vccd1 vccd1 _16940_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_151_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12063_ _20423_/Q _12064_/S _12041_/X _12063_/C1 vssd1 vssd1 vccd1 vccd1 _12063_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1901 _18754_/A vssd1 vssd1 vccd1 vccd1 _18746_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_284_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1912 _18726_/A vssd1 vssd1 vccd1 vccd1 _18724_/A sky130_fd_sc_hd__buf_4
Xfanout1923 _16165_/C1 vssd1 vssd1 vccd1 vccd1 _16087_/B1 sky130_fd_sc_hd__buf_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1934 _18694_/A vssd1 vssd1 vccd1 vccd1 _18698_/A sky130_fd_sc_hd__buf_4
X_11014_ _19160_/Q _12569_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11014_/X sky130_fd_sc_hd__o21ba_1
Xfanout1945 _13890_/C1 vssd1 vssd1 vccd1 vccd1 _17963_/B1 sky130_fd_sc_hd__buf_2
X_16871_ _19230_/Q _16996_/A2 _16996_/B1 _19099_/Q _16870_/X vssd1 vssd1 vccd1 vccd1
+ _16871_/X sky130_fd_sc_hd__o221a_1
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1956 fanout1960/X vssd1 vssd1 vccd1 vccd1 _18422_/A sky130_fd_sc_hd__buf_2
XFILLER_77_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1967 _18905_/A vssd1 vssd1 vccd1 vccd1 _18112_/A sky130_fd_sc_hd__buf_6
XFILLER_78_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout980 _17099_/A1 vssd1 vssd1 vccd1 vccd1 _17692_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1978 _13595_/A vssd1 vssd1 vccd1 vccd1 _18842_/A sky130_fd_sc_hd__clkbuf_8
X_18610_ _18842_/A _18610_/B vssd1 vssd1 vccd1 vccd1 _20925_/D sky130_fd_sc_hd__nor2_1
XFILLER_219_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1989 fanout2002/X vssd1 vssd1 vccd1 vccd1 _17952_/A sky130_fd_sc_hd__buf_8
X_15822_ _15822_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15822_/X sky130_fd_sc_hd__and2_1
Xfanout991 _16964_/B1 vssd1 vssd1 vccd1 vccd1 _16980_/B1 sky130_fd_sc_hd__buf_4
X_19590_ _19590_/CLK _19590_/D vssd1 vssd1 vccd1 vccd1 _19590_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18541_ _18560_/A _18541_/B vssd1 vssd1 vccd1 vccd1 _18541_/X sky130_fd_sc_hd__or2_1
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15753_ _15882_/A1 _15742_/X _15743_/X _15752_/X vssd1 vssd1 vccd1 vccd1 _15753_/X
+ sky130_fd_sc_hd__a22o_4
X_12965_ _14121_/A _14119_/B _14119_/A vssd1 vssd1 vccd1 vccd1 _12965_/X sky130_fd_sc_hd__or3b_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ _16605_/A _17574_/B _14704_/C vssd1 vssd1 vccd1 vccd1 _14704_/X sky130_fd_sc_hd__and3_4
X_11916_ _19292_/Q _20079_/Q _11916_/S vssd1 vssd1 vccd1 vccd1 _11916_/X sky130_fd_sc_hd__mux2_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _18767_/A _18472_/B vssd1 vssd1 vccd1 vccd1 _18472_/X sky130_fd_sc_hd__or2_1
X_15684_ _14815_/S _15547_/X _15548_/Y _16053_/A vssd1 vssd1 vccd1 vccd1 _15684_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12896_ _12896_/A _13209_/A _13221_/A vssd1 vssd1 vccd1 vccd1 _12896_/X sky130_fd_sc_hd__or3b_1
XFILLER_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 _19501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_351 _17917_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _17919_/A _17919_/B _14635_/C vssd1 vssd1 vccd1 vccd1 _14635_/X sky130_fd_sc_hd__and3_4
XANTENNA_362 _10308_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17423_ _20265_/Q _20264_/Q _17446_/A _17423_/D vssd1 vssd1 vccd1 vccd1 _17423_/X
+ sky130_fd_sc_hd__and4_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_373 _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11847_ _19822_/Q _12009_/A2 _11845_/X _12183_/C1 _11846_/X vssd1 vssd1 vccd1 vccd1
+ _11847_/X sky130_fd_sc_hd__o221a_1
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_384 _15338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_395 _15888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _20225_/Q _17356_/A2 _17362_/B1 _20274_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17354_/X sky130_fd_sc_hd__a221o_1
XFILLER_186_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14566_ _17744_/A _17918_/B vssd1 vssd1 vccd1 vccd1 _14567_/C sky130_fd_sc_hd__nor2_1
XFILLER_158_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11319_/X _11778_/B _11778_/C vssd1 vssd1 vccd1 vccd1 _15259_/A sky130_fd_sc_hd__and3b_1
XFILLER_202_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16305_ _19709_/Q _16306_/C _19710_/Q vssd1 vssd1 vccd1 vccd1 _16307_/B sky130_fd_sc_hd__a21oi_1
X_13517_ _13056_/Y _13517_/B vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__nand2b_1
X_17285_ _20200_/Q _17330_/A2 _17291_/B1 _17284_/X vssd1 vssd1 vccd1 vccd1 _17285_/X
+ sky130_fd_sc_hd__a211o_1
X_10729_ _12396_/A1 _19468_/Q _19436_/Q _12397_/S _12371_/C1 vssd1 vssd1 vccd1 vccd1
+ _10729_/X sky130_fd_sc_hd__a221o_1
XFILLER_146_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14497_ _19275_/Q _17894_/A1 _14519_/S vssd1 vssd1 vccd1 vccd1 _19275_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19024_ _18255_/Y _19048_/A2 _18760_/X _12553_/D _19048_/C1 vssd1 vssd1 vccd1 vccd1
+ _19024_/X sky130_fd_sc_hd__a221o_1
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16236_ _16240_/A1 _16235_/X _19695_/D vssd1 vssd1 vccd1 vccd1 _19656_/D sky130_fd_sc_hd__o21a_4
X_13448_ _13448_/A _13448_/B vssd1 vssd1 vccd1 vccd1 _13448_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_103_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap1275 _16066_/A vssd1 vssd1 vccd1 vccd1 _09569_/A sky130_fd_sc_hd__buf_6
X_16167_ _19607_/Q _16170_/S _16166_/Y _16167_/C1 vssd1 vssd1 vccd1 vccd1 _19607_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13379_ _20928_/Q _13602_/A1 _18612_/B vssd1 vssd1 vccd1 vccd1 _13379_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15118_ _15109_/X _15117_/X _15118_/S vssd1 vssd1 vccd1 vccd1 _15983_/B sky130_fd_sc_hd__mux2_4
XFILLER_114_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16098_ _10282_/X _16126_/A2 _16097_/X vssd1 vssd1 vccd1 vccd1 _19573_/D sky130_fd_sc_hd__o21a_1
XFILLER_141_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19926_ _20662_/CLK _19926_/D vssd1 vssd1 vccd1 vccd1 _19926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15049_ _15045_/X _15048_/X _15292_/S vssd1 vssd1 vccd1 vccd1 _15049_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20692_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_268_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19857_ _20017_/CLK _19857_/D vssd1 vssd1 vccd1 vccd1 _19857_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_205_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09610_ _09610_/A _12967_/B _09610_/C vssd1 vssd1 vccd1 vccd1 _09686_/C sky130_fd_sc_hd__and3_2
XFILLER_284_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18808_ _18808_/A _18808_/B vssd1 vssd1 vccd1 vccd1 _20986_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19788_ _20451_/CLK _19788_/D vssd1 vssd1 vccd1 vccd1 _19788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09541_ _12480_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _09541_/Y sky130_fd_sc_hd__nand2_4
X_18739_ _20970_/Q _18280_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18740_/B sky130_fd_sc_hd__mux2_1
XFILLER_271_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20701_ _20701_/CLK _20701_/D vssd1 vssd1 vccd1 vccd1 _20701_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20632_ _20655_/CLK _20632_/D vssd1 vssd1 vccd1 vccd1 _20632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20563_ _20563_/CLK _20563_/D vssd1 vssd1 vccd1 vccd1 _20563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20494_ _20659_/CLK _20494_/D vssd1 vssd1 vccd1 vccd1 _20494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1208 _15095_/X vssd1 vssd1 vccd1 vccd1 _16002_/B1 sky130_fd_sc_hd__buf_6
XFILLER_266_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1219 _13370_/B vssd1 vssd1 vccd1 vccd1 _13397_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_59_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21046_ _21046_/A vssd1 vssd1 vccd1 vccd1 _21046_/X sky130_fd_sc_hd__buf_2
XFILLER_115_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09808_ _09806_/X _09807_/X _12058_/S vssd1 vssd1 vccd1 vccd1 _09808_/X sky130_fd_sc_hd__mux2_1
XFILLER_274_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_15__f_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_15__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09739_ _11291_/A2 _12258_/S _11204_/S _11396_/S vssd1 vssd1 vccd1 vccd1 _09748_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12750_ _12791_/A _12791_/B vssd1 vssd1 vccd1 vccd1 _12750_/Y sky130_fd_sc_hd__nor2_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11701_ _09834_/A _20543_/Q _20511_/Q _10621_/S vssd1 vssd1 vccd1 vccd1 _11701_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12681_ _12479_/A _12582_/C _12682_/B _12680_/Y vssd1 vssd1 vccd1 vccd1 _12681_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _19244_/Q _14438_/A2 _14419_/X _16187_/A vssd1 vssd1 vccd1 vccd1 _19244_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _19417_/Q _12025_/S _11631_/X _09834_/C vssd1 vssd1 vccd1 vccd1 _11632_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ _19517_/Q _14352_/B vssd1 vssd1 vccd1 vccd1 _14361_/A sky130_fd_sc_hd__and2_1
XFILLER_129_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11563_ _11561_/X _11562_/X _11563_/S vssd1 vssd1 vccd1 vccd1 _11563_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13302_ _13334_/A _13300_/X _13301_/Y _13298_/X vssd1 vssd1 vccd1 vccd1 _13302_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10514_ _19672_/Q _20160_/Q _11295_/S vssd1 vssd1 vccd1 vccd1 _10514_/X sky130_fd_sc_hd__mux2_1
X_17070_ _20042_/Q _17872_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20042_/D sky130_fd_sc_hd__mux2_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14282_ _14280_/Y _14282_/B vssd1 vssd1 vccd1 vccd1 _14283_/B sky130_fd_sc_hd__and2b_1
X_11494_ _11495_/A _11734_/B vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__or2_2
X_16021_ _16049_/A1 _16010_/X _16020_/X vssd1 vssd1 vccd1 vccd1 _16021_/X sky130_fd_sc_hd__a21o_4
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ _13233_/A _13233_/B _13233_/C vssd1 vssd1 vccd1 vccd1 _13233_/X sky130_fd_sc_hd__or3_1
X_10445_ _19809_/Q _10502_/A2 _10443_/X _11274_/B2 _10444_/X vssd1 vssd1 vccd1 vccd1
+ _10445_/X sky130_fd_sc_hd__o221a_1
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ _11497_/A _13162_/A _13162_/B _11730_/B _11496_/Y vssd1 vssd1 vccd1 vccd1
+ _13166_/C sky130_fd_sc_hd__a311o_1
X_10376_ _19578_/Q _10375_/X _11243_/S vssd1 vssd1 vccd1 vccd1 _10377_/B sky130_fd_sc_hd__mux2_2
XFILLER_151_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12115_ _11955_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12115_/X sky130_fd_sc_hd__and2b_1
XFILLER_69_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17972_ _18064_/A _17972_/B _17976_/C vssd1 vssd1 vccd1 vccd1 _20728_/D sky130_fd_sc_hd__nor3_1
X_13095_ _20911_/Q _13092_/X _13094_/Y vssd1 vssd1 vccd1 vccd1 _13096_/B sky130_fd_sc_hd__o21a_1
XFILLER_269_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19711_ _20757_/CLK _19711_/D vssd1 vssd1 vccd1 vccd1 _19711_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1720 _12138_/A1 vssd1 vssd1 vccd1 vccd1 _11983_/A1 sky130_fd_sc_hd__buf_8
X_12046_ _10430_/S _12051_/A1 _19360_/Q _12046_/B1 vssd1 vssd1 vccd1 vccd1 _12046_/X
+ sky130_fd_sc_hd__a31o_1
X_16923_ _16981_/A1 _15780_/X _16879_/X _16922_/X vssd1 vssd1 vccd1 vccd1 _16923_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1731 _12312_/A1 vssd1 vssd1 vccd1 vccd1 _12396_/A1 sky130_fd_sc_hd__buf_6
XFILLER_284_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1742 _12519_/C vssd1 vssd1 vccd1 vccd1 _09695_/A sky130_fd_sc_hd__buf_8
XFILLER_266_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1753 _13967_/S vssd1 vssd1 vccd1 vccd1 _14003_/S sky130_fd_sc_hd__buf_8
XFILLER_238_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1764 _14524_/A1 vssd1 vssd1 vccd1 vccd1 _13582_/A sky130_fd_sc_hd__buf_4
X_19642_ _20480_/CLK _19642_/D vssd1 vssd1 vccd1 vccd1 _19642_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1775 output482/A vssd1 vssd1 vccd1 vccd1 _18152_/B sky130_fd_sc_hd__buf_4
X_16854_ _16805_/X _16851_/Y _16853_/X _17008_/A1 vssd1 vssd1 vccd1 vccd1 _16854_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout1786 _18223_/B vssd1 vssd1 vccd1 vccd1 _18248_/B sky130_fd_sc_hd__buf_12
Xfanout1797 _12548_/B vssd1 vssd1 vccd1 vccd1 _12549_/B sky130_fd_sc_hd__buf_4
XFILLER_266_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15805_ _20808_/Q _15941_/A2 _15798_/X _15941_/B2 _15804_/X vssd1 vssd1 vccd1 vccd1
+ _15805_/X sky130_fd_sc_hd__a221o_2
X_19573_ _19574_/CLK _19573_/D vssd1 vssd1 vccd1 vccd1 _19573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13997_ _19198_/Q _14077_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _13997_/X sky130_fd_sc_hd__mux2_1
X_16785_ _20403_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16785_/X sky130_fd_sc_hd__a21o_1
XFILLER_253_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18524_ _20901_/Q _18559_/B _18523_/X _18458_/B vssd1 vssd1 vccd1 vccd1 _18525_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12948_ _20012_/Q _20013_/Q _20014_/Q vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__or3_4
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15736_ _16053_/A _15736_/B vssd1 vssd1 vccd1 vccd1 _15736_/Y sky130_fd_sc_hd__nor2_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_162_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20998_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_261_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18455_ _13479_/A _13478_/A _12589_/C _18472_/B _14110_/A vssd1 vssd1 vccd1 vccd1
+ _18455_/X sky130_fd_sc_hd__o311a_1
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12879_ _19521_/Q _12889_/A vssd1 vssd1 vccd1 vccd1 _12880_/B sky130_fd_sc_hd__nor2_1
XANTENNA_170 _19108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15667_ _20963_/Q _15939_/A2 _15996_/B1 _20835_/Q _15666_/X vssd1 vssd1 vccd1 vccd1
+ _15667_/X sky130_fd_sc_hd__a221o_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_192 _19541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17406_ _17402_/A _17441_/A _17457_/B _20251_/Q vssd1 vssd1 vccd1 vccd1 _17406_/X
+ sky130_fd_sc_hd__a31o_1
X_14618_ _19382_/Q _17902_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19382_/D sky130_fd_sc_hd__mux2_1
X_18386_ _20848_/Q _18385_/B _18385_/Y _18734_/A vssd1 vssd1 vccd1 vccd1 _20848_/D
+ sky130_fd_sc_hd__o211a_1
X_15598_ _20897_/Q _15937_/A2 _15994_/B1 _15597_/X _15937_/C1 vssd1 vssd1 vccd1 vccd1
+ _15598_/X sky130_fd_sc_hd__a221o_1
XFILLER_159_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14549_ _19319_/Q _17592_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19319_/D sky130_fd_sc_hd__mux2_1
X_17337_ _17337_/A _17337_/B vssd1 vssd1 vccd1 vccd1 _17337_/Y sky130_fd_sc_hd__nor2_8
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17268_ _20195_/Q _17268_/A2 _17266_/X _17267_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1
+ _20195_/D sky130_fd_sc_hd__o221a_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19007_ _21023_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _19007_/X sky130_fd_sc_hd__or2_1
X_16219_ _19642_/Q _17696_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19642_/D sky130_fd_sc_hd__mux2_1
X_17199_ _20163_/Q _17199_/A1 _17215_/S vssd1 vssd1 vccd1 vccd1 _20163_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19909_ _20669_/CLK _19909_/D vssd1 vssd1 vccd1 vccd1 _19909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09524_ input45/X vssd1 vssd1 vccd1 vccd1 _09524_/Y sky130_fd_sc_hd__inv_2
XFILLER_271_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20615_ _20683_/CLK _20615_/D vssd1 vssd1 vccd1 vccd1 _20615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20546_ _20646_/CLK _20546_/D vssd1 vssd1 vccd1 vccd1 _20546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20477_ _20573_/CLK _20477_/D vssd1 vssd1 vccd1 vccd1 _20477_/Q sky130_fd_sc_hd__dfxtp_1
X_10230_ _19381_/Q _20672_/Q _10983_/S vssd1 vssd1 vccd1 vccd1 _10230_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10161_ _09689_/A _10153_/X _10160_/X _10144_/X vssd1 vssd1 vccd1 vccd1 _10161_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput380 _13804_/X vssd1 vssd1 vccd1 vccd1 din0[13] sky130_fd_sc_hd__buf_4
Xfanout1005 _16049_/A1 vssd1 vssd1 vccd1 vccd1 _15606_/A1 sky130_fd_sc_hd__buf_12
Xoutput391 _13814_/X vssd1 vssd1 vccd1 vccd1 din0[23] sky130_fd_sc_hd__buf_4
XFILLER_273_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1016 _18974_/A2 vssd1 vssd1 vccd1 vccd1 _18954_/A2 sky130_fd_sc_hd__buf_4
XFILLER_117_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1027 _16963_/A2 vssd1 vssd1 vccd1 vccd1 _17004_/A2 sky130_fd_sc_hd__buf_6
XFILLER_248_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1038 _11247_/X vssd1 vssd1 vccd1 vccd1 _17852_/A1 sky130_fd_sc_hd__buf_4
XFILLER_102_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _20130_/Q _20098_/Q _10092_/S vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__mux2_1
XFILLER_266_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1049 _11049_/B1 vssd1 vssd1 vccd1 vccd1 _17889_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13920_ _18710_/A _13920_/B vssd1 vssd1 vccd1 vccd1 _19125_/D sky130_fd_sc_hd__and2_1
X_21029_ _21029_/CLK _21029_/D vssd1 vssd1 vccd1 vccd1 _21029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ _13847_/X _20249_/Q _17335_/B vssd1 vssd1 vccd1 vccd1 _13851_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ _19515_/Q _12916_/A2 _12801_/X _12916_/B2 vssd1 vssd1 vccd1 vccd1 _12803_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16570_ _19851_/Q _16592_/A2 _16592_/B1 input22/X vssd1 vssd1 vccd1 vccd1 _16571_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_76_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13782_ split3/X _13497_/Y _13509_/Y _16240_/A1 vssd1 vssd1 vccd1 vccd1 _13782_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_222_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10994_ _10989_/X _10993_/X _09621_/A vssd1 vssd1 vccd1 vccd1 _10994_/X sky130_fd_sc_hd__a21o_1
XFILLER_16_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15521_ _12578_/B _12729_/X _15589_/S vssd1 vssd1 vccd1 vccd1 _15521_/Y sky130_fd_sc_hd__o21ai_1
X_12733_ _19506_/Q _12758_/B vssd1 vssd1 vccd1 vccd1 _12736_/C sky130_fd_sc_hd__nand2_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15452_ _17269_/A _15451_/X _15452_/S vssd1 vssd1 vccd1 vccd1 _15452_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18240_ _18514_/B vssd1 vssd1 vccd1 vccd1 _18240_/Y sky130_fd_sc_hd__inv_2
X_12664_ _19496_/Q _19495_/Q _12664_/C vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__nor3_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _19521_/Q _14392_/B _14394_/B vssd1 vssd1 vccd1 vccd1 _14403_/X sky130_fd_sc_hd__a21o_1
X_11615_ _12828_/A _11649_/S _11614_/Y vssd1 vssd1 vccd1 vccd1 _11651_/A sky130_fd_sc_hd__o21a_1
XFILLER_89_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18171_ _20788_/Q _18170_/Y _18236_/S vssd1 vssd1 vccd1 vccd1 _18172_/B sky130_fd_sc_hd__mux2_1
X_15383_ _20858_/Q _15569_/S vssd1 vssd1 vccd1 vccd1 _15383_/X sky130_fd_sc_hd__or2_1
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12595_ _12708_/A _13002_/A vssd1 vssd1 vccd1 vccd1 _12917_/A sky130_fd_sc_hd__nand2_2
XFILLER_204_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17122_ _20090_/Q _17647_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20090_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14334_ _14333_/A _14333_/B _14333_/C vssd1 vssd1 vccd1 vccd1 _14343_/B sky130_fd_sc_hd__a21o_1
XFILLER_184_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11546_ _09986_/A _20541_/Q _20509_/Q _12174_/S vssd1 vssd1 vccd1 vccd1 _11546_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17053_ _20025_/Q _17855_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20025_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14265_ _14397_/A _14397_/B _14265_/C vssd1 vssd1 vccd1 vccd1 _14265_/X sky130_fd_sc_hd__or3_1
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11477_ _12186_/S _11477_/B vssd1 vssd1 vccd1 vccd1 _11477_/X sky130_fd_sc_hd__or2_1
X_16004_ _15526_/B _15987_/X _16003_/X _15526_/Y vssd1 vssd1 vccd1 vccd1 _16004_/X
+ sky130_fd_sc_hd__a22o_1
X_13216_ _13216_/A _13272_/B vssd1 vssd1 vccd1 vccd1 _13216_/Y sky130_fd_sc_hd__nor2_1
X_10428_ _19876_/Q _19777_/Q _10428_/S vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14196_ _20274_/Q _14237_/A2 _14216_/B1 input245/X vssd1 vssd1 vccd1 vccd1 _14198_/B
+ sky130_fd_sc_hd__a22o_4
X_13147_ _15226_/A _13523_/B _10968_/Y vssd1 vssd1 vccd1 vccd1 _13538_/B sky130_fd_sc_hd__a21o_4
XFILLER_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10359_ _10357_/X _10358_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _10359_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _18048_/A _17955_/B _17959_/C vssd1 vssd1 vccd1 vccd1 _20722_/D sky130_fd_sc_hd__nor3_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13029_/Y _13327_/A _13326_/B vssd1 vssd1 vccd1 vccd1 _13303_/C sky130_fd_sc_hd__o21ai_4
XFILLER_39_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1550 fanout1556/X vssd1 vssd1 vccd1 vccd1 _11074_/S sky130_fd_sc_hd__buf_4
XFILLER_211_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12029_ _12192_/A1 _12012_/X _12020_/X _12028_/Y vssd1 vssd1 vccd1 vccd1 _12029_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_16906_ _19234_/Q _16980_/A2 _16980_/B1 _19103_/Q _16905_/X vssd1 vssd1 vccd1 vccd1
+ _16906_/X sky130_fd_sc_hd__o221a_1
Xfanout1561 _10842_/S vssd1 vssd1 vccd1 vccd1 _12323_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_272_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17886_ _20657_/Q _17886_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20657_/D sky130_fd_sc_hd__mux2_1
Xfanout1572 _09624_/Y vssd1 vssd1 vccd1 vccd1 _12072_/C1 sky130_fd_sc_hd__buf_4
XFILLER_254_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1583 _11009_/B2 vssd1 vssd1 vccd1 vccd1 _11353_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19625_ _20463_/CLK _19625_/D vssd1 vssd1 vccd1 vccd1 _19625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1594 _11008_/A3 vssd1 vssd1 vccd1 vccd1 _11363_/A1 sky130_fd_sc_hd__clkbuf_8
X_16837_ _16846_/A input80/X vssd1 vssd1 vccd1 vccd1 _16837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19556_ _19618_/CLK _19556_/D vssd1 vssd1 vccd1 vccd1 _19556_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_280_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16768_ _17008_/A1 _16767_/X _17008_/B1 vssd1 vssd1 vccd1 vccd1 _16768_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_213_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18507_ _18891_/A _18507_/B vssd1 vssd1 vccd1 vccd1 _20895_/D sky130_fd_sc_hd__nor2_1
XFILLER_280_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15719_ _20901_/Q _15322_/A _15994_/B1 _15718_/X _15323_/A vssd1 vssd1 vccd1 vccd1
+ _15719_/X sky130_fd_sc_hd__a221o_1
XFILLER_280_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19487_ _20708_/CLK _19487_/D vssd1 vssd1 vccd1 vccd1 _19487_/Q sky130_fd_sc_hd__dfxtp_1
X_16699_ _19954_/Q _17945_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19954_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18438_ _18734_/A _18438_/B vssd1 vssd1 vccd1 vccd1 _20873_/D sky130_fd_sc_hd__and2_1
XFILLER_178_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18369_ _18532_/B _18385_/B vssd1 vssd1 vccd1 vccd1 _18369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20400_ _20690_/CLK _20400_/D vssd1 vssd1 vccd1 vccd1 _20400_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20331_ _20468_/CLK _20331_/D vssd1 vssd1 vccd1 vccd1 _20331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20262_ _20421_/CLK _20262_/D vssd1 vssd1 vccd1 vccd1 _20262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20193_ _20727_/CLK _20193_/D vssd1 vssd1 vccd1 vccd1 _20193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput108 dout1[10] vssd1 vssd1 vccd1 vccd1 input108/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput119 dout1[20] vssd1 vssd1 vccd1 vccd1 input119/X sky130_fd_sc_hd__clkbuf_2
XFILLER_243_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09507_ _09507_/A vssd1 vssd1 vccd1 vccd1 _09507_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11400_ _11400_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11401_/B sky130_fd_sc_hd__nor2_1
XFILLER_184_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12380_ _20491_/Q _20331_/Q _12381_/S vssd1 vssd1 vccd1 vccd1 _12380_/X sky130_fd_sc_hd__mux2_1
XANTENNA_70 _09504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_81 _09869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _19535_/Q _09594_/X _11325_/X _11330_/Y vssd1 vssd1 vccd1 vccd1 _11331_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_92 _12035_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20529_ _20690_/CLK _20529_/D vssd1 vssd1 vccd1 vccd1 _20529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14050_ _19184_/Q _14082_/A2 _14049_/X _16195_/A vssd1 vssd1 vccd1 vccd1 _19184_/D
+ sky130_fd_sc_hd__o211a_1
X_11262_ _20625_/Q _09688_/B _11261_/X _11274_/B2 vssd1 vssd1 vccd1 vccd1 _11262_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ _19246_/Q _13001_/B vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__xnor2_1
X_10213_ _19477_/Q _09695_/Y _10212_/X _12377_/S vssd1 vssd1 vccd1 vccd1 _10213_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_137_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11193_ _19624_/Q _19930_/Q _19268_/Q _20055_/Q _12346_/S _11391_/C vssd1 vssd1 vccd1
+ vccd1 _11193_/X sky130_fd_sc_hd__mux4_1
XFILLER_133_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10144_ _11101_/A _10142_/X _10143_/X _12311_/C1 vssd1 vssd1 vccd1 vccd1 _10144_/X
+ sky130_fd_sc_hd__a211o_2
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ _20521_/Q _17914_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20521_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14952_ _14958_/A _14973_/B _14966_/C vssd1 vssd1 vccd1 vccd1 _15020_/A sky130_fd_sc_hd__or3_4
XFILLER_153_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10075_ _12073_/C1 _10058_/X _10074_/X _12074_/B1 vssd1 vssd1 vccd1 vccd1 _10075_/X
+ sky130_fd_sc_hd__a211o_2
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13903_ _16241_/A _13943_/S vssd1 vssd1 vccd1 vccd1 _13903_/Y sky130_fd_sc_hd__nor2_4
X_17671_ _20457_/Q _17705_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20457_/D sky130_fd_sc_hd__mux2_1
X_14883_ _14885_/B vssd1 vssd1 vccd1 vccd1 _14883_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19410_ _20701_/CLK _19410_/D vssd1 vssd1 vccd1 vccd1 _19410_/Q sky130_fd_sc_hd__dfxtp_1
X_16622_ _19881_/Q _17936_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19881_/D sky130_fd_sc_hd__mux2_1
XFILLER_235_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13834_ _20004_/Q split1/X _13788_/X split2/X vssd1 vssd1 vccd1 vccd1 _13834_/X sky130_fd_sc_hd__a22o_4
XFILLER_251_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19341_ _20719_/CLK _19341_/D vssd1 vssd1 vccd1 vccd1 _19341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16553_ _16593_/A _16553_/B vssd1 vssd1 vccd1 vccd1 _19842_/D sky130_fd_sc_hd__or2_1
XFILLER_188_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _13765_/A _13765_/B vssd1 vssd1 vccd1 vccd1 _13765_/X sky130_fd_sc_hd__and2_2
XFILLER_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10977_ _19562_/Q _11061_/A _09659_/X _10976_/Y vssd1 vssd1 vccd1 vccd1 _10977_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15504_ _15504_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _15504_/Y sky130_fd_sc_hd__nand2_1
X_19272_ _20085_/CLK _19272_/D vssd1 vssd1 vccd1 vccd1 _19272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12716_ _14894_/A _12716_/B vssd1 vssd1 vccd1 vccd1 _12716_/Y sky130_fd_sc_hd__nand2_1
XFILLER_280_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13696_ _13697_/B vssd1 vssd1 vccd1 vccd1 _13696_/Y sky130_fd_sc_hd__inv_2
X_16484_ _19793_/Q _17947_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19793_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18223_ _19540_/Q _18223_/B vssd1 vssd1 vccd1 vccd1 _18223_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_188_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12647_ _12647_/A _12647_/B vssd1 vssd1 vccd1 vccd1 _12647_/X sky130_fd_sc_hd__or2_1
X_15435_ _15108_/X _15112_/X _15577_/S vssd1 vssd1 vccd1 vccd1 _15435_/X sky130_fd_sc_hd__mux2_1
XFILLER_248_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18154_ _18323_/B _18154_/B vssd1 vssd1 vccd1 vccd1 _18390_/A sky130_fd_sc_hd__nand2_2
X_15366_ _15326_/A _15351_/Y _15365_/X _15349_/X vssd1 vssd1 vccd1 vccd1 _15366_/X
+ sky130_fd_sc_hd__o31a_1
X_12578_ _12578_/A _12578_/B _15326_/A vssd1 vssd1 vccd1 vccd1 _14809_/A sky130_fd_sc_hd__and3_1
XFILLER_200_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17105_ _20075_/Q _17835_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20075_/D sky130_fd_sc_hd__mux2_1
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11529_ _12140_/C1 _11528_/X _11525_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _11529_/X
+ sky130_fd_sc_hd__o211a_1
X_14317_ _13373_/A _14316_/X _13307_/Y vssd1 vssd1 vccd1 vccd1 _14318_/C sky130_fd_sc_hd__o21a_1
X_18085_ _20769_/Q _20768_/Q _18085_/C vssd1 vssd1 vccd1 vccd1 _18087_/B sky130_fd_sc_hd__and3_1
XFILLER_172_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15297_ _15297_/A vssd1 vssd1 vccd1 vccd1 _15297_/Y sky130_fd_sc_hd__inv_2
X_17036_ _20014_/Q input200/X _17038_/S vssd1 vssd1 vccd1 vccd1 _20014_/D sky130_fd_sc_hd__mux2_1
X_14248_ _19507_/Q _14249_/B vssd1 vssd1 vccd1 vccd1 _14260_/A sky130_fd_sc_hd__nand2_1
XFILLER_259_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ _19499_/Q _14171_/B _14170_/B vssd1 vssd1 vccd1 vccd1 _14179_/X sky130_fd_sc_hd__o21a_1
XFILLER_171_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 _18864_/B1 vssd1 vssd1 vccd1 vccd1 _18974_/B1 sky130_fd_sc_hd__buf_2
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18987_ _21013_/Q _18997_/B vssd1 vssd1 vccd1 vccd1 _18987_/X sky130_fd_sc_hd__or2_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _20707_/Q _17938_/A1 _17946_/S vssd1 vssd1 vccd1 vccd1 _20707_/D sky130_fd_sc_hd__mux2_1
XFILLER_239_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1380 _11860_/B2 vssd1 vssd1 vccd1 vccd1 _11947_/S sky130_fd_sc_hd__buf_6
Xfanout1391 _11848_/S0 vssd1 vssd1 vccd1 vccd1 _12165_/S sky130_fd_sc_hd__buf_6
XFILLER_254_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17869_ _20642_/Q _17869_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20642_/D sky130_fd_sc_hd__mux2_1
XFILLER_213_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19608_ _19609_/CLK _19608_/D vssd1 vssd1 vccd1 vccd1 _19608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20880_ _21000_/CLK _20880_/D vssd1 vssd1 vccd1 vccd1 _20880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19539_ _19541_/CLK _19539_/D vssd1 vssd1 vccd1 vccd1 _19539_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_241_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20314_ _20692_/CLK _20314_/D vssd1 vssd1 vccd1 vccd1 _20314_/Q sky130_fd_sc_hd__dfxtp_1
Xinput90 dout0[52] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20245_ _20296_/CLK _20245_/D vssd1 vssd1 vccd1 vccd1 _20245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ _19818_/Q _12009_/A2 _09985_/X _11563_/S _09986_/X vssd1 vssd1 vccd1 vccd1
+ _09987_/X sky130_fd_sc_hd__o221a_1
XFILLER_27_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20176_ _20715_/CLK _20176_/D vssd1 vssd1 vccd1 vccd1 _20176_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10900_ _11266_/A1 _20661_/Q _11270_/A2 _11256_/S vssd1 vssd1 vccd1 vccd1 _10900_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11880_ _11880_/A _11880_/B vssd1 vssd1 vccd1 vccd1 _11883_/D sky130_fd_sc_hd__xnor2_2
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ _10829_/X _10830_/X _10831_/S vssd1 vssd1 vccd1 vccd1 _10831_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ _13064_/X _13564_/B _13549_/Y _18760_/B vssd1 vssd1 vccd1 vccd1 _13550_/X
+ sky130_fd_sc_hd__o31a_1
X_10762_ _12245_/A1 _17926_/A1 _12401_/B1 vssd1 vssd1 vccd1 vccd1 _10762_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12501_ _19160_/Q _19159_/Q _19158_/Q _19157_/Q vssd1 vssd1 vccd1 vccd1 _12502_/C
+ sky130_fd_sc_hd__or4_1
X_13481_ _13481_/A _17041_/B vssd1 vssd1 vccd1 vccd1 _16598_/C sky130_fd_sc_hd__or2_4
X_10693_ _19373_/Q _12412_/A2 _10691_/X _12412_/B2 _10692_/X vssd1 vssd1 vccd1 vccd1
+ _10693_/X sky130_fd_sc_hd__o221a_1
XFILLER_13_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15220_ _15220_/A _15220_/B vssd1 vssd1 vccd1 vccd1 _15220_/X sky130_fd_sc_hd__or2_4
X_12432_ _12423_/X _12431_/Y _11201_/A _12415_/X vssd1 vssd1 vccd1 vccd1 _12432_/X
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_157_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15151_ _16133_/C _15148_/Y _15149_/X _15150_/X vssd1 vssd1 vccd1 vccd1 _15151_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12363_ _12440_/A _14882_/A vssd1 vssd1 vccd1 vccd1 _12449_/A sky130_fd_sc_hd__or2_2
XFILLER_193_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _19210_/Q _14106_/A2 _14101_/X _16129_/B1 vssd1 vssd1 vccd1 vccd1 _19210_/D
+ sky130_fd_sc_hd__o211a_1
X_11314_ _11313_/B _11312_/X _11313_/Y vssd1 vssd1 vccd1 vccd1 _11783_/B sky130_fd_sc_hd__o21ai_4
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15082_ _21013_/Q _20981_/Q _15309_/S vssd1 vssd1 vccd1 vccd1 _15082_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12294_ _20556_/Q _12313_/S vssd1 vssd1 vccd1 vccd1 _12294_/X sky130_fd_sc_hd__or2_1
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14033_ _19210_/Q _14101_/C _14039_/S vssd1 vssd1 vccd1 vccd1 _14033_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18910_ _21001_/Q _18971_/B vssd1 vssd1 vccd1 vccd1 _18910_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11245_ _15103_/A1 _11240_/X _11244_/X vssd1 vssd1 vccd1 vccd1 _11245_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19890_ _20077_/CLK _19890_/D vssd1 vssd1 vccd1 vccd1 _19890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18841_ _18499_/X _18840_/B _18839_/X _18840_/Y vssd1 vssd1 vccd1 vccd1 _18842_/B
+ sky130_fd_sc_hd__o211a_1
X_11176_ _09618_/A _11174_/X _11175_/X _09621_/A vssd1 vssd1 vccd1 vccd1 _11176_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_268_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10127_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10127_/Y sky130_fd_sc_hd__nand2_2
X_18772_ _18808_/A _18772_/B vssd1 vssd1 vccd1 vccd1 _20980_/D sky130_fd_sc_hd__nor2_1
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15984_ _12283_/B _15984_/A2 _15984_/B1 _12281_/Y _16030_/D1 vssd1 vssd1 vccd1 vccd1
+ _15984_/X sky130_fd_sc_hd__a221o_1
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17723_ _20504_/Q split4/A _17738_/S vssd1 vssd1 vccd1 vccd1 _20504_/D sky130_fd_sc_hd__mux2_1
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14935_ _15314_/C _14948_/A vssd1 vssd1 vccd1 vccd1 _14935_/Y sky130_fd_sc_hd__nor2_8
XFILLER_236_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10058_ _10048_/X _10051_/X _10054_/X _10057_/X _12058_/S _12059_/A1 vssd1 vssd1
+ vccd1 vccd1 _10058_/X sky130_fd_sc_hd__mux4_2
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17654_ _20440_/Q _17931_/A1 _17669_/S vssd1 vssd1 vccd1 vccd1 _20440_/D sky130_fd_sc_hd__mux2_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ _11223_/B _12443_/B _14870_/S vssd1 vssd1 vccd1 vccd1 _15039_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16605_ _16605_/A _17574_/B _16605_/C vssd1 vssd1 vccd1 vccd1 _16605_/X sky130_fd_sc_hd__and3_4
XFILLER_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13817_ _13822_/A1 _13755_/B split9/A input233/X vssd1 vssd1 vccd1 vccd1 _13817_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17585_ _20343_/Q _17896_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20343_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14797_ _19523_/Q _14797_/B vssd1 vssd1 vccd1 vccd1 _14797_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_69_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20658_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19324_ _20479_/CLK _19324_/D vssd1 vssd1 vccd1 vccd1 _19324_/Q sky130_fd_sc_hd__dfxtp_1
X_16536_ _19834_/Q _16578_/A2 _16578_/B1 input35/X vssd1 vssd1 vccd1 vccd1 _16537_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13748_ _13670_/Y _13741_/B _13741_/Y _13671_/Y _13747_/X vssd1 vssd1 vccd1 vccd1
+ _13749_/B sky130_fd_sc_hd__o221a_4
XFILLER_232_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19255_ _20273_/CLK _19255_/D vssd1 vssd1 vccd1 vccd1 _19255_/Q sky130_fd_sc_hd__dfxtp_1
X_16467_ _19776_/Q _17930_/A1 _16471_/S vssd1 vssd1 vccd1 vccd1 _19776_/D sky130_fd_sc_hd__mux2_1
X_13679_ _16598_/C _13679_/B vssd1 vssd1 vccd1 vccd1 _13679_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18206_ _20795_/Q _18205_/Y _18236_/S vssd1 vssd1 vccd1 vccd1 _18207_/B sky130_fd_sc_hd__mux2_1
X_15418_ _20923_/Q _15567_/A2 _15417_/X vssd1 vssd1 vccd1 vccd1 _15418_/X sky130_fd_sc_hd__o21a_1
X_19186_ _21044_/CLK _19186_/D vssd1 vssd1 vccd1 vccd1 _19186_/Q sky130_fd_sc_hd__dfxtp_1
X_16398_ _19744_/Q _16396_/B _16397_/Y vssd1 vssd1 vccd1 vccd1 _19744_/D sky130_fd_sc_hd__o21a_1
XFILLER_191_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18137_ _18134_/A _18152_/B _18152_/C _18136_/Y vssd1 vssd1 vccd1 vccd1 _18138_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15349_ _12578_/A _13568_/A _15348_/X _10935_/B vssd1 vssd1 vccd1 vccd1 _15349_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18068_ _20762_/Q _18069_/C _20763_/Q vssd1 vssd1 vccd1 vccd1 _18070_/B sky130_fd_sc_hd__a21oi_1
XFILLER_145_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17019_ _19997_/Q input206/X _17849_/S vssd1 vssd1 vccd1 vccd1 _19997_/D sky130_fd_sc_hd__mux2_1
X_09910_ _19819_/Q _12009_/A2 _09908_/X _12183_/C1 _09909_/X vssd1 vssd1 vccd1 vccd1
+ _09910_/X sky130_fd_sc_hd__o221a_1
XFILLER_259_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout606 _14601_/X vssd1 vssd1 vccd1 vccd1 _14632_/S sky130_fd_sc_hd__buf_6
X_20030_ _20658_/CLK _20030_/D vssd1 vssd1 vccd1 vccd1 _20030_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout617 _14488_/X vssd1 vssd1 vccd1 vccd1 _14520_/S sky130_fd_sc_hd__buf_12
X_09841_ _19684_/Q _20172_/Q _10400_/S vssd1 vssd1 vccd1 vccd1 _09841_/X sky130_fd_sc_hd__mux2_1
Xfanout628 _13902_/Y vssd1 vssd1 vccd1 vccd1 _14004_/B1 sky130_fd_sc_hd__buf_6
Xfanout639 _16707_/X vssd1 vssd1 vccd1 vccd1 _16876_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_59_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09772_ _09770_/X _09771_/X _11945_/S vssd1 vssd1 vccd1 vccd1 _09772_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20932_ _20998_/CLK _20932_/D vssd1 vssd1 vccd1 vccd1 _20932_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20863_ _20863_/CLK _20863_/D vssd1 vssd1 vccd1 vccd1 _20863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20794_ _20794_/CLK _20794_/D vssd1 vssd1 vccd1 vccd1 _20794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11030_ _11024_/X _11029_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _11030_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20228_ _21013_/CLK _20228_/D vssd1 vssd1 vccd1 vccd1 _20228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_249_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20159_ _20679_/CLK _20159_/D vssd1 vssd1 vccd1 vccd1 _20159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _13140_/B vssd1 vssd1 vccd1 vccd1 _13902_/A sky130_fd_sc_hd__clkinv_2
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14720_ _19477_/Q _17692_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19477_/D sky130_fd_sc_hd__mux2_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11932_ _20422_/Q _20358_/Q _20650_/Q _20614_/Q _11932_/S0 _12008_/C vssd1 vssd1
+ vccd1 vccd1 _11932_/X sky130_fd_sc_hd__mux4_1
XFILLER_233_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_500 _20004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_511 input218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_522 _13627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14651_ _19413_/Q _17935_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19413_/D sky130_fd_sc_hd__mux2_1
XANTENNA_533 _13637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _11949_/S _11858_/X _11862_/Y _12020_/C1 vssd1 vssd1 vccd1 vccd1 _11872_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_544 _11537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_555 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _20466_/Q _20306_/Q _12389_/S vssd1 vssd1 vccd1 vccd1 _10814_/X sky130_fd_sc_hd__mux2_1
XFILLER_214_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_566 _13472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13602_ _13602_/A1 _13449_/B _13599_/Y _12982_/B vssd1 vssd1 vccd1 vccd1 _13603_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_577 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17370_ _20233_/Q _17378_/A2 _17370_/B1 _20282_/Q _17370_/C1 vssd1 vssd1 vccd1 vccd1
+ _17370_/X sky130_fd_sc_hd__a221o_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_588 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14582_ _19348_/Q _17934_/A1 _14599_/S vssd1 vssd1 vccd1 vccd1 _19348_/D sky130_fd_sc_hd__mux2_1
X_11794_ _13420_/A _11794_/B _11794_/C vssd1 vssd1 vccd1 vccd1 _15652_/B sky130_fd_sc_hd__nand3_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_599 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16321_ _19715_/Q _16322_/C _19716_/Q vssd1 vssd1 vccd1 vccd1 _16323_/B sky130_fd_sc_hd__a21oi_1
X_10745_ _12383_/A _10731_/Y _09502_/A vssd1 vssd1 vccd1 vccd1 _10745_/Y sky130_fd_sc_hd__a21oi_1
X_13533_ _13064_/C _13055_/Y _13062_/Y _13564_/B vssd1 vssd1 vccd1 vccd1 _13533_/X
+ sky130_fd_sc_hd__a31o_1
X_19040_ _18295_/Y _19048_/A2 _19017_/X _12552_/B _19048_/C1 vssd1 vssd1 vccd1 vccd1
+ _19040_/X sky130_fd_sc_hd__a221o_1
X_16252_ _19668_/Q _17926_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19668_/D sky130_fd_sc_hd__mux2_1
X_13464_ _20011_/Q _20009_/Q _20010_/Q _20008_/Q vssd1 vssd1 vccd1 vccd1 _13464_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_199_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10676_ _11094_/S _10675_/X _10674_/X _12398_/C1 vssd1 vssd1 vccd1 vccd1 _10676_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_173_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15203_ _15396_/A1 _15189_/X _15202_/X vssd1 vssd1 vccd1 vccd1 _16754_/B sky130_fd_sc_hd__a21oi_4
X_12415_ _12409_/X _12414_/X _12415_/S vssd1 vssd1 vccd1 vccd1 _12415_/X sky130_fd_sc_hd__mux2_2
X_16183_ _17432_/A _16183_/B vssd1 vssd1 vccd1 vccd1 _19615_/D sky130_fd_sc_hd__and2_1
X_13395_ _13395_/A _13395_/B vssd1 vssd1 vccd1 vccd1 _13395_/Y sky130_fd_sc_hd__nor2_1
X_12346_ _19429_/Q _20588_/Q _12346_/S vssd1 vssd1 vccd1 vccd1 _12346_/X sky130_fd_sc_hd__mux2_1
X_15134_ _15314_/D _15134_/B vssd1 vssd1 vccd1 vccd1 _15140_/S sky130_fd_sc_hd__or2_4
XFILLER_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19942_ _20181_/CLK _19942_/D vssd1 vssd1 vccd1 vccd1 _19942_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_116_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21018_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15065_ _15057_/X _15064_/X _15577_/S vssd1 vssd1 vccd1 vccd1 _15065_/X sky130_fd_sc_hd__mux2_4
X_12277_ _12277_/A1 _17949_/A1 _12276_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _15988_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_5_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14016_ _12584_/B _14043_/A2 _14034_/B1 _14015_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1
+ _19172_/D sky130_fd_sc_hd__o221a_1
X_11228_ _11228_/A1 _14038_/A2 _11227_/X _11228_/B1 _19855_/Q vssd1 vssd1 vccd1 vccd1
+ _11228_/X sky130_fd_sc_hd__o32a_1
XFILLER_141_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19873_ _20718_/CLK _19873_/D vssd1 vssd1 vccd1 vccd1 _19873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18824_ _19126_/Q _12533_/B _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18824_/Y sky130_fd_sc_hd__a21oi_1
X_11159_ _12230_/A1 _20658_/Q _10842_/S _19367_/Q _12398_/C1 vssd1 vssd1 vccd1 vccd1
+ _11159_/X sky130_fd_sc_hd__o221a_1
XFILLER_268_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18755_ _18755_/A _18755_/B vssd1 vssd1 vccd1 vccd1 _18756_/B sky130_fd_sc_hd__nor2_2
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ _20942_/Q _16044_/A2 _15966_/X vssd1 vssd1 vccd1 vccd1 _15967_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput280 versionID[0] vssd1 vssd1 vccd1 vccd1 input280/X sky130_fd_sc_hd__buf_2
XFILLER_64_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17706_ _20490_/Q _17706_/A1 _17706_/S vssd1 vssd1 vccd1 vccd1 _20490_/D sky130_fd_sc_hd__mux2_1
X_14918_ _14917_/A _10308_/S _14917_/Y vssd1 vssd1 vccd1 vccd1 _15022_/B sky130_fd_sc_hd__a21o_2
XFILLER_247_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18686_ _20945_/Q _18686_/B vssd1 vssd1 vccd1 vccd1 _18686_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ _15898_/A _15925_/B vssd1 vssd1 vccd1 vccd1 _15898_/Y sky130_fd_sc_hd__nand2_1
XFILLER_264_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17637_ _20393_/Q _17914_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20393_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14849_ _11414_/B _11734_/B _15983_/A vssd1 vssd1 vccd1 vccd1 _14849_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17568_ _20328_/Q _17704_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20328_/D sky130_fd_sc_hd__mux2_1
XFILLER_205_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19307_ _20662_/CLK _19307_/D vssd1 vssd1 vccd1 vccd1 _19307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16519_ _19826_/Q _17705_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19826_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17499_ _17505_/A1 _17498_/Y _18104_/A vssd1 vssd1 vccd1 vccd1 _20284_/D sky130_fd_sc_hd__a21oi_1
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19238_ _20291_/CLK _19238_/D vssd1 vssd1 vccd1 vccd1 _19238_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_176_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19169_ _20659_/CLK _19169_/D vssd1 vssd1 vccd1 vccd1 _19169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20013_ _20014_/CLK _20013_/D vssd1 vssd1 vccd1 vccd1 _20013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09824_ _09809_/X _09823_/X _12074_/B1 vssd1 vssd1 vccd1 vccd1 _09824_/X sky130_fd_sc_hd__a21o_2
XFILLER_259_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_14__f_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_99_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09755_ _09753_/X _09754_/X _12006_/S vssd1 vssd1 vccd1 vccd1 _09755_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09686_ _09686_/A _12976_/B _09686_/C _09686_/D vssd1 vssd1 vccd1 vccd1 _09686_/Y
+ sky130_fd_sc_hd__nor4_4
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20915_ _20980_/CLK _20915_/D vssd1 vssd1 vccd1 vccd1 _20915_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20846_ _21040_/CLK _20846_/D vssd1 vssd1 vccd1 vccd1 _20846_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20777_ _21029_/CLK _20777_/D vssd1 vssd1 vccd1 vccd1 _20777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10530_ _10528_/X _10529_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _10530_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _11234_/A _11234_/B _10460_/X vssd1 vssd1 vccd1 vccd1 _10461_/X sky130_fd_sc_hd__or3b_1
XFILLER_136_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ _12200_/A vssd1 vssd1 vccd1 vccd1 _13183_/A sky130_fd_sc_hd__clkinv_4
X_13180_ _16054_/A _13180_/B vssd1 vssd1 vccd1 vccd1 _13181_/B sky130_fd_sc_hd__xnor2_4
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10392_ _20472_/Q _11708_/B _12103_/A1 vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__a21o_1
XFILLER_136_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12131_ _19957_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _12131_/X sky130_fd_sc_hd__or2_1
XFILLER_269_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12062_ _12071_/S _12061_/X _12060_/X _12072_/A1 vssd1 vssd1 vccd1 vccd1 _12062_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout1902 _14482_/A vssd1 vssd1 vccd1 vccd1 _18754_/A sky130_fd_sc_hd__clkbuf_4
Xfanout1913 _18714_/A vssd1 vssd1 vccd1 vccd1 _14758_/C1 sky130_fd_sc_hd__buf_4
X_11013_ _12245_/A1 _11049_/B1 _11012_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _13648_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1924 _16143_/A vssd1 vssd1 vccd1 vccd1 _16165_/C1 sky130_fd_sc_hd__buf_4
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1935 _14185_/C1 vssd1 vssd1 vccd1 vccd1 _18694_/A sky130_fd_sc_hd__clkbuf_4
X_16870_ _20412_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16870_/X sky130_fd_sc_hd__a21o_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1946 fanout1960/X vssd1 vssd1 vccd1 vccd1 _13890_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1957 _18414_/A vssd1 vssd1 vccd1 vccd1 _17974_/B1 sky130_fd_sc_hd__buf_4
Xfanout1968 _17532_/A vssd1 vssd1 vccd1 vccd1 _18905_/A sky130_fd_sc_hd__buf_4
Xfanout970 _17095_/A1 vssd1 vssd1 vccd1 vccd1 _17931_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout981 _17901_/A1 vssd1 vssd1 vccd1 vccd1 _17099_/A1 sky130_fd_sc_hd__buf_4
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _15819_/Y _15820_/X _15817_/X vssd1 vssd1 vccd1 vccd1 _15821_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_65_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1979 _16278_/A vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout992 _16719_/X vssd1 vssd1 vccd1 vccd1 _16964_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18540_ _18932_/A _18540_/B vssd1 vssd1 vccd1 vccd1 _20906_/D sky130_fd_sc_hd__nor2_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _19754_/Q _15999_/A2 _15751_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15752_/X
+ sky130_fd_sc_hd__a211o_1
X_12964_ _19249_/Q _12964_/A2 _16716_/A _19997_/Q vssd1 vssd1 vccd1 vccd1 _14119_/B
+ sky130_fd_sc_hd__a22o_4
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14703_ _17744_/A _16604_/B vssd1 vssd1 vccd1 vccd1 _14704_/C sky130_fd_sc_hd__nor2_1
XFILLER_166_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _18760_/B _18471_/B vssd1 vssd1 vccd1 vccd1 _18473_/A sky130_fd_sc_hd__or2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _20047_/Q _19922_/Q _11915_/S vssd1 vssd1 vccd1 vccd1 _11915_/X sky130_fd_sc_hd__mux2_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15683_ _13419_/A _12565_/B _15682_/X vssd1 vssd1 vccd1 vccd1 _15683_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_330 _20259_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _13199_/B _13233_/B vssd1 vssd1 vccd1 vccd1 _12896_/A sky130_fd_sc_hd__nand2_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_341 _19501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_352 _17706_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17422_ _20265_/Q _20264_/Q vssd1 vssd1 vccd1 vccd1 _17446_/B sky130_fd_sc_hd__nand2_2
XFILLER_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14634_ _17850_/A _17918_/B vssd1 vssd1 vccd1 vccd1 _14635_/C sky130_fd_sc_hd__nor2_1
XANTENNA_363 output482/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_374 _18765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11846_ _12008_/A _19326_/Q _11846_/C vssd1 vssd1 vccd1 vccd1 _11846_/X sky130_fd_sc_hd__or3_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_385 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_396 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17353_ _20225_/Q _17363_/A2 _17352_/X _18692_/A vssd1 vssd1 vccd1 vccd1 _20225_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _16243_/B _14668_/B _17538_/C vssd1 vssd1 vccd1 vccd1 _17918_/B sky130_fd_sc_hd__or3_2
X_11777_ _13523_/A _11779_/B _11776_/Y vssd1 vssd1 vccd1 vccd1 _11778_/C sky130_fd_sc_hd__a21o_1
XFILLER_159_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16304_ _19709_/Q _16306_/C _16303_/Y vssd1 vssd1 vccd1 vccd1 _19709_/D sky130_fd_sc_hd__o21a_1
X_10728_ _10127_/A _10723_/Y _10727_/X _10721_/X vssd1 vssd1 vccd1 vccd1 _10728_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_186_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13516_ _20918_/Q _13598_/A2 _13513_/Y _13515_/X _14110_/A vssd1 vssd1 vccd1 vccd1
+ _13516_/X sky130_fd_sc_hd__a2111o_1
XFILLER_147_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17284_ _17284_/A _17290_/B _17290_/C vssd1 vssd1 vccd1 vccd1 _17284_/X sky130_fd_sc_hd__and3_1
X_14496_ _19274_/Q _17859_/A1 _14519_/S vssd1 vssd1 vccd1 vccd1 _19274_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19023_ _21030_/Q _19015_/B _19022_/X _18728_/A vssd1 vssd1 vccd1 vccd1 _21030_/D
+ sky130_fd_sc_hd__o211a_1
X_16235_ _13441_/X _16235_/B vssd1 vssd1 vccd1 vccd1 _16235_/X sky130_fd_sc_hd__and2b_1
X_10659_ _20468_/Q _20308_/Q _12381_/S vssd1 vssd1 vccd1 vccd1 _10659_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13447_ _13600_/A _13600_/B _12771_/C vssd1 vssd1 vccd1 vccd1 _13448_/B sky130_fd_sc_hd__o21a_1
XFILLER_256_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16166_ _16878_/B _16190_/S vssd1 vssd1 vccd1 vccd1 _16166_/Y sky130_fd_sc_hd__nand2_1
X_13378_ _19229_/Q _13378_/B vssd1 vssd1 vccd1 vccd1 _13378_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15117_ _15407_/S _15112_/X _15116_/X vssd1 vssd1 vccd1 vccd1 _15117_/X sky130_fd_sc_hd__a21o_1
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12329_ _11726_/S _11367_/B _12708_/A vssd1 vssd1 vccd1 vccd1 _12329_/Y sky130_fd_sc_hd__a21oi_1
X_16097_ _19573_/Q _16077_/B _16097_/B1 vssd1 vssd1 vccd1 vccd1 _16097_/X sky130_fd_sc_hd__o21a_1
XFILLER_173_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19925_ _20681_/CLK _19925_/D vssd1 vssd1 vccd1 vccd1 _19925_/Q sky130_fd_sc_hd__dfxtp_1
X_15048_ _15046_/X _15170_/B _15170_/A vssd1 vssd1 vccd1 vccd1 _15048_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19856_ _20014_/CLK _19856_/D vssd1 vssd1 vccd1 vccd1 _19856_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_229_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18807_ _18483_/X _18819_/B _18805_/X _18806_/Y vssd1 vssd1 vccd1 vccd1 _18808_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19787_ _20710_/CLK _19787_/D vssd1 vssd1 vccd1 vccd1 _19787_/Q sky130_fd_sc_hd__dfxtp_1
X_16999_ input66/X input101/X _17009_/S vssd1 vssd1 vccd1 vccd1 _16999_/X sky130_fd_sc_hd__mux2_8
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_84_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _20410_/CLK sky130_fd_sc_hd__clkbuf_16
X_09540_ _12480_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _09540_/X sky130_fd_sc_hd__and2_1
XFILLER_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18738_ _18748_/A _18738_/B vssd1 vssd1 vccd1 vccd1 _20969_/D sky130_fd_sc_hd__and2_1
XFILLER_224_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20711_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_236_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18669_ _18966_/A _18669_/B vssd1 vssd1 vccd1 vccd1 _20940_/D sky130_fd_sc_hd__nor2_1
XFILLER_92_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20700_ _20711_/CLK _20700_/D vssd1 vssd1 vccd1 vccd1 _20700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20631_ _20663_/CLK _20631_/D vssd1 vssd1 vccd1 vccd1 _20631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20562_ _20694_/CLK _20562_/D vssd1 vssd1 vccd1 vccd1 _20562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20493_ _20657_/CLK _20493_/D vssd1 vssd1 vccd1 vccd1 _20493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1209 _15095_/X vssd1 vssd1 vccd1 vccd1 _15457_/B1 sky130_fd_sc_hd__buf_2
XFILLER_247_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09807_ _10057_/S _09793_/X _09794_/X vssd1 vssd1 vccd1 vccd1 _09807_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09738_ _09738_/A _11213_/B vssd1 vssd1 vccd1 vccd1 _09738_/Y sky130_fd_sc_hd__nand2_8
XFILLER_228_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09669_ _18163_/B _11235_/A vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__or2_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11718_/S _11697_/X _11699_/X vssd1 vssd1 vccd1 vccd1 _11700_/X sky130_fd_sc_hd__a21o_1
XFILLER_243_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12680_ _19498_/Q _12680_/B vssd1 vssd1 vccd1 vccd1 _12680_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _20576_/Q _11708_/B vssd1 vssd1 vccd1 vccd1 _11631_/X sky130_fd_sc_hd__or2_1
X_20829_ _21023_/CLK _20829_/D vssd1 vssd1 vccd1 vccd1 _20829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14350_ _20289_/Q _14431_/A2 _14431_/B1 input230/X vssd1 vssd1 vccd1 vccd1 _14352_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _09986_/A _19814_/Q _19318_/Q _09928_/S vssd1 vssd1 vccd1 vccd1 _11562_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10513_ _20128_/Q _20096_/Q _11295_/S vssd1 vssd1 vccd1 vccd1 _10513_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13301_ _13300_/B _13300_/C _13300_/A vssd1 vssd1 vccd1 vccd1 _13301_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_156_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14281_ _19510_/Q _14281_/B vssd1 vssd1 vccd1 vccd1 _14282_/B sky130_fd_sc_hd__nand2_1
X_11493_ _19511_/Q _15659_/A _11726_/S vssd1 vssd1 vccd1 vccd1 _11734_/B sky130_fd_sc_hd__mux2_4
X_16020_ _19732_/Q _16039_/B _16012_/X _16019_/X vssd1 vssd1 vccd1 vccd1 _16020_/X
+ sky130_fd_sc_hd__o22a_1
X_13232_ _20939_/Q _13366_/C1 _13323_/C _13231_/X _18687_/B vssd1 vssd1 vccd1 vccd1
+ _13232_/X sky130_fd_sc_hd__a221o_1
X_10444_ _11266_/A1 _19313_/Q _11270_/A2 _11256_/S vssd1 vssd1 vccd1 vccd1 _10444_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ _11497_/A _13162_/A _13162_/B _11496_/Y vssd1 vssd1 vccd1 vccd1 _13419_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_123_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10375_ _11242_/A1 _14011_/A2 _10374_/X _11242_/B1 _19850_/Q vssd1 vssd1 vccd1 vccd1
+ _10375_/X sky130_fd_sc_hd__o32a_1
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ _12110_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__nand2b_1
XFILLER_269_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17971_ _20728_/Q _20727_/Q _17971_/C vssd1 vssd1 vccd1 vccd1 _17976_/C sky130_fd_sc_hd__and3_1
X_13094_ _20911_/Q _13092_/X _13272_/B vssd1 vssd1 vccd1 vccd1 _13094_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19710_ _20757_/CLK _19710_/D vssd1 vssd1 vccd1 vccd1 _19710_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1710 _12270_/B1 vssd1 vssd1 vccd1 vccd1 _11378_/S sky130_fd_sc_hd__buf_6
X_16922_ _19236_/Q _16980_/A2 _16980_/B1 _19105_/Q _16921_/X vssd1 vssd1 vccd1 vccd1
+ _16922_/X sky130_fd_sc_hd__o221a_1
X_12045_ _19424_/Q _12053_/S _12044_/X _12051_/C1 vssd1 vssd1 vccd1 vccd1 _12045_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout1721 _12752_/A vssd1 vssd1 vccd1 vccd1 _12138_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout1732 _12312_/A1 vssd1 vssd1 vccd1 vccd1 _12371_/A1 sky130_fd_sc_hd__buf_6
XFILLER_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1743 _09503_/Y vssd1 vssd1 vccd1 vccd1 _12519_/C sky130_fd_sc_hd__buf_12
XFILLER_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1754 _14042_/S vssd1 vssd1 vccd1 vccd1 _14036_/S sky130_fd_sc_hd__buf_6
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19641_ _20679_/CLK _19641_/D vssd1 vssd1 vccd1 vccd1 _19641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16853_ _19228_/Q _16996_/A2 _16996_/B1 _19097_/Q _16852_/X vssd1 vssd1 vccd1 vccd1
+ _16853_/X sky130_fd_sc_hd__o221a_1
Xfanout1765 _09488_/Y vssd1 vssd1 vccd1 vccd1 _14524_/A1 sky130_fd_sc_hd__buf_6
XFILLER_266_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1776 _20721_/Q vssd1 vssd1 vccd1 vccd1 output482/A sky130_fd_sc_hd__buf_12
Xfanout1787 _18209_/A1 vssd1 vssd1 vccd1 vccd1 _18223_/B sky130_fd_sc_hd__buf_12
XFILLER_281_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15804_ _16017_/C1 _15803_/X _15799_/X vssd1 vssd1 vccd1 vccd1 _15804_/X sky130_fd_sc_hd__o21a_2
XFILLER_19_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1798 _20182_/Q vssd1 vssd1 vccd1 vccd1 _12548_/B sky130_fd_sc_hd__clkbuf_4
X_19572_ _20341_/CLK _19572_/D vssd1 vssd1 vccd1 vccd1 _19572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16784_ _16869_/A _16784_/B vssd1 vssd1 vccd1 vccd1 _16784_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13996_ _14035_/A1 _14011_/A2 _11241_/X _14035_/B1 _19847_/Q vssd1 vssd1 vccd1 vccd1
+ _14077_/C sky130_fd_sc_hd__o32a_1
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18523_ _18671_/B _18523_/B vssd1 vssd1 vccd1 vccd1 _18523_/X sky130_fd_sc_hd__or2_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15735_ _13417_/A _15981_/B _15219_/Y vssd1 vssd1 vccd1 vccd1 _15735_/Y sky130_fd_sc_hd__o21ai_1
X_12947_ _19263_/Q _12950_/B2 _16716_/A _20011_/Q vssd1 vssd1 vccd1 vccd1 _16714_/B
+ sky130_fd_sc_hd__a22o_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18454_ _18746_/A _18454_/B vssd1 vssd1 vccd1 vccd1 _20881_/D sky130_fd_sc_hd__and2_1
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15666_ _20931_/Q _15995_/A2 _15665_/X vssd1 vssd1 vccd1 vccd1 _15666_/X sky130_fd_sc_hd__o21a_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12878_ _13233_/A _12878_/B vssd1 vssd1 vccd1 vccd1 _13199_/B sky130_fd_sc_hd__nor2_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 _13780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_171 _19108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_182 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17405_ _17402_/Y _17404_/X _17403_/X _17434_/A vssd1 vssd1 vccd1 vccd1 _20250_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14617_ _19381_/Q _17099_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19381_/D sky130_fd_sc_hd__mux2_1
XANTENNA_193 _19541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ _09901_/S _11828_/X _11827_/X _12140_/C1 vssd1 vssd1 vccd1 vccd1 _11829_/X
+ sky130_fd_sc_hd__a211o_1
X_18385_ _18556_/B _18385_/B vssd1 vssd1 vccd1 vccd1 _18385_/Y sky130_fd_sc_hd__nand2_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15597_ _21027_/Q _20995_/Q _15993_/S vssd1 vssd1 vccd1 vccd1 _15597_/X sky130_fd_sc_hd__mux2_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17336_ _17337_/A _17336_/B vssd1 vssd1 vccd1 vccd1 _17336_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14548_ _19318_/Q _17202_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19318_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17267_ _20194_/Q _17330_/A2 _17279_/C1 vssd1 vssd1 vccd1 vccd1 _17267_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_131_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21015_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14479_ _20235_/Q _19264_/Q _14483_/S vssd1 vssd1 vccd1 vccd1 _14480_/B sky130_fd_sc_hd__mux2_1
X_19006_ _18210_/Y _18982_/B _19016_/B1 _19005_/X vssd1 vssd1 vccd1 vccd1 _21022_/D
+ sky130_fd_sc_hd__o211a_1
X_16218_ _19641_/Q _17870_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19641_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17198_ _20162_/Q _17932_/A1 _17215_/S vssd1 vssd1 vccd1 vccd1 _20162_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16149_ _19598_/Q _16196_/S _16148_/Y _16197_/A vssd1 vssd1 vccd1 vccd1 _19598_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_216_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19908_ _20539_/CLK _19908_/D vssd1 vssd1 vccd1 vccd1 _19908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19839_ _20621_/CLK _19839_/D vssd1 vssd1 vccd1 vccd1 _19839_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09523_ input44/X vssd1 vssd1 vccd1 vccd1 _09523_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20614_ _20717_/CLK _20614_/D vssd1 vssd1 vccd1 vccd1 _20614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20545_ _20585_/CLK _20545_/D vssd1 vssd1 vccd1 vccd1 _20545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20476_ _20702_/CLK _20476_/D vssd1 vssd1 vccd1 vccd1 _20476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10160_ _11363_/A1 _10156_/X _10159_/X _09689_/C vssd1 vssd1 vccd1 vccd1 _10160_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput370 _13477_/X vssd1 vssd1 vccd1 vccd1 core_wb_stb_o sky130_fd_sc_hd__buf_4
XFILLER_121_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1006 _14904_/X vssd1 vssd1 vccd1 vccd1 _16049_/A1 sky130_fd_sc_hd__clkbuf_16
Xoutput381 _13805_/X vssd1 vssd1 vccd1 vccd1 din0[14] sky130_fd_sc_hd__buf_4
XFILLER_248_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput392 _13815_/X vssd1 vssd1 vccd1 vccd1 din0[24] sky130_fd_sc_hd__buf_4
X_10091_ _19674_/Q _20162_/Q _10092_/S vssd1 vssd1 vccd1 vccd1 _10091_/X sky130_fd_sc_hd__mux2_1
Xfanout1017 _18864_/A2 vssd1 vssd1 vccd1 vccd1 _18974_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_273_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1028 _16711_/Y vssd1 vssd1 vccd1 vccd1 _16963_/A2 sky130_fd_sc_hd__buf_6
Xfanout1039 _17051_/A1 vssd1 vssd1 vccd1 vccd1 _17678_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21028_ _21030_/CLK _21028_/D vssd1 vssd1 vccd1 vccd1 _21028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ _17421_/A _17451_/B vssd1 vssd1 vccd1 vccd1 _17231_/A sky130_fd_sc_hd__nor2_2
XFILLER_75_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _12483_/Y _12800_/X _15768_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12801_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_216_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10993_ _11336_/A _20089_/Q _10983_/S _10991_/X _10992_/X vssd1 vssd1 vccd1 vccd1
+ _10993_/X sky130_fd_sc_hd__a311o_1
XFILLER_16_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13781_ _13612_/A split3/X _15127_/A _13493_/Y _13244_/X vssd1 vssd1 vccd1 vccd1
+ _13781_/X sky130_fd_sc_hd__a32o_4
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15520_ _15495_/X _15503_/Y _15519_/X _15520_/B2 vssd1 vssd1 vccd1 vccd1 _15520_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12730_/X _12731_/Y _12716_/B vssd1 vssd1 vccd1 vccd1 _12736_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _17302_/A _15482_/A2 _15016_/A _20796_/Q _15450_/X vssd1 vssd1 vccd1 vccd1
+ _15451_/X sky130_fd_sc_hd__a221o_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _19159_/Q _12479_/X _12578_/B _09621_/A vssd1 vssd1 vccd1 vccd1 _12674_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14402_ _14400_/Y _14402_/B vssd1 vssd1 vccd1 vccd1 _14405_/A sky130_fd_sc_hd__nand2b_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18170_ _18466_/B vssd1 vssd1 vccd1 vccd1 _18170_/Y sky130_fd_sc_hd__inv_2
X_11614_ _11922_/A1 _13717_/A _12158_/B1 vssd1 vssd1 vccd1 vccd1 _11614_/Y sky130_fd_sc_hd__o21ai_1
X_15382_ _20730_/Q _15445_/A2 _15445_/B1 _20762_/Q vssd1 vssd1 vccd1 vccd1 _15382_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12708_/A _13002_/A vssd1 vssd1 vccd1 vccd1 _12628_/A sky130_fd_sc_hd__and2_1
XFILLER_204_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ _20089_/Q _17189_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20089_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14333_ _14333_/A _14333_/B _14333_/C vssd1 vssd1 vccd1 vccd1 _14335_/B sky130_fd_sc_hd__and3_1
X_11545_ _11563_/S _11542_/X _11544_/X vssd1 vssd1 vccd1 vccd1 _11545_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _20024_/Q _17679_/A1 _17080_/S vssd1 vssd1 vccd1 vccd1 _20024_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11476_ _20414_/Q _20350_/Q _12165_/S vssd1 vssd1 vccd1 vccd1 _11477_/B sky130_fd_sc_hd__mux2_1
X_14264_ _14275_/A1 _14263_/X _13386_/Y vssd1 vssd1 vccd1 vccd1 _14265_/C sky130_fd_sc_hd__o21a_1
XFILLER_100_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ _15246_/A _16001_/Y _16002_/Y _15981_/A _12578_/A vssd1 vssd1 vccd1 vccd1
+ _16003_/X sky130_fd_sc_hd__o32a_1
XFILLER_100_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13215_ _13011_/Y _13012_/X _13086_/A _13227_/A vssd1 vssd1 vccd1 vccd1 _13215_/X
+ sky130_fd_sc_hd__a211o_1
X_10427_ _10425_/X _10426_/X _10585_/S vssd1 vssd1 vccd1 vccd1 _10427_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _19222_/Q _14205_/A2 _14194_/X _18710_/A vssd1 vssd1 vccd1 vccd1 _19222_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13146_ _11055_/B _13145_/A _13145_/B _11053_/Y vssd1 vssd1 vccd1 vccd1 _13523_/B
+ sky130_fd_sc_hd__a31o_4
X_10358_ _19637_/Q _19943_/Q _19281_/Q _20068_/Q _11292_/S0 _11290_/C vssd1 vssd1
+ vccd1 vccd1 _10358_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17954_ _21044_/Q _20722_/Q vssd1 vssd1 vccd1 vccd1 _17959_/C sky130_fd_sc_hd__and2b_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _20963_/Q _20897_/Q _13076_/X vssd1 vssd1 vccd1 vccd1 _13327_/A sky130_fd_sc_hd__o21ai_4
X_10289_ _19589_/Q _10288_/X _11240_/S vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__mux2_2
XFILLER_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1540 _10137_/C vssd1 vssd1 vccd1 vccd1 _11257_/S sky130_fd_sc_hd__buf_6
XFILLER_39_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16905_ _20416_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16905_/X sky130_fd_sc_hd__a21o_1
X_12028_ _12850_/A1 _12027_/X _09729_/Y vssd1 vssd1 vccd1 vccd1 _12028_/Y sky130_fd_sc_hd__a21oi_1
Xfanout1551 _12219_/S vssd1 vssd1 vccd1 vccd1 _12381_/S sky130_fd_sc_hd__buf_6
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17885_ _17919_/A _17885_/B _17885_/C vssd1 vssd1 vccd1 vccd1 _17885_/X sky130_fd_sc_hd__and3_4
Xfanout1562 _11161_/S vssd1 vssd1 vccd1 vccd1 _12316_/S sky130_fd_sc_hd__buf_6
XFILLER_78_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1573 _09624_/Y vssd1 vssd1 vccd1 vccd1 _09689_/C sky130_fd_sc_hd__buf_8
XFILLER_254_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1584 _11597_/C1 vssd1 vssd1 vccd1 vccd1 _11009_/B2 sky130_fd_sc_hd__clkbuf_8
XFILLER_93_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19624_ _20670_/CLK _19624_/D vssd1 vssd1 vccd1 vccd1 _19624_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1595 _11600_/C1 vssd1 vssd1 vccd1 vccd1 _11008_/A3 sky130_fd_sc_hd__buf_6
X_16836_ _16805_/X _16833_/Y _16835_/X _16932_/A1 vssd1 vssd1 vccd1 vccd1 _16836_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19555_ _20263_/CLK _19555_/D vssd1 vssd1 vccd1 vccd1 _19555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16767_ _17006_/A1 _15243_/X _16766_/X vssd1 vssd1 vccd1 vccd1 _16767_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13979_ _19192_/Q _14065_/C _14003_/S vssd1 vssd1 vccd1 vccd1 _13979_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18506_ _20895_/Q _18474_/S _18505_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18507_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15718_ _21031_/Q _20999_/Q _15993_/S vssd1 vssd1 vccd1 vccd1 _15718_/X sky130_fd_sc_hd__mux2_1
X_19486_ _20713_/CLK _19486_/D vssd1 vssd1 vccd1 vccd1 _19486_/Q sky130_fd_sc_hd__dfxtp_1
X_16698_ _19953_/Q _17876_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19953_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18437_ _20873_/Q _18275_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18438_/B sky130_fd_sc_hd__mux2_1
XFILLER_278_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15649_ _15649_/A1 _16063_/A2 _13427_/C _15922_/B2 vssd1 vssd1 vccd1 vccd1 _15650_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18368_ _20839_/Q _18385_/B _18367_/Y _18740_/A vssd1 vssd1 vccd1 vccd1 _20839_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_193_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17319_ _20212_/Q _17232_/X _17318_/X _17974_/B1 vssd1 vssd1 vccd1 vccd1 _20212_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18299_ _18299_/A1 _14406_/B _18298_/Y vssd1 vssd1 vccd1 vccd1 _18550_/B sky130_fd_sc_hd__o21ai_4
XFILLER_119_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20330_ _20491_/CLK _20330_/D vssd1 vssd1 vccd1 vccd1 _20330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20261_ _20261_/CLK _20261_/D vssd1 vssd1 vccd1 vccd1 _20261_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_134_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20192_ _20428_/CLK _20192_/D vssd1 vssd1 vccd1 vccd1 _20192_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput109 dout1[11] vssd1 vssd1 vccd1 vccd1 input109/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09506_ _11384_/S vssd1 vssd1 vccd1 vccd1 _10525_/S sky130_fd_sc_hd__inv_2
XFILLER_53_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_60 _17336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_71 _09504_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11326_/X _11329_/X _10127_/A vssd1 vssd1 vccd1 vccd1 _11330_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_166_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_82 _09946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20528_ _20667_/CLK _20528_/D vssd1 vssd1 vccd1 vccd1 _20528_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_93 _12040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11261_ _11268_/A _20589_/Q _11261_/C vssd1 vssd1 vccd1 vccd1 _11261_/X sky130_fd_sc_hd__and3_1
X_20459_ _20468_/CLK _20459_/D vssd1 vssd1 vccd1 vccd1 _20459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10212_ _11336_/A _19445_/Q _10217_/S vssd1 vssd1 vccd1 vccd1 _10212_/X sky130_fd_sc_hd__and3_1
X_13000_ _19245_/Q _13104_/B vssd1 vssd1 vccd1 vccd1 _13001_/B sky130_fd_sc_hd__nand2_1
XFILLER_97_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11192_ _19799_/Q _11192_/A2 _11190_/X _15129_/A0 _11191_/X vssd1 vssd1 vccd1 vccd1
+ _11192_/X sky130_fd_sc_hd__o221a_1
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10143_ _12513_/C _10135_/X _10139_/X _09621_/A vssd1 vssd1 vccd1 vccd1 _10143_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ _14951_/A _14951_/B _14951_/C _14973_/C vssd1 vssd1 vccd1 vccd1 _14966_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10074_ _12072_/C1 _10062_/X _10065_/X _10073_/X vssd1 vssd1 vccd1 vccd1 _10074_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13902_ _13902_/A _13902_/B vssd1 vssd1 vccd1 vccd1 _13902_/Y sky130_fd_sc_hd__nand2_4
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17670_ _20456_/Q _17947_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20456_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14882_ _14882_/A _14882_/B _15494_/B vssd1 vssd1 vccd1 vccd1 _14885_/B sky130_fd_sc_hd__and3_4
XFILLER_235_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16621_ _19880_/Q _17935_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19880_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ _20003_/Q split1/X _13787_/X _16279_/B vssd1 vssd1 vccd1 vccd1 _13833_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_251_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19340_ _20718_/CLK _19340_/D vssd1 vssd1 vccd1 vccd1 _19340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16552_ _19842_/Q _16576_/A2 _16576_/B1 input12/X vssd1 vssd1 vccd1 vccd1 _16553_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_204_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13764_ _13764_/A _13764_/B vssd1 vssd1 vccd1 vccd1 _13765_/B sky130_fd_sc_hd__nor2_8
X_10976_ _11061_/A _16075_/A vssd1 vssd1 vccd1 vccd1 _10976_/Y sky130_fd_sc_hd__nor2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15503_ _15258_/A _15498_/Y _15502_/X vssd1 vssd1 vccd1 vccd1 _15503_/Y sky130_fd_sc_hd__o21ai_1
X_19271_ _20690_/CLK _19271_/D vssd1 vssd1 vccd1 vccd1 _19271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12715_ _12726_/A _12726_/B vssd1 vssd1 vccd1 vccd1 _12715_/Y sky130_fd_sc_hd__nor2_1
X_16483_ _19792_/Q _17806_/A1 _16483_/S vssd1 vssd1 vccd1 vccd1 _19792_/D sky130_fd_sc_hd__mux2_1
XFILLER_241_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13695_ _13740_/A _13693_/X _13694_/X _13740_/B vssd1 vssd1 vccd1 vccd1 _13697_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18222_ _18416_/A _18222_/B vssd1 vssd1 vccd1 vccd1 _20798_/D sky130_fd_sc_hd__and2_1
XFILLER_204_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15434_ _15442_/B _15127_/B _15220_/A vssd1 vssd1 vccd1 vccd1 _15434_/X sky130_fd_sc_hd__a21o_1
XFILLER_231_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ _19498_/Q _12680_/B _19499_/Q vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__a21oi_1
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18153_ _18136_/Y _18152_/X _18138_/A vssd1 vssd1 vccd1 vccd1 _18154_/B sky130_fd_sc_hd__o21a_1
XFILLER_7_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15365_ _15365_/A _15365_/B _15365_/C vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__and3_1
XFILLER_178_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12577_ _12577_/A _12577_/B vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__or2_2
XFILLER_8_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17104_ _20074_/Q _17872_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20074_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _14325_/A _14312_/B _14315_/X vssd1 vssd1 vccd1 vccd1 _14316_/X sky130_fd_sc_hd__a21bo_1
XFILLER_117_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18084_ _20768_/Q _18085_/C _20769_/Q vssd1 vssd1 vccd1 vccd1 _18086_/B sky130_fd_sc_hd__a21oi_1
X_11528_ _11526_/X _11527_/X _11528_/S vssd1 vssd1 vccd1 vccd1 _11528_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15296_ _15066_/S _15295_/X _15548_/B1 vssd1 vssd1 vccd1 vccd1 _15297_/A sky130_fd_sc_hd__o21ai_1
X_17035_ _20013_/Q input199/X _17038_/S vssd1 vssd1 vccd1 vccd1 _20013_/D sky130_fd_sc_hd__mux2_1
X_14247_ _20279_/Q _14267_/A2 _14267_/B1 input219/X vssd1 vssd1 vccd1 vccd1 _14249_/B
+ sky130_fd_sc_hd__a22o_4
X_11459_ _19415_/Q _20574_/Q _12185_/S vssd1 vssd1 vccd1 vccd1 _11459_/X sky130_fd_sc_hd__mux2_1
XFILLER_264_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14178_ _14176_/Y _14178_/B vssd1 vssd1 vccd1 vccd1 _14181_/A sky130_fd_sc_hd__nand2b_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13106_/B _12909_/X _12629_/Y vssd1 vssd1 vccd1 vccd1 _13129_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18986_ _18160_/Y _18982_/B _18984_/X _19016_/B1 vssd1 vssd1 vccd1 vccd1 _21012_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _20706_/Q _17937_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20706_/D sky130_fd_sc_hd__mux2_1
XFILLER_285_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1370 _14267_/A2 vssd1 vssd1 vccd1 vccd1 _14117_/A sky130_fd_sc_hd__buf_6
XFILLER_39_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1381 _09931_/S vssd1 vssd1 vccd1 vccd1 _09928_/S sky130_fd_sc_hd__buf_4
X_17868_ _20641_/Q _17902_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20641_/D sky130_fd_sc_hd__mux2_1
Xfanout1392 _11848_/S0 vssd1 vssd1 vccd1 vccd1 _12185_/S sky130_fd_sc_hd__buf_6
XFILLER_253_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19607_ _19607_/CLK _19607_/D vssd1 vssd1 vccd1 vccd1 _19607_/Q sky130_fd_sc_hd__dfxtp_1
X_16819_ _16846_/A input78/X vssd1 vssd1 vccd1 vccd1 _16819_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17799_ _20576_/Q _17939_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20576_/D sky130_fd_sc_hd__mux2_1
XFILLER_241_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19538_ _19603_/CLK _19538_/D vssd1 vssd1 vccd1 vccd1 _19538_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_241_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19469_ _20468_/CLK _19469_/D vssd1 vssd1 vccd1 vccd1 _19469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20313_ _20701_/CLK _20313_/D vssd1 vssd1 vccd1 vccd1 _20313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput80 dout0[43] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput91 dout0[53] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20244_ _20296_/CLK _20244_/D vssd1 vssd1 vccd1 vccd1 _20244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20175_ _20482_/CLK _20175_/D vssd1 vssd1 vccd1 vccd1 _20175_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ _09986_/A _19322_/Q _09986_/C vssd1 vssd1 vccd1 vccd1 _09986_/X sky130_fd_sc_hd__or3_1
XFILLER_249_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10830_ _09618_/A _10816_/X _10817_/X vssd1 vssd1 vccd1 vccd1 _10830_/X sky130_fd_sc_hd__o21a_1
XFILLER_198_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10761_ _12400_/A1 _10753_/X _10760_/X _10746_/X vssd1 vssd1 vccd1 vccd1 _10761_/X
+ sky130_fd_sc_hd__o31a_4
XFILLER_158_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12500_ _19156_/Q _19155_/Q _19154_/Q _12500_/D vssd1 vssd1 vccd1 vccd1 _15095_/B
+ sky130_fd_sc_hd__and4_4
XFILLER_12_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10692_ _10692_/A _20664_/Q _12406_/C vssd1 vssd1 vccd1 vccd1 _10692_/X sky130_fd_sc_hd__or3_1
XFILLER_197_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13480_ _19661_/D _17041_/B vssd1 vssd1 vccd1 vccd1 _13480_/Y sky130_fd_sc_hd__nor2_2
XFILLER_240_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12431_ _12431_/A1 _12430_/X _12275_/A vssd1 vssd1 vccd1 vccd1 _12431_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15150_ _12486_/Y _12666_/A _15127_/A _15442_/A _15150_/C1 vssd1 vssd1 vccd1 vccd1
+ _15150_/X sky130_fd_sc_hd__a221o_2
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ _19525_/Q _12361_/Y _15949_/A vssd1 vssd1 vccd1 vccd1 _14882_/A sky130_fd_sc_hd__mux2_8
XFILLER_32_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14101_ _14105_/A _14107_/B _14101_/C vssd1 vssd1 vccd1 vccd1 _14101_/X sky130_fd_sc_hd__or3_1
XFILLER_153_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ _19494_/Q _11313_/B vssd1 vssd1 vccd1 vccd1 _11313_/Y sky130_fd_sc_hd__nand2_1
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15081_ _15081_/A _15133_/B vssd1 vssd1 vccd1 vccd1 _15081_/X sky130_fd_sc_hd__and2_1
X_12293_ _10127_/A _12292_/X _12291_/X vssd1 vssd1 vccd1 vccd1 _12293_/X sky130_fd_sc_hd__a21o_2
XFILLER_126_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14032_ _14041_/A1 _14041_/A2 _10038_/X _14041_/B1 _19859_/Q vssd1 vssd1 vccd1 vccd1
+ _14101_/C sky130_fd_sc_hd__o32a_1
X_11244_ _10553_/A _10553_/B _11243_/X _18163_/B vssd1 vssd1 vccd1 vccd1 _11244_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_162_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11175_ _18765_/A _19463_/Q _19431_/Q _11174_/S _09695_/A vssd1 vssd1 vccd1 vccd1
+ _11175_/X sky130_fd_sc_hd__a221o_1
X_18840_ _20991_/Q _18840_/B vssd1 vssd1 vccd1 vccd1 _18840_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10126_ _10035_/Y _10120_/X _10125_/X _10118_/X _10024_/X vssd1 vssd1 vccd1 vccd1
+ _10127_/B sky130_fd_sc_hd__a32o_1
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18771_ _18570_/B _18768_/X _18770_/X vssd1 vssd1 vccd1 vccd1 _18772_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15983_ _15983_/A _15983_/B vssd1 vssd1 vccd1 vccd1 _15983_/Y sky130_fd_sc_hd__nand2_1
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17722_ _20503_/Q _17896_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20503_/D sky130_fd_sc_hd__mux2_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14934_ _14980_/B _14973_/B vssd1 vssd1 vccd1 vccd1 _14948_/A sky130_fd_sc_hd__nand2b_4
X_10057_ _10055_/X _10056_/X _10057_/S vssd1 vssd1 vccd1 vccd1 _10057_/X sky130_fd_sc_hd__mux2_1
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _20439_/Q _17687_/A1 _17657_/S vssd1 vssd1 vccd1 vccd1 _20439_/D sky130_fd_sc_hd__mux2_1
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ _14859_/X _14864_/Y _15170_/A vssd1 vssd1 vccd1 vccd1 _14865_/X sky130_fd_sc_hd__mux2_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ _17850_/A _16604_/B vssd1 vssd1 vccd1 vccd1 _16605_/C sky130_fd_sc_hd__nor2_1
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13816_ _13816_/A1 _13750_/B _13816_/B1 input232/X vssd1 vssd1 vccd1 vccd1 _13816_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17584_ _20342_/Q _17895_/A1 _17601_/S vssd1 vssd1 vccd1 vccd1 _20342_/D sky130_fd_sc_hd__mux2_1
X_14796_ _19145_/Q _14802_/A2 _14795_/X _17536_/D vssd1 vssd1 vccd1 vccd1 _19522_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19323_ _20645_/CLK _19323_/D vssd1 vssd1 vccd1 vccd1 _19323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16535_ _16557_/A _16535_/B vssd1 vssd1 vccd1 vccd1 _19833_/D sky130_fd_sc_hd__or2_1
XFILLER_17_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13747_ _13777_/A _13747_/B vssd1 vssd1 vccd1 vccd1 _13747_/X sky130_fd_sc_hd__or2_1
X_10959_ _20154_/Q _11379_/B _11212_/S vssd1 vssd1 vccd1 vccd1 _10959_/X sky130_fd_sc_hd__o21a_1
XFILLER_204_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19254_ _20818_/CLK _19254_/D vssd1 vssd1 vccd1 vccd1 _19254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16466_ _19775_/Q _17929_/A1 _16483_/S vssd1 vssd1 vccd1 vccd1 _19775_/D sky130_fd_sc_hd__mux2_1
XFILLER_231_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13678_ _13679_/B vssd1 vssd1 vccd1 vccd1 _13678_/Y sky130_fd_sc_hd__inv_2
X_18205_ _18493_/B vssd1 vssd1 vccd1 vccd1 _18205_/Y sky130_fd_sc_hd__clkinv_4
X_15417_ _20891_/Q _14971_/A _15566_/B1 _15416_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15417_/X sky130_fd_sc_hd__a221o_1
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19185_ _19574_/CLK _19185_/D vssd1 vssd1 vccd1 vccd1 _19185_/Q sky130_fd_sc_hd__dfxtp_1
X_12629_ _13106_/A _12629_/B vssd1 vssd1 vccd1 vccd1 _12629_/Y sky130_fd_sc_hd__nand2_1
X_16397_ _18080_/A _16402_/C vssd1 vssd1 vccd1 vccd1 _16397_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18136_ _18136_/A _18136_/B vssd1 vssd1 vccd1 vccd1 _18136_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20701_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15348_ _15246_/A _15346_/X _15347_/Y _12630_/Y _15348_/B2 vssd1 vssd1 vccd1 vccd1
+ _15348_/X sky130_fd_sc_hd__o32a_1
XFILLER_156_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18067_ _20762_/Q _18069_/C _18066_/Y vssd1 vssd1 vccd1 vccd1 _20762_/D sky130_fd_sc_hd__o21a_1
X_15279_ _19739_/Q _15453_/A2 _15269_/X _15396_/A1 _15278_/X vssd1 vssd1 vccd1 vccd1
+ _15279_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17018_ _19996_/Q input201/X _17849_/S vssd1 vssd1 vccd1 vccd1 _19996_/D sky130_fd_sc_hd__mux2_1
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout607 _14594_/S vssd1 vssd1 vccd1 vccd1 _14596_/S sky130_fd_sc_hd__buf_12
X_09840_ _20140_/Q _20108_/Q _10397_/S vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__mux2_1
Xfanout618 _14488_/X vssd1 vssd1 vccd1 vccd1 _14519_/S sky130_fd_sc_hd__buf_6
XFILLER_217_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout629 _13900_/A2 vssd1 vssd1 vccd1 vccd1 _13896_/B1 sky130_fd_sc_hd__buf_4
XFILLER_59_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_13__f_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ _20141_/Q _20109_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _09771_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18969_ _19147_/Q _18976_/A2 _18767_/B vssd1 vssd1 vccd1 vccd1 _18969_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_246_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20931_ _20998_/CLK _20931_/D vssd1 vssd1 vccd1 vccd1 _20931_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20862_ _20862_/CLK _20862_/D vssd1 vssd1 vccd1 vccd1 _20862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20793_ _20863_/CLK _20793_/D vssd1 vssd1 vccd1 vccd1 _20793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20227_ _21018_/CLK _20227_/D vssd1 vssd1 vccd1 vccd1 _20227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20158_ _20559_/CLK _20158_/D vssd1 vssd1 vccd1 vccd1 _20158_/Q sky130_fd_sc_hd__dfxtp_1
X_09969_ _09901_/S _09968_/X _09967_/X _12151_/A1 vssd1 vssd1 vccd1 vccd1 _09969_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20089_ _20565_/CLK _20089_/D vssd1 vssd1 vccd1 vccd1 _20089_/Q sky130_fd_sc_hd__dfxtp_1
X_12980_ _13575_/C _14110_/C vssd1 vssd1 vccd1 vccd1 _13140_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11931_ _19391_/Q _12085_/A2 _11929_/X _11641_/S _11930_/X vssd1 vssd1 vccd1 vccd1
+ _11931_/X sky130_fd_sc_hd__o221a_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_501 _20621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_512 input220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _19412_/Q _17934_/A1 _14650_/S vssd1 vssd1 vccd1 vccd1 _19412_/D sky130_fd_sc_hd__mux2_1
XANTENNA_523 _13584_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _11949_/S _11862_/B vssd1 vssd1 vccd1 vccd1 _11862_/Y sky130_fd_sc_hd__nand2_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_534 _15323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_545 _12513_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_556 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13601_ _12664_/C _13600_/X _12982_/B vssd1 vssd1 vccd1 vccd1 _13603_/A sky130_fd_sc_hd__a21oi_1
XFILLER_261_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10813_ _10127_/A _10808_/Y _10812_/X _10806_/X vssd1 vssd1 vccd1 vccd1 _10813_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_567 _13666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _19347_/Q _17199_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19347_/D sky130_fd_sc_hd__mux2_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_578 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ _11764_/Y _11765_/X _11789_/X _15551_/A _11792_/X vssd1 vssd1 vccd1 vccd1
+ _11793_/X sky130_fd_sc_hd__a2111o_2
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_589 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16320_ _19715_/Q _16322_/C _16319_/Y vssd1 vssd1 vccd1 vccd1 _19715_/D sky130_fd_sc_hd__o21a_1
X_13532_ _13064_/C _13055_/Y _13062_/Y vssd1 vssd1 vccd1 vccd1 _13532_/Y sky130_fd_sc_hd__a21oi_1
X_10744_ _12383_/A _10744_/B vssd1 vssd1 vccd1 vccd1 _10744_/X sky130_fd_sc_hd__or2_1
XFILLER_213_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16251_ _19667_/Q _17925_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19667_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13463_ split3/A _13463_/B _13463_/C vssd1 vssd1 vccd1 vccd1 _13463_/X sky130_fd_sc_hd__and3_4
X_10675_ _19274_/Q _20061_/Q _12219_/S vssd1 vssd1 vccd1 vccd1 _10675_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15202_ _19705_/Q _15201_/X _15454_/S vssd1 vssd1 vccd1 vccd1 _15202_/X sky130_fd_sc_hd__mux2_2
X_12414_ _12412_/X _12413_/X _12414_/S vssd1 vssd1 vccd1 vccd1 _12414_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16182_ _19615_/Q _15861_/X _16190_/S vssd1 vssd1 vccd1 vccd1 _16183_/B sky130_fd_sc_hd__mux2_1
X_13394_ _13021_/Y _13394_/B vssd1 vssd1 vccd1 vccd1 _13395_/B sky130_fd_sc_hd__nand2b_1
XFILLER_126_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15133_ _15133_/A _15133_/B vssd1 vssd1 vccd1 vccd1 _15133_/X sky130_fd_sc_hd__and2_1
XFILLER_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ _12343_/X _12344_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _12345_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19941_ _20472_/CLK _19941_/D vssd1 vssd1 vccd1 vccd1 _19941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15064_ _15063_/X _15060_/X _15292_/S vssd1 vssd1 vccd1 vccd1 _15064_/X sky130_fd_sc_hd__mux2_1
X_12276_ _11201_/A _12258_/X _12275_/X vssd1 vssd1 vccd1 vccd1 _12276_/X sky130_fd_sc_hd__o21a_2
XFILLER_175_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14015_ _19204_/Q _14089_/C _14039_/S vssd1 vssd1 vccd1 vccd1 _14015_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11227_ input123/X input158/X _11241_/S vssd1 vssd1 vccd1 vccd1 _11227_/X sky130_fd_sc_hd__mux2_8
X_19872_ _20468_/CLK _19872_/D vssd1 vssd1 vccd1 vccd1 _19872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_268_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18823_ _18830_/A _18823_/B vssd1 vssd1 vccd1 vccd1 _18823_/Y sky130_fd_sc_hd__nand2_1
X_11158_ _11353_/C1 _11156_/X _11157_/X _11359_/S vssd1 vssd1 vccd1 vccd1 _11158_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_150_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_156_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21026_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_95_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10109_ _12107_/A1 _17898_/A1 _10108_/X _12194_/B2 vssd1 vssd1 vccd1 vccd1 _15504_/A
+ sky130_fd_sc_hd__a22o_2
X_11089_ _19625_/Q _11090_/S _11072_/X _11094_/S vssd1 vssd1 vccd1 vccd1 _11089_/X
+ sky130_fd_sc_hd__o211a_1
X_15966_ _20910_/Q _16043_/A2 _16043_/B1 _15965_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _15966_/X sky130_fd_sc_hd__a221o_1
X_18754_ _18754_/A _18754_/B vssd1 vssd1 vccd1 vccd1 _20977_/D sky130_fd_sc_hd__and2_1
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput270 partID[15] vssd1 vssd1 vccd1 vccd1 input270/X sky130_fd_sc_hd__clkbuf_2
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput281 versionID[1] vssd1 vssd1 vccd1 vccd1 _15081_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14917_ _14917_/A _16711_/A vssd1 vssd1 vccd1 vccd1 _14917_/Y sky130_fd_sc_hd__nor2_1
X_17705_ _20489_/Q _17705_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20489_/D sky130_fd_sc_hd__mux2_1
XFILLER_252_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18685_ _18973_/A _18685_/B vssd1 vssd1 vccd1 vccd1 _20944_/D sky130_fd_sc_hd__nor2_1
X_15897_ _19552_/Q _15980_/A2 _15895_/X _15896_/X _16185_/A vssd1 vssd1 vccd1 vccd1
+ _19552_/D sky130_fd_sc_hd__o221a_1
XFILLER_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17636_ _20392_/Q _17947_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20392_/D sky130_fd_sc_hd__mux2_1
X_14848_ _14844_/X _14847_/X _15170_/A vssd1 vssd1 vccd1 vccd1 _14848_/X sky130_fd_sc_hd__mux2_1
XFILLER_251_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17567_ _20327_/Q _17806_/A1 _17567_/S vssd1 vssd1 vccd1 vccd1 _20327_/D sky130_fd_sc_hd__mux2_1
XFILLER_211_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14779_ _19514_/Q _14797_/B vssd1 vssd1 vccd1 vccd1 _14779_/X sky130_fd_sc_hd__or2_1
XFILLER_189_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19306_ _20690_/CLK _19306_/D vssd1 vssd1 vccd1 vccd1 _19306_/Q sky130_fd_sc_hd__dfxtp_1
X_16518_ _19825_/Q _17111_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19825_/D sky130_fd_sc_hd__mux2_1
X_17498_ _20284_/Q _17502_/B vssd1 vssd1 vccd1 vccd1 _17498_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16449_ _19763_/Q _16450_/C _19764_/Q vssd1 vssd1 vccd1 vccd1 _16451_/B sky130_fd_sc_hd__a21oi_1
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19237_ _19246_/CLK _19237_/D vssd1 vssd1 vccd1 vccd1 _19237_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19168_ _19560_/CLK _19168_/D vssd1 vssd1 vccd1 vccd1 _19168_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_164_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18119_ _20782_/Q _18122_/C vssd1 vssd1 vccd1 vccd1 _18120_/B sky130_fd_sc_hd__and2_1
XFILLER_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19099_ _19620_/CLK _19099_/D vssd1 vssd1 vccd1 vccd1 _19099_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_172_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20012_ _20014_/CLK _20012_/D vssd1 vssd1 vccd1 vccd1 _20012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09823_ _12073_/A1 _09812_/X _09815_/X _09822_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1
+ _09823_/X sky130_fd_sc_hd__a311o_1
XFILLER_235_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09754_ _19646_/Q _19952_/Q _19290_/Q _20077_/Q _11932_/S0 _12003_/C vssd1 vssd1
+ vccd1 vccd1 _09754_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09685_ _09676_/Y _12039_/A1 split7/A vssd1 vssd1 vccd1 vccd1 _09685_/X sky130_fd_sc_hd__a21o_4
XFILLER_215_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20914_ _20980_/CLK _20914_/D vssd1 vssd1 vccd1 vccd1 _20914_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20845_ _21043_/CLK _20845_/D vssd1 vssd1 vccd1 vccd1 _20845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20776_ _21029_/CLK _20776_/D vssd1 vssd1 vccd1 vccd1 _20776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10460_ _19569_/Q _10459_/X _11240_/S vssd1 vssd1 vccd1 vccd1 _10460_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10391_ _09829_/A _20376_/Q _20440_/Q _10397_/S _12100_/B1 vssd1 vssd1 vccd1 vccd1
+ _10391_/X sky130_fd_sc_hd__a221o_1
XFILLER_151_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12130_ _20553_/Q _12139_/S vssd1 vssd1 vccd1 vccd1 _12130_/X sky130_fd_sc_hd__or2_1
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ _20651_/Q _20615_/Q _12070_/S vssd1 vssd1 vccd1 vccd1 _12061_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1903 _14482_/A vssd1 vssd1 vccd1 vccd1 _18730_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ _11012_/A _11012_/B _11012_/C vssd1 vssd1 vccd1 vccd1 _11012_/X sky130_fd_sc_hd__or3_2
Xfanout1914 _18352_/C1 vssd1 vssd1 vccd1 vccd1 _18714_/A sky130_fd_sc_hd__buf_2
Xfanout1925 _14070_/C1 vssd1 vssd1 vccd1 vccd1 _16143_/A sky130_fd_sc_hd__clkbuf_8
Xfanout1936 _18396_/A vssd1 vssd1 vccd1 vccd1 _18700_/A sky130_fd_sc_hd__clkbuf_4
Xfanout1947 _14104_/C1 vssd1 vssd1 vccd1 vccd1 _14088_/C1 sky130_fd_sc_hd__buf_4
Xfanout1958 _18416_/A vssd1 vssd1 vccd1 vccd1 _18414_/A sky130_fd_sc_hd__buf_4
Xfanout960 _11397_/A2 vssd1 vssd1 vccd1 vccd1 _17058_/A1 sky130_fd_sc_hd__clkbuf_2
X_15820_ _14843_/S _15373_/X _15376_/Y _15258_/A vssd1 vssd1 vccd1 vccd1 _15820_/X
+ sky130_fd_sc_hd__o22a_2
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout971 _17095_/A1 vssd1 vssd1 vccd1 vccd1 _17163_/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout1969 _13595_/A vssd1 vssd1 vccd1 vccd1 _17532_/A sky130_fd_sc_hd__buf_8
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout982 _10207_/X vssd1 vssd1 vccd1 vccd1 _17901_/A1 sky130_fd_sc_hd__buf_6
XFILLER_265_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout993 _17005_/A2 vssd1 vssd1 vccd1 vccd1 _16996_/B1 sky130_fd_sc_hd__buf_4
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _20806_/Q _15941_/A2 _15744_/X _15941_/B2 _15750_/X vssd1 vssd1 vccd1 vccd1
+ _15751_/X sky130_fd_sc_hd__a221o_1
X_12963_ _16719_/A _18136_/A _16710_/A _12963_/D vssd1 vssd1 vccd1 vccd1 _14121_/A
+ sky130_fd_sc_hd__or4_4
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14702_ _19461_/Q _17708_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19461_/D sky130_fd_sc_hd__mux2_1
XFILLER_234_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18470_ _18760_/B _18471_/B vssd1 vssd1 vccd1 vccd1 _18470_/Y sky130_fd_sc_hd__nor2_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _11513_/S _11913_/X _11912_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _11914_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_73_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15682_ _11730_/B _15984_/A2 _15984_/B1 _13166_/B _15890_/A vssd1 vssd1 vccd1 vccd1
+ _15682_/X sky130_fd_sc_hd__a221o_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_320 _13479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12894_ _13209_/B _12894_/B vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__and2_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 _20260_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17421_/A _17421_/B vssd1 vssd1 vccd1 vccd1 _17421_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_342 _19502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14633_ _19397_/Q _17917_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19397_/D sky130_fd_sc_hd__mux2_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11845_ _11851_/A _19921_/Q _12165_/S _20046_/Q vssd1 vssd1 vccd1 vccd1 _11845_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_353 _17178_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_364 _12708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_375 _18765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_386 _15387_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _20224_/Q _17356_/A2 _17362_/B1 _20273_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17352_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_397 _16000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14564_ _19091_/Q _16454_/B vssd1 vssd1 vccd1 vccd1 _17744_/A sky130_fd_sc_hd__or2_4
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _15264_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _19709_/Q _16306_/C _18054_/A vssd1 vssd1 vccd1 vccd1 _16303_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13515_ _19219_/Q _13499_/A _13514_/Y vssd1 vssd1 vccd1 vccd1 _13515_/X sky130_fd_sc_hd__o21a_1
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17283_ _20200_/Q _17331_/A2 _17281_/X _17282_/X _17331_/C1 vssd1 vssd1 vccd1 vccd1
+ _20200_/D sky130_fd_sc_hd__o221a_1
X_10727_ _19565_/Q _11061_/A _09659_/X _10726_/Y vssd1 vssd1 vccd1 vccd1 _10727_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14495_ _19273_/Q _17683_/A1 _14519_/S vssd1 vssd1 vccd1 vccd1 _19273_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19022_ _18250_/Y _19048_/A2 _19048_/B1 _12552_/D _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19022_/X sky130_fd_sc_hd__a221o_1
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16234_ _16240_/A1 _16233_/X _19695_/D vssd1 vssd1 vccd1 vccd1 _19655_/D sky130_fd_sc_hd__o21a_2
X_13446_ _13463_/B _13446_/B vssd1 vssd1 vccd1 vccd1 _16232_/B sky130_fd_sc_hd__nand2_8
X_10658_ _20029_/Q _12219_/S vssd1 vssd1 vccd1 vccd1 _10658_/X sky130_fd_sc_hd__or2_1
XFILLER_139_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16165_ _19606_/Q _16164_/B _16164_/Y _16165_/C1 vssd1 vssd1 vccd1 vccd1 _19606_/D
+ sky130_fd_sc_hd__o211a_1
X_13377_ _13377_/A _13377_/B vssd1 vssd1 vccd1 vccd1 _13377_/Y sky130_fd_sc_hd__nor2_2
X_10589_ _10587_/X _10588_/X _12056_/S vssd1 vssd1 vccd1 vccd1 _10589_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15116_ _11137_/A _15113_/X _15114_/Y _15115_/Y _15545_/A vssd1 vssd1 vccd1 vccd1
+ _15116_/X sky130_fd_sc_hd__o221a_1
X_12328_ _11012_/A _12326_/X _12327_/X vssd1 vssd1 vccd1 vccd1 _12328_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_86_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16096_ _10116_/X _16126_/A2 _16095_/X vssd1 vssd1 vccd1 vccd1 _19572_/D sky130_fd_sc_hd__o21a_1
XFILLER_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19924_ _20438_/CLK _19924_/D vssd1 vssd1 vccd1 vccd1 _19924_/Q sky130_fd_sc_hd__dfxtp_1
X_15047_ _14842_/X _14846_/X _15062_/S vssd1 vssd1 vccd1 vccd1 _15170_/B sky130_fd_sc_hd__mux2_1
X_12259_ _20147_/Q _20115_/Q _12428_/S vssd1 vssd1 vccd1 vccd1 _12259_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19855_ _20017_/CLK _19855_/D vssd1 vssd1 vccd1 vccd1 _19855_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18806_ _20986_/Q _18819_/B vssd1 vssd1 vccd1 vccd1 _18806_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19786_ _20712_/CLK _19786_/D vssd1 vssd1 vccd1 vccd1 _19786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16998_ _17008_/A1 _16997_/X _17008_/B1 vssd1 vssd1 vccd1 vccd1 _16998_/Y sky130_fd_sc_hd__o21ai_2
X_18737_ _20969_/Q _18275_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18738_/B sky130_fd_sc_hd__mux2_1
XFILLER_271_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15949_ _15949_/A _15949_/B vssd1 vssd1 vccd1 vccd1 _15949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18668_ _18544_/X _18684_/A2 _18666_/Y _18667_/Y vssd1 vssd1 vccd1 vccd1 _18669_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17619_ _20375_/Q _17687_/A1 _17623_/S vssd1 vssd1 vccd1 vccd1 _20375_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18599_ _20923_/Q _18619_/B vssd1 vssd1 vccd1 vccd1 _18599_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_53_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20467_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20630_ _20630_/CLK _20630_/D vssd1 vssd1 vccd1 vccd1 _20630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20561_ _20561_/CLK _20561_/D vssd1 vssd1 vccd1 vccd1 _20561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20492_ _20687_/CLK _20492_/D vssd1 vssd1 vccd1 vccd1 _20492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21044_ _21044_/CLK _21044_/D vssd1 vssd1 vccd1 vccd1 _21044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09806_ _09791_/X _09792_/X _09806_/S vssd1 vssd1 vccd1 vccd1 _09806_/X sky130_fd_sc_hd__mux2_1
XFILLER_275_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09737_ _19165_/Q _13863_/A vssd1 vssd1 vccd1 vccd1 _09737_/Y sky130_fd_sc_hd__nand2_2
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09668_ _09680_/B _09680_/C _09638_/Y vssd1 vssd1 vccd1 vccd1 _09678_/C sky130_fd_sc_hd__a21oi_1
XFILLER_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09599_ _16454_/A _16454_/B vssd1 vssd1 vccd1 vccd1 _17850_/A sky130_fd_sc_hd__nand2b_4
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _12192_/A1 _11619_/X _11623_/X _11629_/X vssd1 vssd1 vccd1 vccd1 _11646_/A
+ sky130_fd_sc_hd__a31o_1
X_20828_ _21022_/CLK _20828_/D vssd1 vssd1 vccd1 vccd1 _20828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ _09986_/A _20038_/Q _19913_/Q _09928_/S vssd1 vssd1 vccd1 vccd1 _11561_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20759_ _20759_/CLK _20759_/D vssd1 vssd1 vccd1 vccd1 _20759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ _13300_/A _13300_/B _13300_/C vssd1 vssd1 vccd1 vccd1 _13300_/X sky130_fd_sc_hd__and3_1
X_10512_ _09507_/A _10510_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14280_ _19510_/Q _14281_/B vssd1 vssd1 vccd1 vccd1 _14280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11492_ _12194_/A1 _17937_/A1 _11491_/X _12194_/B2 vssd1 vssd1 vccd1 vccd1 _15659_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_155_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13231_ _19240_/Q _13231_/B vssd1 vssd1 vccd1 vccd1 _13231_/X sky130_fd_sc_hd__xor2_1
X_10443_ _11266_/A1 _19908_/Q _10324_/S _20033_/Q vssd1 vssd1 vccd1 vccd1 _10443_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13162_ _13162_/A _13162_/B vssd1 vssd1 vccd1 vccd1 _13420_/B sky130_fd_sc_hd__nand2_2
X_10374_ input117/X input153/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10374_/X sky130_fd_sc_hd__mux2_8
XFILLER_124_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12113_ _11804_/A _11804_/B _12112_/X vssd1 vssd1 vccd1 vccd1 _12202_/A sky130_fd_sc_hd__a21o_2
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17970_ _20727_/Q _17971_/C _20728_/Q vssd1 vssd1 vccd1 vccd1 _17972_/B sky130_fd_sc_hd__a21oi_1
X_13093_ _20947_/Q _18472_/B _20946_/Q vssd1 vssd1 vccd1 vccd1 _13305_/B sky130_fd_sc_hd__or3b_4
XFILLER_269_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1700 _12254_/A vssd1 vssd1 vccd1 vccd1 _12337_/A sky130_fd_sc_hd__buf_6
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16921_ _20418_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16921_/X sky130_fd_sc_hd__a21o_2
X_12044_ _20583_/Q _12044_/B vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__or2_1
XFILLER_278_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1711 _12270_/B1 vssd1 vssd1 vccd1 vccd1 _11212_/S sky130_fd_sc_hd__buf_6
XFILLER_266_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1722 _10581_/A1 vssd1 vssd1 vccd1 vccd1 _12051_/A1 sky130_fd_sc_hd__buf_6
Xfanout1733 _12312_/A1 vssd1 vssd1 vccd1 vccd1 _12230_/A1 sky130_fd_sc_hd__buf_6
Xfanout1744 _12059_/A1 vssd1 vssd1 vccd1 vccd1 _11981_/C1 sky130_fd_sc_hd__buf_8
Xfanout1755 _14042_/S vssd1 vssd1 vccd1 vccd1 _14039_/S sky130_fd_sc_hd__clkbuf_4
X_19640_ _20075_/CLK _19640_/D vssd1 vssd1 vccd1 vccd1 _19640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16852_ _20410_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16852_/X sky130_fd_sc_hd__a21o_1
Xfanout1766 _09488_/A vssd1 vssd1 vccd1 vccd1 _13205_/A sky130_fd_sc_hd__buf_6
XFILLER_78_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1777 _17441_/A vssd1 vssd1 vccd1 vccd1 _17446_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_281_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1788 _18209_/A1 vssd1 vssd1 vccd1 vccd1 _18213_/B sky130_fd_sc_hd__buf_12
Xfanout790 _12857_/B vssd1 vssd1 vccd1 vccd1 _12916_/A2 sky130_fd_sc_hd__buf_4
X_15803_ _20968_/Q _16045_/A2 _16016_/S _20840_/Q _15802_/X vssd1 vssd1 vccd1 vccd1
+ _15803_/X sky130_fd_sc_hd__a221o_1
Xfanout1799 _16769_/S vssd1 vssd1 vccd1 vccd1 _16799_/S sky130_fd_sc_hd__clkbuf_8
X_19571_ _20341_/CLK _19571_/D vssd1 vssd1 vccd1 vccd1 _19571_/Q sky130_fd_sc_hd__dfxtp_1
X_16783_ _19966_/Q _16849_/A _16782_/Y _16451_/A vssd1 vssd1 vccd1 vccd1 _19966_/D
+ sky130_fd_sc_hd__a211o_1
X_13995_ _19165_/Q _19050_/S _14043_/B1 _13994_/X _16129_/B1 vssd1 vssd1 vccd1 vccd1
+ _19165_/D sky130_fd_sc_hd__o221a_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15734_ _15734_/A _15734_/B _15981_/B vssd1 vssd1 vccd1 vccd1 _15734_/X sky130_fd_sc_hd__and3_1
X_18522_ _18891_/A _18522_/B vssd1 vssd1 vccd1 vccd1 _20900_/D sky130_fd_sc_hd__nor2_1
X_12946_ _16711_/A _12946_/B _16720_/B _16720_/C vssd1 vssd1 vccd1 vccd1 _16719_/A
+ sky130_fd_sc_hd__or4_2
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _20881_/Q _18315_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18454_/B sky130_fd_sc_hd__mux2_1
X_15665_ _20899_/Q _15937_/A2 _15994_/B1 _15664_/X _15937_/C1 vssd1 vssd1 vccd1 vccd1
+ _15665_/X sky130_fd_sc_hd__a221o_1
XFILLER_244_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12877_ _12911_/A _12877_/B vssd1 vssd1 vccd1 vccd1 _12878_/B sky130_fd_sc_hd__nor2_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_150 _13755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _13780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _19380_/Q _17866_/A1 _14628_/S vssd1 vssd1 vccd1 vccd1 _19380_/D sky130_fd_sc_hd__mux2_1
X_17404_ _20257_/Q _17236_/A _17442_/A vssd1 vssd1 vccd1 vccd1 _17404_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 _19110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ _20649_/Q _20613_/Q _12139_/S vssd1 vssd1 vccd1 vccd1 _11828_/X sky130_fd_sc_hd__mux2_1
XANTENNA_183 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18384_ _20847_/Q _18387_/B _18383_/Y _18754_/A vssd1 vssd1 vccd1 vccd1 _20847_/D
+ sky130_fd_sc_hd__o211a_1
X_15596_ _20737_/Q _16041_/A2 _16041_/B1 _20769_/Q vssd1 vssd1 vccd1 vccd1 _15596_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_194 _19542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17402_/A _17335_/B _17336_/B vssd1 vssd1 vccd1 vccd1 _17335_/X sky130_fd_sc_hd__and3_4
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _19317_/Q _17099_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19317_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11759_ _11758_/B _15734_/A _13415_/A vssd1 vssd1 vccd1 vccd1 _15763_/B sky130_fd_sc_hd__a21o_1
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17266_ _17266_/A _17275_/B _17269_/C vssd1 vssd1 vccd1 vccd1 _17266_/X sky130_fd_sc_hd__and3_1
XFILLER_146_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14478_ _18718_/A _14478_/B vssd1 vssd1 vccd1 vccd1 _19263_/D sky130_fd_sc_hd__and2_1
X_19005_ _21022_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _19005_/X sky130_fd_sc_hd__or2_1
X_16217_ _19640_/Q _17869_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19640_/D sky130_fd_sc_hd__mux2_1
X_13429_ _15816_/A _13429_/B _13414_/Y vssd1 vssd1 vccd1 vccd1 _13430_/A sky130_fd_sc_hd__or3b_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17197_ _20161_/Q _17931_/A1 _17215_/S vssd1 vssd1 vccd1 vccd1 _20161_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16148_ _16794_/B _16196_/S vssd1 vssd1 vccd1 vccd1 _16148_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_171_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20969_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_100_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20757_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16079_ _16079_/A _16079_/B vssd1 vssd1 vccd1 vccd1 _16079_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19907_ _20657_/CLK _19907_/D vssd1 vssd1 vccd1 vccd1 _19907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19838_ _19978_/CLK _19838_/D vssd1 vssd1 vccd1 vccd1 _19838_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 coreIndex[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
X_19769_ _20565_/CLK _19769_/D vssd1 vssd1 vccd1 vccd1 _19769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09522_ _09522_/A vssd1 vssd1 vccd1 vccd1 _09522_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20613_ _20681_/CLK _20613_/D vssd1 vssd1 vccd1 vccd1 _20613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20544_ _20676_/CLK _20544_/D vssd1 vssd1 vccd1 vccd1 _20544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20475_ _20703_/CLK _20475_/D vssd1 vssd1 vccd1 vccd1 _20475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput360 _13652_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[4] sky130_fd_sc_hd__buf_4
Xoutput371 _09531_/X vssd1 vssd1 vccd1 vccd1 core_wb_we_o sky130_fd_sc_hd__buf_4
Xoutput382 _13806_/X vssd1 vssd1 vccd1 vccd1 din0[15] sky130_fd_sc_hd__buf_4
Xfanout1007 _14903_/Y vssd1 vssd1 vccd1 vccd1 _15314_/B sky130_fd_sc_hd__buf_4
X_10090_ _09507_/A _10089_/X _10088_/X vssd1 vssd1 vccd1 vccd1 _10090_/X sky130_fd_sc_hd__o21a_1
XFILLER_160_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput393 _13816_/X vssd1 vssd1 vccd1 vccd1 din0[25] sky130_fd_sc_hd__buf_4
Xfanout1018 _18785_/A2 vssd1 vssd1 vccd1 vccd1 _18864_/A2 sky130_fd_sc_hd__buf_2
Xfanout1029 _15527_/Y vssd1 vssd1 vccd1 vccd1 _15976_/B2 sky130_fd_sc_hd__buf_4
XFILLER_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21027_ _21027_/CLK _21027_/D vssd1 vssd1 vccd1 vccd1 _21027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12800_ _12804_/B _12800_/B vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__or2_1
X_13780_ _13780_/A _13780_/B vssd1 vssd1 vccd1 vccd1 _13780_/X sky130_fd_sc_hd__and2_1
XFILLER_262_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10992_ _11336_/A _11258_/A1 _20121_/Q _11345_/S vssd1 vssd1 vccd1 vccd1 _10992_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_28_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _15504_/A _12731_/B vssd1 vssd1 vccd1 vccd1 _12731_/Y sky130_fd_sc_hd__nand2_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15450_ _20860_/Q _15449_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15450_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12662_ _12662_/A _12662_/B _12662_/C vssd1 vssd1 vccd1 vccd1 _13501_/B sky130_fd_sc_hd__and3_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14401_ _19522_/Q _14406_/B vssd1 vssd1 vccd1 vccd1 _14402_/B sky130_fd_sc_hd__nand2_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _12157_/A1 _17905_/A1 _11609_/X _12153_/B1 vssd1 vssd1 vccd1 vccd1 _13717_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15381_ _19710_/Q _15475_/A2 _15475_/B1 _19742_/Q vssd1 vssd1 vccd1 vccd1 _15381_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_212_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12593_ _19864_/Q _19863_/Q vssd1 vssd1 vccd1 vccd1 _16598_/A sky130_fd_sc_hd__or2_4
XFILLER_129_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17120_ _20088_/Q _17922_/A1 _17132_/S vssd1 vssd1 vccd1 vccd1 _20088_/D sky130_fd_sc_hd__mux2_1
X_14332_ _19515_/Q _14332_/B vssd1 vssd1 vccd1 vccd1 _14333_/C sky130_fd_sc_hd__xnor2_1
XFILLER_129_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11544_ _09986_/C _11543_/X _12006_/S vssd1 vssd1 vccd1 vccd1 _11544_/X sky130_fd_sc_hd__a21o_1
XFILLER_183_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _20023_/Q _17051_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20023_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _14262_/A _14259_/B _14262_/X vssd1 vssd1 vccd1 vccd1 _14263_/X sky130_fd_sc_hd__a21bo_1
XFILLER_184_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11475_ _19383_/Q _20674_/Q _12165_/S vssd1 vssd1 vccd1 vccd1 _11475_/X sky130_fd_sc_hd__mux2_1
X_16002_ _16002_/A1 _15988_/Y _16002_/B1 vssd1 vssd1 vccd1 vccd1 _16002_/Y sky130_fd_sc_hd__a21oi_1
X_13214_ _13002_/A _13209_/Y _13210_/X _13213_/X vssd1 vssd1 vccd1 vccd1 _13218_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10426_ _20376_/Q _20440_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _10426_/X sky130_fd_sc_hd__mux2_1
X_14194_ _14204_/A _16068_/B _14194_/C vssd1 vssd1 vccd1 vccd1 _14194_/X sky130_fd_sc_hd__or3_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13145_ _13145_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _13495_/B sky130_fd_sc_hd__nand2_2
XFILLER_152_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10357_ _19812_/Q _11291_/A2 _10355_/X _11291_/B2 _10356_/X vssd1 vssd1 vccd1 vccd1
+ _10357_/X sky130_fd_sc_hd__o221a_1
XFILLER_3_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _20722_/Q _21044_/Q vssd1 vssd1 vccd1 vccd1 _17955_/B sky130_fd_sc_hd__and2b_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _20963_/Q _20897_/Q _13340_/A vssd1 vssd1 vccd1 vccd1 _13076_/X sky130_fd_sc_hd__a21o_1
XFILLER_285_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10288_ _09672_/A _14038_/A2 _10287_/X _11228_/B1 _19861_/Q vssd1 vssd1 vccd1 vccd1
+ _10288_/X sky130_fd_sc_hd__o32a_1
XFILLER_250_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16904_ _19979_/Q _16876_/A _16903_/Y _18126_/A vssd1 vssd1 vccd1 vccd1 _19979_/D
+ sky130_fd_sc_hd__a211o_1
X_12027_ _12023_/X _12026_/X _12828_/A vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__mux2_1
Xfanout1530 _10425_/S vssd1 vssd1 vccd1 vccd1 _12070_/S sky130_fd_sc_hd__buf_6
XFILLER_266_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1541 _10137_/C vssd1 vssd1 vccd1 vccd1 _10986_/B sky130_fd_sc_hd__buf_6
XFILLER_39_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1552 fanout1556/X vssd1 vssd1 vccd1 vccd1 _12219_/S sky130_fd_sc_hd__clkbuf_4
X_17884_ _17884_/A _17918_/A vssd1 vssd1 vccd1 vccd1 _17885_/C sky130_fd_sc_hd__nor2_1
Xfanout1563 _11161_/S vssd1 vssd1 vccd1 vccd1 _12313_/S sky130_fd_sc_hd__clkbuf_4
Xfanout1574 _09624_/Y vssd1 vssd1 vccd1 vccd1 _12399_/C1 sky130_fd_sc_hd__buf_6
X_19623_ _20657_/CLK _19623_/D vssd1 vssd1 vccd1 vccd1 _19623_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1585 _09622_/Y vssd1 vssd1 vccd1 vccd1 _11597_/C1 sky130_fd_sc_hd__buf_8
X_16835_ _19226_/Q _17003_/B _16964_/B1 _19095_/Q _16834_/X vssd1 vssd1 vccd1 vccd1
+ _16835_/X sky130_fd_sc_hd__o221a_1
XFILLER_254_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1596 _09621_/Y vssd1 vssd1 vccd1 vccd1 _11600_/C1 sky130_fd_sc_hd__buf_6
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19554_ _19617_/CLK _19554_/D vssd1 vssd1 vccd1 vccd1 _19554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_280_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13978_ _14002_/A1 _13978_/A2 _10458_/X _14002_/B1 _19841_/Q vssd1 vssd1 vccd1 vccd1
+ _14065_/C sky130_fd_sc_hd__o32a_2
X_16766_ _19219_/Q _16996_/A2 _16713_/X _16765_/X vssd1 vssd1 vccd1 vccd1 _16766_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18505_ _18616_/B _18505_/B vssd1 vssd1 vccd1 vccd1 _18505_/X sky130_fd_sc_hd__or2_2
X_12929_ _13466_/B _14117_/B vssd1 vssd1 vccd1 vccd1 _12930_/B sky130_fd_sc_hd__nor2_8
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15717_ _20869_/Q _16018_/A2 fanout819/X vssd1 vssd1 vccd1 vccd1 _15717_/X sky130_fd_sc_hd__o21ba_1
XFILLER_262_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19485_ _20712_/CLK _19485_/D vssd1 vssd1 vccd1 vccd1 _19485_/Q sky130_fd_sc_hd__dfxtp_1
X_16697_ _19952_/Q _17107_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19952_/D sky130_fd_sc_hd__mux2_1
XFILLER_234_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18436_ _18734_/A _18436_/B vssd1 vssd1 vccd1 vccd1 _20872_/D sky130_fd_sc_hd__and2_1
XFILLER_34_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15648_ _15977_/A1 _12855_/X _15647_/X _15703_/B2 vssd1 vssd1 vccd1 vccd1 _15650_/A
+ sky130_fd_sc_hd__o22a_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18367_ _18529_/B _18385_/B vssd1 vssd1 vccd1 vccd1 _18367_/Y sky130_fd_sc_hd__nand2_1
X_15579_ _15610_/A1 _15065_/X _15610_/B1 vssd1 vssd1 vccd1 vccd1 _15654_/B sky130_fd_sc_hd__o21ai_4
XFILLER_203_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17318_ _20211_/Q _17321_/A2 _17305_/C _17317_/X _17330_/C1 vssd1 vssd1 vccd1 vccd1
+ _17318_/X sky130_fd_sc_hd__a221o_1
XFILLER_193_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18298_ _19555_/Q _18308_/B vssd1 vssd1 vccd1 vccd1 _18298_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_174_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17249_ _20188_/Q _17235_/Y _17279_/C1 vssd1 vssd1 vccd1 vccd1 _17249_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20260_ _20685_/CLK _20260_/D vssd1 vssd1 vccd1 vccd1 _20260_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_134_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20191_ _20428_/CLK _20191_/D vssd1 vssd1 vccd1 vccd1 _20191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ _12430_/S vssd1 vssd1 vccd1 vccd1 _09505_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_50 _16927_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 _17813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 _09607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20527_ _20686_/CLK _20527_/D vssd1 vssd1 vccd1 vccd1 _20527_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_83 _10714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_94 _12154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11260_ _11250_/X _11253_/X _11256_/X _11259_/X _12513_/C _09621_/A vssd1 vssd1 vccd1
+ vccd1 _11260_/X sky130_fd_sc_hd__mux4_2
X_20458_ _20491_/CLK _20458_/D vssd1 vssd1 vccd1 vccd1 _20458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10211_ _19880_/Q _19781_/Q _10217_/S vssd1 vssd1 vccd1 vccd1 _10211_/X sky130_fd_sc_hd__mux2_1
XFILLER_279_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11191_ _11191_/A _19303_/Q _11191_/C vssd1 vssd1 vccd1 vccd1 _11191_/X sky130_fd_sc_hd__or3_1
X_20389_ _21046_/A _20389_/D vssd1 vssd1 vccd1 vccd1 _20389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ _10140_/X _10141_/X _12377_/S vssd1 vssd1 vccd1 vccd1 _10142_/X sky130_fd_sc_hd__mux2_1
XFILLER_267_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14950_ _14950_/A _14950_/B vssd1 vssd1 vccd1 vccd1 _14973_/C sky130_fd_sc_hd__nand2_1
X_10073_ _12073_/A1 _10069_/X _10072_/X _12059_/C1 vssd1 vssd1 vccd1 vccd1 _10073_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13901_ _13902_/A _16133_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _13901_/X sky130_fd_sc_hd__and3_1
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14881_ _14881_/A _14881_/B vssd1 vssd1 vccd1 vccd1 _14881_/X sky130_fd_sc_hd__or2_1
XFILLER_263_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16620_ _19879_/Q _17657_/A1 _16620_/S vssd1 vssd1 vccd1 vccd1 _19879_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13832_ _20002_/Q split1/X _13786_/X _16279_/B vssd1 vssd1 vccd1 vccd1 _13832_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_90_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16551_ _16551_/A _16551_/B vssd1 vssd1 vccd1 vccd1 _19841_/D sky130_fd_sc_hd__or2_1
XFILLER_244_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13763_ _13684_/Y _13741_/B _13741_/Y _13685_/Y _13762_/X vssd1 vssd1 vccd1 vccd1
+ _13764_/B sky130_fd_sc_hd__o221a_4
X_10975_ _11239_/A1 _13969_/A2 _10974_/X _11228_/B1 _19834_/Q vssd1 vssd1 vccd1 vccd1
+ _16075_/A sky130_fd_sc_hd__o32ai_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12714_ _12709_/X _12711_/Y _12706_/Y _12707_/X vssd1 vssd1 vccd1 vccd1 _12714_/X
+ sky130_fd_sc_hd__a211o_1
X_15502_ _14843_/S _15499_/X _15501_/Y _15526_/B vssd1 vssd1 vccd1 vccd1 _15502_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_280_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19270_ _20379_/CLK _19270_/D vssd1 vssd1 vccd1 vccd1 _19270_/Q sky130_fd_sc_hd__dfxtp_1
X_16482_ _19791_/Q _17945_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19791_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13694_ _13694_/A _14878_/A _13694_/C vssd1 vssd1 vccd1 vccd1 _13694_/X sky130_fd_sc_hd__and3_2
X_18221_ _20798_/Q _18220_/Y _18311_/S vssd1 vssd1 vccd1 vccd1 _18222_/B sky130_fd_sc_hd__mux2_1
X_15433_ _15433_/A _15433_/B _15494_/B vssd1 vssd1 vccd1 vccd1 _15433_/X sky130_fd_sc_hd__and3_1
X_12645_ _12698_/B _12698_/C vssd1 vssd1 vccd1 vccd1 _12645_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_203_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18152_ _18163_/A _18152_/B _18152_/C vssd1 vssd1 vccd1 vccd1 _18152_/X sky130_fd_sc_hd__and3_1
X_15364_ _15258_/A _15359_/X _15363_/X _14843_/S vssd1 vssd1 vccd1 vccd1 _15365_/C
+ sky130_fd_sc_hd__o22a_2
XFILLER_8_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12576_ _12577_/A _12577_/B vssd1 vssd1 vccd1 vccd1 _12576_/Y sky130_fd_sc_hd__nor2_1
XFILLER_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17103_ _20073_/Q _17939_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20073_/D sky130_fd_sc_hd__mux2_1
X_14315_ _14325_/A _14315_/B _14323_/B vssd1 vssd1 vccd1 vccd1 _14315_/X sky130_fd_sc_hd__or3b_1
XFILLER_117_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18083_ _20768_/Q _18085_/C _18082_/Y vssd1 vssd1 vccd1 vccd1 _20768_/D sky130_fd_sc_hd__o21a_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11527_ _19283_/Q _20070_/Q _11527_/S vssd1 vssd1 vccd1 vccd1 _11527_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15295_ _15407_/S _15057_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _15295_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17034_ _20012_/Q input198/X _17040_/S vssd1 vssd1 vccd1 vccd1 _20012_/D sky130_fd_sc_hd__mux2_1
X_14246_ _19227_/Q _14256_/A2 _14245_/X _18352_/C1 vssd1 vssd1 vccd1 vccd1 _19227_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11458_ _19165_/Q _19914_/Q _12464_/C vssd1 vssd1 vccd1 vccd1 _11458_/X sky130_fd_sc_hd__and3_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10409_ _10409_/A _10409_/B vssd1 vssd1 vccd1 vccd1 _10409_/X sky130_fd_sc_hd__or2_1
Xclkbuf_3_4_0_wb_clk_i ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_14177_ _19500_/Q _14177_/B vssd1 vssd1 vccd1 vccd1 _14178_/B sky130_fd_sc_hd__nand2_2
X_11389_ _11387_/X _11388_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _11389_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13104_/B _13127_/Y _13334_/A vssd1 vssd1 vccd1 vccd1 _13128_/X sky130_fd_sc_hd__o21a_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_12__f_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19214_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18985_ _18985_/A _18985_/B vssd1 vssd1 vccd1 vccd1 _18985_/X sky130_fd_sc_hd__and2_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13059_ _20949_/Q _20883_/Q vssd1 vssd1 vccd1 vccd1 _13060_/D sky130_fd_sc_hd__or2_1
X_17936_ _20705_/Q _17936_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20705_/D sky130_fd_sc_hd__mux2_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1360 _14038_/B1 vssd1 vssd1 vccd1 vccd1 _14041_/B1 sky130_fd_sc_hd__buf_4
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1371 _12921_/X vssd1 vssd1 vccd1 vccd1 _14267_/A2 sky130_fd_sc_hd__buf_6
X_17867_ _20640_/Q _17901_/A1 _17883_/S vssd1 vssd1 vccd1 vccd1 _20640_/D sky130_fd_sc_hd__mux2_1
Xfanout1382 _11860_/B2 vssd1 vssd1 vccd1 vccd1 _09931_/S sky130_fd_sc_hd__buf_6
XFILLER_227_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1393 _09736_/Y vssd1 vssd1 vccd1 vccd1 _11848_/S0 sky130_fd_sc_hd__buf_4
XFILLER_253_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19606_ _19606_/CLK _19606_/D vssd1 vssd1 vccd1 vccd1 _19606_/Q sky130_fd_sc_hd__dfxtp_1
X_16818_ _16805_/X _16815_/Y _16817_/X _16932_/A1 vssd1 vssd1 vccd1 vccd1 _16818_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_253_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17798_ _20575_/Q _17938_/A1 _17806_/S vssd1 vssd1 vccd1 vccd1 _20575_/D sky130_fd_sc_hd__mux2_1
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19537_ _19620_/CLK _19537_/D vssd1 vssd1 vccd1 vccd1 _19537_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_207_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16749_ _16799_/S input70/X vssd1 vssd1 vccd1 vccd1 _16749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_146_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19468_ _20084_/CLK _19468_/D vssd1 vssd1 vccd1 vccd1 _19468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18419_ _20864_/Q _18230_/Y _18419_/S vssd1 vssd1 vccd1 vccd1 _18420_/B sky130_fd_sc_hd__mux2_1
XFILLER_195_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19399_ _20638_/CLK _19399_/D vssd1 vssd1 vccd1 vccd1 _19399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20312_ _20472_/CLK _20312_/D vssd1 vssd1 vccd1 vccd1 _20312_/Q sky130_fd_sc_hd__dfxtp_1
Xinput70 dout0[34] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_2
XFILLER_238_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput81 dout0[44] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__clkbuf_2
Xinput92 dout0[54] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20243_ _20296_/CLK _20243_/D vssd1 vssd1 vccd1 vccd1 _20243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20174_ _20481_/CLK _20174_/D vssd1 vssd1 vccd1 vccd1 _20174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09985_ _09986_/A _19917_/Q _12188_/S _20042_/Q vssd1 vssd1 vccd1 vccd1 _09985_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20715_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_232_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10760_ _12399_/A1 _10756_/X _10759_/X _12399_/C1 vssd1 vssd1 vccd1 vccd1 _10760_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_201_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10691_ _12411_/A _20500_/Q _12334_/S0 _20532_/Q vssd1 vssd1 vccd1 vccd1 _10691_/X
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_203_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20446_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12430_ _12426_/X _12429_/X _12430_/S vssd1 vssd1 vccd1 vccd1 _12430_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ _16037_/A vssd1 vssd1 vccd1 vccd1 _12361_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14100_ _19209_/Q _14104_/A2 _14099_/X _16127_/B1 vssd1 vssd1 vccd1 vccd1 _19209_/D
+ sky130_fd_sc_hd__o211a_1
X_11312_ _12433_/A1 _17852_/A1 _11311_/Y _09750_/Y vssd1 vssd1 vccd1 vccd1 _11312_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_154_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15080_ _20723_/Q _15445_/A2 _15445_/B1 _20755_/Q vssd1 vssd1 vccd1 vccd1 _15080_/X
+ sky130_fd_sc_hd__a22o_1
X_12292_ _10203_/A _11326_/A _11236_/B split7/X vssd1 vssd1 vccd1 vccd1 _12292_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14031_ _19177_/Q _14031_/A2 _14040_/B1 _14030_/X _16127_/B1 vssd1 vssd1 vccd1 vccd1
+ _19177_/D sky130_fd_sc_hd__o221a_1
X_11243_ _19575_/Q _11242_/X _11243_/S vssd1 vssd1 vccd1 vccd1 _11243_/X sky130_fd_sc_hd__mux2_4
XFILLER_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11174_ _19866_/Q _19767_/Q _11174_/S vssd1 vssd1 vccd1 vccd1 _11174_/X sky130_fd_sc_hd__mux2_1
XFILLER_267_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10125_ _10037_/Y _10124_/Y _09669_/X vssd1 vssd1 vccd1 vccd1 _10125_/X sky130_fd_sc_hd__a21o_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18770_ _18459_/Y _20980_/Q _18840_/B vssd1 vssd1 vccd1 vccd1 _18770_/X sky130_fd_sc_hd__mux2_1
XFILLER_283_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15982_ _15982_/A _15982_/B _15982_/C vssd1 vssd1 vccd1 vccd1 _15982_/X sky130_fd_sc_hd__or3_1
XFILLER_283_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17721_ _20502_/Q _17861_/A1 _17738_/S vssd1 vssd1 vccd1 vccd1 _20502_/D sky130_fd_sc_hd__mux2_1
X_14933_ _14945_/A _15314_/C vssd1 vssd1 vccd1 vccd1 _14933_/Y sky130_fd_sc_hd__nor2_8
X_10056_ _12060_/A1 _19474_/Q _19442_/Q _10428_/S vssd1 vssd1 vccd1 vccd1 _10056_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ _20438_/Q _17686_/A1 _17669_/S vssd1 vssd1 vccd1 vccd1 _20438_/D sky130_fd_sc_hd__mux2_1
XFILLER_264_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14864_ _15114_/B vssd1 vssd1 vccd1 vccd1 _14864_/Y sky130_fd_sc_hd__inv_2
XFILLER_251_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16603_ _19864_/Q _16597_/X _16602_/Y vssd1 vssd1 vccd1 vccd1 _19864_/D sky130_fd_sc_hd__o21a_1
XFILLER_223_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13815_ _13816_/A1 _13745_/B _13816_/B1 input231/X vssd1 vssd1 vccd1 vccd1 _13815_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17583_ _20341_/Q _17894_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20341_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14795_ _19522_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14795_/X sky130_fd_sc_hd__or2_1
X_19322_ _20677_/CLK _19322_/D vssd1 vssd1 vccd1 vccd1 _19322_/Q sky130_fd_sc_hd__dfxtp_1
X_16534_ _19833_/Q _16578_/A2 _16578_/B1 input32/X vssd1 vssd1 vccd1 vccd1 _16535_/B
+ sky130_fd_sc_hd__o22a_1
X_13746_ _11921_/Y _13742_/B _13663_/A vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__o21a_2
X_10958_ _19666_/Q _11377_/S vssd1 vssd1 vccd1 vccd1 _10958_/X sky130_fd_sc_hd__or2_1
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19253_ _20273_/CLK _19253_/D vssd1 vssd1 vccd1 vccd1 _19253_/Q sky130_fd_sc_hd__dfxtp_1
X_16465_ _19774_/Q _17928_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19774_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13677_ _13718_/A _13675_/Y _13676_/Y _13655_/A vssd1 vssd1 vccd1 vccd1 _13679_/B
+ sky130_fd_sc_hd__a211o_4
X_10889_ _10553_/B _10041_/Y _10888_/X _10028_/X vssd1 vssd1 vccd1 vccd1 _10889_/Y
+ sky130_fd_sc_hd__o211ai_2
X_18204_ _18209_/A1 _14208_/B _18203_/Y vssd1 vssd1 vccd1 vccd1 _18493_/B sky130_fd_sc_hd__o21ai_4
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15416_ _21021_/Q _20989_/Q _15508_/S vssd1 vssd1 vccd1 vccd1 _15416_/X sky130_fd_sc_hd__mux2_1
X_12628_ _12628_/A _12628_/B vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__or2_1
X_16396_ _19744_/Q _16396_/B vssd1 vssd1 vccd1 vccd1 _16402_/C sky130_fd_sc_hd__and2_2
X_19184_ _19621_/CLK _19184_/D vssd1 vssd1 vccd1 vccd1 _19184_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18135_ _18322_/A _18322_/C vssd1 vssd1 vccd1 vccd1 _18138_/A sky130_fd_sc_hd__nor2_1
X_15347_ _16002_/A1 _15331_/Y _15457_/B1 vssd1 vssd1 vccd1 vccd1 _15347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12559_ _13636_/A _13694_/A vssd1 vssd1 vccd1 vccd1 _12561_/A sky130_fd_sc_hd__and2_2
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15278_ _17254_/A _15277_/X _15452_/S vssd1 vssd1 vccd1 vccd1 _15278_/X sky130_fd_sc_hd__mux2_1
X_18066_ _20762_/Q _18069_/C _18056_/A vssd1 vssd1 vccd1 vccd1 _18066_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17017_ _19995_/Q input190/X _17849_/S vssd1 vssd1 vccd1 vccd1 _19995_/D sky130_fd_sc_hd__mux2_1
X_14229_ _19505_/Q _14229_/B vssd1 vssd1 vccd1 vccd1 _14230_/B sky130_fd_sc_hd__or2_1
XFILLER_256_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_78_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19577_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout608 _14567_/X vssd1 vssd1 vccd1 vccd1 _14594_/S sky130_fd_sc_hd__buf_6
XFILLER_259_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout619 _14398_/A2 vssd1 vssd1 vccd1 vccd1 _14438_/A2 sky130_fd_sc_hd__buf_6
XFILLER_99_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09770_ _19685_/Q _20173_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _09770_/X sky130_fd_sc_hd__mux2_1
X_18968_ _18968_/A _18968_/B vssd1 vssd1 vccd1 vccd1 _18968_/Y sky130_fd_sc_hd__nand2_4
XFILLER_239_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17919_ _17919_/A _17919_/B _17919_/C vssd1 vssd1 vccd1 vccd1 _17919_/X sky130_fd_sc_hd__and3_4
X_18899_ _19104_/Q _18954_/A2 _18974_/B1 _13428_/B vssd1 vssd1 vccd1 vccd1 _18899_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1190 _10561_/A vssd1 vssd1 vccd1 vccd1 _10385_/A sky130_fd_sc_hd__buf_4
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20930_ _20930_/CLK _20930_/D vssd1 vssd1 vccd1 vccd1 _20930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20861_ _20861_/CLK _20861_/D vssd1 vssd1 vccd1 vccd1 _20861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20792_ _20856_/CLK _20792_/D vssd1 vssd1 vccd1 vccd1 _20792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20226_ _20818_/CLK _20226_/D vssd1 vssd1 vccd1 vccd1 _20226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20157_ _20179_/CLK _20157_/D vssd1 vssd1 vccd1 vccd1 _20157_/Q sky130_fd_sc_hd__dfxtp_1
X_09968_ _20645_/Q _20609_/Q _12149_/S vssd1 vssd1 vccd1 vccd1 _09968_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20088_ _20559_/CLK _20088_/D vssd1 vssd1 vccd1 vccd1 _20088_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ _20043_/Q _19918_/Q _12149_/S vssd1 vssd1 vccd1 vccd1 _09899_/X sky130_fd_sc_hd__mux2_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _12003_/A _20682_/Q _12003_/C vssd1 vssd1 vccd1 vccd1 _11930_/X sky130_fd_sc_hd__or3_1
XFILLER_100_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_502 _20621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _11948_/A1 _11859_/X _11860_/X vssd1 vssd1 vccd1 vccd1 _11862_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_513 input220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_524 _13192_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_535 _18949_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_546 _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ _13600_/A _13600_/B vssd1 vssd1 vccd1 vccd1 _13600_/X sky130_fd_sc_hd__xor2_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _19564_/Q _11061_/A _09659_/X _10811_/Y vssd1 vssd1 vccd1 vccd1 _10812_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_557 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14580_ _19346_/Q _17932_/A1 _14599_/S vssd1 vssd1 vccd1 vccd1 _19346_/D sky130_fd_sc_hd__mux2_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_568 _13716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11792_ _11794_/C _11792_/B vssd1 vssd1 vccd1 vccd1 _11792_/X sky130_fd_sc_hd__and2_1
XFILLER_220_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_579 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13531_ _13589_/A1 _13526_/X _13527_/Y _13530_/X vssd1 vssd1 vccd1 vccd1 _13531_/X
+ sky130_fd_sc_hd__a31o_1
X_10743_ _10741_/X _10742_/X _12391_/S vssd1 vssd1 vccd1 vccd1 _10744_/B sky130_fd_sc_hd__mux2_1
XFILLER_213_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16250_ _19666_/Q _17647_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19666_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13462_ _16232_/B _13462_/B vssd1 vssd1 vccd1 vccd1 _13462_/X sky130_fd_sc_hd__or2_1
X_10674_ _12396_/A1 _19904_/Q _12391_/S _10658_/X vssd1 vssd1 vccd1 vccd1 _10674_/X
+ sky130_fd_sc_hd__o211a_1
X_15201_ _19737_/Q _15604_/A2 _15190_/X _15396_/A1 _15200_/X vssd1 vssd1 vccd1 vccd1
+ _15201_/X sky130_fd_sc_hd__a221o_1
X_12413_ _20427_/Q _20363_/Q _20655_/Q _20619_/Q _12352_/S _12411_/C vssd1 vssd1 vccd1
+ vccd1 _12413_/X sky130_fd_sc_hd__mux4_1
XFILLER_201_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16181_ _17432_/A _16181_/B vssd1 vssd1 vccd1 vccd1 _19614_/D sky130_fd_sc_hd__and2_1
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13393_ _13002_/A _13253_/C _13389_/X _13392_/X vssd1 vssd1 vccd1 vccd1 _13393_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_194_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15132_ _21014_/Q _20982_/Q _15508_/S vssd1 vssd1 vccd1 vccd1 _15132_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12344_ _19693_/Q _20181_/Q _12344_/S vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19940_ _20669_/CLK _19940_/D vssd1 vssd1 vccd1 vccd1 _19940_/Q sky130_fd_sc_hd__dfxtp_1
X_15063_ _15061_/X _15062_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _15063_/X sky130_fd_sc_hd__mux2_1
X_12275_ _12275_/A _12275_/B _12274_/X vssd1 vssd1 vccd1 vccd1 _12275_/X sky130_fd_sc_hd__or3b_4
XFILLER_181_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14014_ _14041_/A1 _09672_/B _09786_/X _14041_/B1 _19853_/Q vssd1 vssd1 vccd1 vccd1
+ _14089_/C sky130_fd_sc_hd__o32a_1
X_11226_ _09643_/A _09686_/D _11225_/Y _09586_/Y vssd1 vssd1 vccd1 vccd1 _11226_/X
+ sky130_fd_sc_hd__o211a_1
X_19871_ _20084_/CLK _19871_/D vssd1 vssd1 vccd1 vccd1 _19871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18822_ _19093_/Q _12589_/B _12592_/C _13596_/X vssd1 vssd1 vccd1 vccd1 _18823_/B
+ sky130_fd_sc_hd__a22o_1
X_11157_ _13192_/A _19268_/Q _20055_/Q _12295_/B _11363_/A1 vssd1 vssd1 vccd1 vccd1
+ _11157_/X sky130_fd_sc_hd__o221a_1
XFILLER_150_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10108_ _10087_/X _10095_/X _10101_/X _10107_/X vssd1 vssd1 vccd1 vccd1 _10108_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_249_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18753_ _20977_/Q _18315_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18754_/B sky130_fd_sc_hd__mux2_1
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11088_ _12399_/A1 _11087_/X _11084_/X _12392_/C1 vssd1 vssd1 vccd1 vccd1 _11088_/X
+ sky130_fd_sc_hd__o211a_2
X_15965_ _21040_/Q _21008_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _15965_/X sky130_fd_sc_hd__mux2_1
Xinput260 manufacturerID[6] vssd1 vssd1 vccd1 vccd1 _17257_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput271 partID[1] vssd1 vssd1 vccd1 vccd1 _17275_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_248_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17704_ _20488_/Q _17704_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20488_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput282 versionID[2] vssd1 vssd1 vccd1 vccd1 _15133_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10039_ _09672_/A _14041_/A2 _10038_/X _11228_/B1 _19859_/Q vssd1 vssd1 vccd1 vccd1
+ _10039_/X sky130_fd_sc_hd__o32a_1
X_14916_ _14917_/A _12513_/B _14915_/X vssd1 vssd1 vccd1 vccd1 _14981_/A sky130_fd_sc_hd__a21o_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18684_ _18556_/X _18684_/A2 _18682_/Y _18683_/Y vssd1 vssd1 vccd1 vccd1 _18685_/B
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_196_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20574_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_252_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15896_ _12513_/B _15978_/A2 _15980_/A2 vssd1 vssd1 vccd1 vccd1 _15896_/X sky130_fd_sc_hd__a21bo_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17635_ _20391_/Q _17946_/A1 _17635_/S vssd1 vssd1 vccd1 vccd1 _20391_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_125_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20624_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14847_ _14845_/X _14846_/X _15058_/S vssd1 vssd1 vccd1 vccd1 _14847_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17566_ _20326_/Q _17805_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20326_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14778_ _19136_/Q _14798_/A2 _14777_/X _14794_/C1 vssd1 vssd1 vccd1 vccd1 _19513_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_251_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19305_ _20660_/CLK _19305_/D vssd1 vssd1 vccd1 vccd1 _19305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16517_ _19824_/Q _17178_/A1 _16517_/S vssd1 vssd1 vccd1 vccd1 _19824_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13729_ _13780_/A _13729_/B vssd1 vssd1 vccd1 vccd1 _13729_/X sky130_fd_sc_hd__and2_1
X_17497_ _17505_/A1 _17496_/Y _18104_/A vssd1 vssd1 vccd1 vccd1 _20283_/D sky130_fd_sc_hd__a21oi_1
XFILLER_220_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19236_ _19520_/CLK _19236_/D vssd1 vssd1 vccd1 vccd1 _19236_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_177_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16448_ _19763_/Q _16450_/C _16447_/Y vssd1 vssd1 vccd1 vccd1 _19763_/D sky130_fd_sc_hd__o21a_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19167_ _20426_/CLK _19167_/D vssd1 vssd1 vccd1 vccd1 _19167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16379_ _18054_/A _16379_/B _16380_/B vssd1 vssd1 vccd1 vccd1 _19737_/D sky130_fd_sc_hd__nor3_1
XFILLER_158_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18118_ _18905_/A _18118_/B _18122_/C vssd1 vssd1 vccd1 vccd1 _20781_/D sky130_fd_sc_hd__nor3_1
XFILLER_191_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19098_ _20721_/CLK _19098_/D vssd1 vssd1 vccd1 vccd1 _19098_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18049_ _20755_/Q _18047_/B _18048_/Y vssd1 vssd1 vccd1 vccd1 _20755_/D sky130_fd_sc_hd__o21a_1
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20011_ _20014_/CLK _20011_/D vssd1 vssd1 vccd1 vccd1 _20011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _12072_/A1 _09821_/X _09818_/X _12072_/C1 vssd1 vssd1 vccd1 vccd1 _09822_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09753_ _19821_/Q _12009_/A2 _09751_/X _11563_/S _09752_/X vssd1 vssd1 vccd1 vccd1
+ _09753_/X sky130_fd_sc_hd__o221a_1
XFILLER_227_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09684_ _09684_/A _11326_/A vssd1 vssd1 vccd1 vccd1 _09684_/X sky130_fd_sc_hd__and2_1
XFILLER_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20913_ _20913_/CLK _20913_/D vssd1 vssd1 vccd1 vccd1 _20913_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ _21006_/CLK _20844_/D vssd1 vssd1 vccd1 vccd1 _20844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20775_ _21029_/CLK _20775_/D vssd1 vssd1 vccd1 vccd1 _20775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10390_ _10387_/X _10388_/X _10389_/X _09507_/A _10516_/S vssd1 vssd1 vccd1 vccd1
+ _10390_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12060_ _12060_/A1 _20519_/Q _10585_/S _12042_/X vssd1 vssd1 vccd1 vccd1 _12060_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11011_ _09689_/C _10999_/X _11002_/X _11010_/X vssd1 vssd1 vccd1 vccd1 _11012_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_145_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1904 fanout1905/X vssd1 vssd1 vccd1 vccd1 _14482_/A sky130_fd_sc_hd__buf_2
XFILLER_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20209_ _20766_/CLK _20209_/D vssd1 vssd1 vccd1 vccd1 _20209_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1915 _18726_/A vssd1 vssd1 vccd1 vccd1 _18352_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1926 _16193_/A vssd1 vssd1 vccd1 vccd1 _16197_/A sky130_fd_sc_hd__buf_4
XFILLER_77_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1937 _14185_/C1 vssd1 vssd1 vccd1 vccd1 _18396_/A sky130_fd_sc_hd__buf_2
Xfanout1948 fanout1960/X vssd1 vssd1 vccd1 vccd1 _14104_/C1 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout950 _10933_/Y vssd1 vssd1 vccd1 vccd1 _15610_/A1 sky130_fd_sc_hd__buf_12
Xfanout1959 fanout1960/X vssd1 vssd1 vccd1 vccd1 _18416_/A sky130_fd_sc_hd__buf_4
Xfanout961 _11331_/X vssd1 vssd1 vccd1 vccd1 _11397_/A2 sky130_fd_sc_hd__buf_6
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout972 split4/A vssd1 vssd1 vccd1 vccd1 _17095_/A1 sky130_fd_sc_hd__buf_4
XFILLER_93_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout983 _17199_/A1 vssd1 vssd1 vccd1 vccd1 _17933_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout994 _16719_/X vssd1 vssd1 vccd1 vccd1 _17005_/A2 sky130_fd_sc_hd__buf_4
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _12960_/X _12961_/X _12962_/S vssd1 vssd1 vccd1 vccd1 _12963_/D sky130_fd_sc_hd__mux2_4
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _16017_/C1 _15749_/X _15745_/X vssd1 vssd1 vccd1 vccd1 _15750_/X sky130_fd_sc_hd__o21a_2
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _19460_/Q _17707_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19460_/D sky130_fd_sc_hd__mux2_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _19823_/Q _19327_/Q _11915_/S vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12893_ _12911_/A _12893_/B vssd1 vssd1 vccd1 vccd1 _12894_/B sky130_fd_sc_hd__or2_1
XANTENNA_310 input238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15681_ _11752_/X _15981_/B _15680_/X vssd1 vssd1 vccd1 vccd1 _15681_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 _13494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_332 _20261_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17420_ _17420_/A _17432_/A vssd1 vssd1 vccd1 vccd1 _20256_/D sky130_fd_sc_hd__and2_1
XFILLER_61_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _19396_/Q _17916_/A1 _14632_/S vssd1 vssd1 vccd1 vccd1 _19396_/D sky130_fd_sc_hd__mux2_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_343 _19502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ _09501_/Y _16063_/B2 _11843_/X vssd1 vssd1 vccd1 vccd1 _11877_/A sky130_fd_sc_hd__a21oi_2
XFILLER_260_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_354 _17905_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_365 _11367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_376 _12504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _19333_/Q _17674_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19333_/D sky130_fd_sc_hd__mux2_1
X_17351_ _20224_/Q _17363_/A2 _17350_/X _18692_/A vssd1 vssd1 vccd1 vccd1 _20224_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_387 _16815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_398 _16018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11775_ _13541_/A _11775_/B vssd1 vssd1 vccd1 vccd1 _11787_/A sky130_fd_sc_hd__xnor2_1
XFILLER_199_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16306_/C _16302_/B vssd1 vssd1 vccd1 vccd1 _19708_/D sky130_fd_sc_hd__nor2_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _11061_/A _16081_/A vssd1 vssd1 vccd1 vccd1 _10726_/Y sky130_fd_sc_hd__nor2_1
X_13514_ _19219_/Q _13499_/A _14110_/B vssd1 vssd1 vccd1 vccd1 _13514_/Y sky130_fd_sc_hd__a21oi_1
X_17282_ _20199_/Q _17330_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17282_/X sky130_fd_sc_hd__a21o_1
X_14494_ _19272_/Q _17751_/A1 _14519_/S vssd1 vssd1 vccd1 vccd1 _19272_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19021_ _21029_/Q _19015_/B _19020_/X _18728_/A vssd1 vssd1 vccd1 vccd1 _21029_/D
+ sky130_fd_sc_hd__o211a_1
X_16233_ _13441_/X _16233_/B vssd1 vssd1 vccd1 vccd1 _16233_/X sky130_fd_sc_hd__and2b_1
X_13445_ split3/X _13463_/C _19695_/Q vssd1 vssd1 vccd1 vccd1 _13446_/B sky130_fd_sc_hd__a21oi_4
X_10657_ _20532_/Q _12323_/S vssd1 vssd1 vccd1 vccd1 _10657_/X sky130_fd_sc_hd__or2_1
XFILLER_277_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16164_ _16869_/B _16164_/B vssd1 vssd1 vccd1 vccd1 _16164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13376_ _13377_/A _13377_/B vssd1 vssd1 vccd1 vccd1 _13376_/X sky130_fd_sc_hd__and2_1
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10588_ _19807_/Q _19311_/Q _11682_/S vssd1 vssd1 vccd1 vccd1 _10588_/X sky130_fd_sc_hd__mux2_1
X_12327_ _12402_/A1 _17951_/A1 _12401_/B1 vssd1 vssd1 vccd1 vccd1 _12327_/X sky130_fd_sc_hd__o21a_1
X_15115_ _15167_/S _14872_/A _15254_/S vssd1 vssd1 vccd1 vccd1 _15115_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16095_ _19572_/Q _16079_/B _16107_/B1 vssd1 vssd1 vccd1 vccd1 _16095_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15046_ _14843_/X _14852_/X _15058_/S vssd1 vssd1 vccd1 vccd1 _15046_/X sky130_fd_sc_hd__mux2_1
X_19923_ _20669_/CLK _19923_/D vssd1 vssd1 vccd1 vccd1 _19923_/Q sky130_fd_sc_hd__dfxtp_1
X_12258_ _12252_/X _12257_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _12258_/X sky130_fd_sc_hd__mux2_2
XFILLER_170_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11209_ _12430_/S _11204_/X _11208_/Y _11384_/S vssd1 vssd1 vccd1 vccd1 _11209_/X
+ sky130_fd_sc_hd__o211a_1
X_19854_ _20017_/CLK _19854_/D vssd1 vssd1 vccd1 vccd1 _19854_/Q sky130_fd_sc_hd__dfxtp_4
X_12189_ _12189_/A _12189_/B vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__or2_1
XFILLER_284_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18805_ _18589_/Y _18818_/A2 _18803_/Y _18804_/Y vssd1 vssd1 vccd1 vccd1 _18805_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19785_ _20081_/CLK _19785_/D vssd1 vssd1 vccd1 vccd1 _19785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16997_ _17006_/A1 _16021_/X _16945_/X _16996_/X vssd1 vssd1 vccd1 vccd1 _16997_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18736_ _18736_/A _18736_/B vssd1 vssd1 vccd1 vccd1 _20968_/D sky130_fd_sc_hd__and2_1
XFILLER_95_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ _15948_/A1 _12880_/X _15947_/X _12832_/B vssd1 vssd1 vccd1 vccd1 _15948_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_236_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18667_ _19520_/Q _18667_/B vssd1 vssd1 vccd1 vccd1 _18667_/Y sky130_fd_sc_hd__nand2_1
X_15879_ _16017_/C1 _15878_/X _15874_/X vssd1 vssd1 vccd1 vccd1 _15879_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17618_ _20374_/Q _17686_/A1 _17635_/S vssd1 vssd1 vccd1 vccd1 _20374_/D sky130_fd_sc_hd__mux2_1
XFILLER_212_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18598_ _18598_/A _18598_/B vssd1 vssd1 vccd1 vccd1 _20922_/D sky130_fd_sc_hd__nor2_1
XFILLER_212_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17549_ _20309_/Q _17928_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20309_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20560_ _20565_/CLK _20560_/D vssd1 vssd1 vccd1 vccd1 _20560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19219_ _19219_/CLK _19219_/D vssd1 vssd1 vccd1 vccd1 _19219_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_93_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20663_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20491_ _20491_/CLK _20491_/D vssd1 vssd1 vccd1 vccd1 _20491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_wb_clk_i _20408_/CLK vssd1 vssd1 vccd1 vccd1 _20666_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_192_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21043_ _21043_/CLK _21043_/D vssd1 vssd1 vccd1 vccd1 _21043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09805_ _09796_/X _09798_/X _09804_/X _12058_/S _12136_/B1 vssd1 vssd1 vccd1 vccd1
+ _09805_/X sky130_fd_sc_hd__o221a_1
XFILLER_189_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09736_ _10937_/A _14112_/B vssd1 vssd1 vccd1 vccd1 _09736_/Y sky130_fd_sc_hd__nor2_8
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09667_ _11242_/A1 _13978_/A2 _09664_/C _09665_/X _11243_/S vssd1 vssd1 vccd1 vccd1
+ _09680_/C sky130_fd_sc_hd__o311ai_4
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09598_ _09609_/A _19092_/Q vssd1 vssd1 vccd1 vccd1 _16454_/B sky130_fd_sc_hd__nand2b_4
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20827_ _21021_/CLK _20827_/D vssd1 vssd1 vccd1 vccd1 _20827_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11560_ _12190_/C1 _11557_/X _11559_/X vssd1 vssd1 vccd1 vccd1 _11560_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20758_ _20759_/CLK _20758_/D vssd1 vssd1 vccd1 vccd1 _20758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ _10356_/A _19344_/Q _20699_/Q _10518_/S _11304_/S vssd1 vssd1 vccd1 vccd1
+ _10511_/X sky130_fd_sc_hd__a221o_1
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ _12012_/S _11482_/X _11490_/X _11474_/X vssd1 vssd1 vccd1 vccd1 _11491_/X
+ sky130_fd_sc_hd__a31o_1
X_20689_ _20704_/CLK _20689_/D vssd1 vssd1 vccd1 vccd1 _20689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13230_ _13139_/A _19241_/Q _13229_/X vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__a21o_2
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10442_ _19634_/Q _10502_/A2 _10439_/X _10440_/X _10441_/X vssd1 vssd1 vccd1 vccd1
+ _10442_/X sky130_fd_sc_hd__o221a_1
X_13161_ _11415_/A _13422_/B _11575_/B _10276_/Y vssd1 vssd1 vccd1 vccd1 _13162_/B
+ sky130_fd_sc_hd__a211o_2
X_10373_ _10373_/A _11234_/B _10372_/X vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__or3b_1
XFILLER_151_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12112_ _12112_/A _13431_/A _13432_/A vssd1 vssd1 vccd1 vccd1 _12112_/X sky130_fd_sc_hd__or3b_1
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13092_ _20976_/Q _20910_/Q _13091_/X vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16920_ _19981_/Q _16876_/A _16919_/Y _18704_/A vssd1 vssd1 vccd1 vccd1 _19981_/D
+ sky130_fd_sc_hd__a211o_1
X_12043_ _19955_/Q _12043_/B vssd1 vssd1 vccd1 vccd1 _12043_/X sky130_fd_sc_hd__or2_1
Xfanout1701 _12254_/A vssd1 vssd1 vccd1 vccd1 _11391_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_46_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1712 _12270_/B1 vssd1 vssd1 vccd1 vccd1 _12347_/C1 sky130_fd_sc_hd__buf_4
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1723 _10581_/A1 vssd1 vssd1 vccd1 vccd1 _12060_/A1 sky130_fd_sc_hd__buf_6
XFILLER_120_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1734 _09504_/Y vssd1 vssd1 vccd1 vccd1 _12312_/A1 sky130_fd_sc_hd__buf_6
X_16851_ _16869_/A _16851_/B vssd1 vssd1 vccd1 vccd1 _16851_/Y sky130_fd_sc_hd__nand2_1
Xfanout1745 _09502_/Y vssd1 vssd1 vccd1 vccd1 _12059_/A1 sky130_fd_sc_hd__buf_8
XFILLER_265_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1756 _13967_/S vssd1 vssd1 vccd1 vccd1 _14042_/S sky130_fd_sc_hd__buf_6
XFILLER_266_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1767 _13275_/A1 vssd1 vssd1 vccd1 vccd1 _09488_/A sky130_fd_sc_hd__buf_6
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout780 _14110_/A vssd1 vssd1 vccd1 vccd1 _18589_/B sky130_fd_sc_hd__buf_4
Xfanout1778 _20263_/Q vssd1 vssd1 vccd1 vccd1 _17441_/A sky130_fd_sc_hd__buf_4
X_15802_ _20936_/Q _16044_/A2 _15801_/X vssd1 vssd1 vccd1 vccd1 _15802_/X sky130_fd_sc_hd__o21a_1
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout791 _12744_/B vssd1 vssd1 vccd1 vccd1 _12857_/B sky130_fd_sc_hd__clkbuf_4
X_19570_ _20341_/CLK _19570_/D vssd1 vssd1 vccd1 vccd1 _19570_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1789 _18163_/A vssd1 vssd1 vccd1 vccd1 _18134_/A sky130_fd_sc_hd__buf_6
XFILLER_219_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16782_ _16778_/Y _16781_/X _17011_/B1 vssd1 vssd1 vccd1 vccd1 _16782_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_77_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13994_ _19197_/Q _14075_/C _14042_/S vssd1 vssd1 vccd1 vccd1 _13994_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18521_ _20900_/Q _18559_/B _18520_/X _18458_/B vssd1 vssd1 vccd1 vccd1 _18522_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_219_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _19546_/Q _16036_/A2 _15732_/X _16185_/A vssd1 vssd1 vccd1 vccd1 _19546_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12945_ _12945_/A _14921_/B _12945_/C vssd1 vssd1 vccd1 vccd1 _16720_/C sky130_fd_sc_hd__or3_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _18740_/A _18452_/B vssd1 vssd1 vccd1 vccd1 _20880_/D sky130_fd_sc_hd__and2_1
XFILLER_283_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _21029_/Q _20997_/Q _15993_/S vssd1 vssd1 vccd1 vccd1 _15664_/X sky130_fd_sc_hd__mux2_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12876_ _12911_/A _12877_/B vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__and2_1
XANTENNA_140 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 _13760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 _13839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17403_ _17402_/A _17441_/A _17457_/B _20250_/Q vssd1 vssd1 vccd1 vccd1 _17403_/X
+ sky130_fd_sc_hd__a31o_1
X_14615_ _19379_/Q _17899_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19379_/D sky130_fd_sc_hd__mux2_1
XANTENNA_173 _19111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11827_ _12752_/A _20517_/Q _12143_/S _11809_/X vssd1 vssd1 vccd1 vccd1 _11827_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_184 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18383_ _18553_/B _18387_/B vssd1 vssd1 vccd1 vccd1 _18383_/Y sky130_fd_sc_hd__nand2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _19717_/Q _15595_/A2 _15595_/B1 _19749_/Q vssd1 vssd1 vccd1 vccd1 _15595_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _19542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17333_/X _17334_/B vssd1 vssd1 vccd1 vccd1 _20217_/D sky130_fd_sc_hd__and2b_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _19316_/Q _17934_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19316_/D sky130_fd_sc_hd__mux2_1
X_11758_ _13415_/A _11758_/B _15734_/A vssd1 vssd1 vccd1 vccd1 _15763_/A sky130_fd_sc_hd__nand3_1
XFILLER_53_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ _12427_/A1 _19341_/Q _20696_/Q _12417_/S _12419_/C1 vssd1 vssd1 vccd1 vccd1
+ _10709_/X sky130_fd_sc_hd__a221o_1
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17265_ _20194_/Q _17268_/A2 _17263_/X _17264_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1
+ _20194_/D sky130_fd_sc_hd__o221a_1
X_14477_ _20234_/Q _19263_/Q _14477_/S vssd1 vssd1 vccd1 vccd1 _14478_/B sky130_fd_sc_hd__mux2_1
X_11689_ _10561_/A _11687_/X _11688_/X vssd1 vssd1 vccd1 vccd1 _11689_/X sky130_fd_sc_hd__a21o_1
X_19004_ _18205_/Y _18982_/B _19016_/B1 _19003_/X vssd1 vssd1 vccd1 vccd1 _21021_/D
+ sky130_fd_sc_hd__o211a_1
X_16216_ _19639_/Q _17202_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19639_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13428_ _15762_/A _13428_/B _13428_/C _13428_/D vssd1 vssd1 vccd1 vccd1 _13429_/B
+ sky130_fd_sc_hd__or4_1
X_17196_ _20160_/Q _17687_/A1 _17215_/S vssd1 vssd1 vccd1 vccd1 _20160_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16147_ _19597_/Q _16194_/S _16146_/Y _16195_/A vssd1 vssd1 vccd1 vccd1 _19597_/D
+ sky130_fd_sc_hd__o211a_1
X_13359_ _13359_/A vssd1 vssd1 vccd1 vccd1 _13359_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16078_ _19563_/Q _16077_/B _16077_/Y _16097_/B1 vssd1 vssd1 vccd1 vccd1 _19563_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15029_ _15442_/A _13658_/A _15023_/Y _15028_/Y vssd1 vssd1 vccd1 vccd1 _15029_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19906_ _20438_/CLK _19906_/D vssd1 vssd1 vccd1 vccd1 _19906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_269_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19837_ _20751_/CLK _19837_/D vssd1 vssd1 vccd1 vccd1 _19837_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_57_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_140_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19697_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 coreIndex[1] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_6
X_19768_ _20720_/CLK _19768_/D vssd1 vssd1 vccd1 vccd1 _19768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09521_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09521_/Y sky130_fd_sc_hd__inv_2
XFILLER_272_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18719_ _20960_/Q _18230_/Y _18719_/S vssd1 vssd1 vccd1 vccd1 _18720_/B sky130_fd_sc_hd__mux2_1
XFILLER_271_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19699_ _19701_/CLK _19699_/D vssd1 vssd1 vccd1 vccd1 _19699_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20612_ _20717_/CLK _20612_/D vssd1 vssd1 vccd1 vccd1 _20612_/Q sky130_fd_sc_hd__dfxtp_1
X_20543_ _20675_/CLK _20543_/D vssd1 vssd1 vccd1 vccd1 _20543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20474_ _20692_/CLK _20474_/D vssd1 vssd1 vccd1 vccd1 _20474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput350 _13745_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[24] sky130_fd_sc_hd__buf_4
XFILLER_133_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput361 _13656_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[5] sky130_fd_sc_hd__buf_4
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput372 _13476_/X vssd1 vssd1 vccd1 vccd1 csb0[0] sky130_fd_sc_hd__buf_4
Xoutput383 _13807_/X vssd1 vssd1 vccd1 vccd1 din0[16] sky130_fd_sc_hd__buf_4
XFILLER_120_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput394 _13817_/X vssd1 vssd1 vccd1 vccd1 din0[26] sky130_fd_sc_hd__buf_4
Xfanout1008 _15982_/C vssd1 vssd1 vccd1 vccd1 _15925_/B sky130_fd_sc_hd__buf_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1019 _18785_/A2 vssd1 vssd1 vccd1 vccd1 _12589_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_248_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21026_ _21026_/CLK _21026_/D vssd1 vssd1 vccd1 vccd1 _21026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09719_ _20045_/Q _19920_/Q _11889_/S vssd1 vssd1 vccd1 vccd1 _09719_/X sky130_fd_sc_hd__mux2_1
XFILLER_274_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10991_ _19665_/Q _10217_/S _10990_/X _11338_/A1 vssd1 vssd1 vccd1 vccd1 _10991_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_216_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12479_/A _12730_/A2 _12731_/B _12729_/X vssd1 vssd1 vccd1 vccd1 _12730_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12661_ _12662_/B _12662_/C _12662_/A vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__a21oi_2
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14400_ _19522_/Q _14406_/B vssd1 vssd1 vccd1 vccd1 _14400_/Y sky130_fd_sc_hd__nor2_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11612_ _12156_/A1 _11610_/X _11611_/X vssd1 vssd1 vccd1 vccd1 _11612_/X sky130_fd_sc_hd__a21o_1
XFILLER_168_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12592_/A _12592_/B _12592_/C _12557_/Y vssd1 vssd1 vccd1 vccd1 _12592_/X
+ sky130_fd_sc_hd__or4b_4
X_15380_ _15380_/A _16009_/B vssd1 vssd1 vccd1 vccd1 _15380_/Y sky130_fd_sc_hd__nand2_1
XFILLER_212_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14331_ _19515_/Q _14332_/B vssd1 vssd1 vccd1 vccd1 _14343_/A sky130_fd_sc_hd__nand2_1
X_11543_ _09986_/A _20134_/Q _20102_/Q _09928_/S vssd1 vssd1 vccd1 vccd1 _11543_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17050_ _20022_/Q _17852_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20022_/D sky130_fd_sc_hd__mux2_1
X_14262_ _14262_/A _14262_/B _14271_/B vssd1 vssd1 vccd1 vccd1 _14262_/X sky130_fd_sc_hd__or3b_1
X_11474_ _12192_/A1 _11469_/X _11473_/X _10409_/A _11466_/X vssd1 vssd1 vccd1 vccd1
+ _11474_/X sky130_fd_sc_hd__o311a_1
XFILLER_183_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13213_ _20941_/Q _13366_/C1 _13212_/X _18687_/B vssd1 vssd1 vccd1 vccd1 _13213_/X
+ sky130_fd_sc_hd__a211o_1
X_16001_ _16050_/A1 _16000_/X _15988_/Y vssd1 vssd1 vccd1 vccd1 _16001_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_109_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _20472_/Q _20312_/Q _10425_/S vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14193_ _13582_/A _14192_/X _13565_/X vssd1 vssd1 vccd1 vccd1 _14194_/C sky130_fd_sc_hd__a21bo_1
X_13144_ _15075_/A _15061_/S _11783_/B _15071_/S _11140_/A vssd1 vssd1 vccd1 vccd1
+ _13145_/B sky130_fd_sc_hd__a311o_2
X_10356_ _10356_/A _19316_/Q _11290_/C vssd1 vssd1 vccd1 vccd1 _10356_/X sky130_fd_sc_hd__or3_1
XFILLER_3_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_11__f_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_74_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17952_ _17952_/A _17952_/B vssd1 vssd1 vccd1 vccd1 _20721_/D sky130_fd_sc_hd__nor2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13075_ _13031_/Y _13354_/A _13353_/B vssd1 vssd1 vccd1 vccd1 _13340_/A sky130_fd_sc_hd__o21ai_2
XFILLER_250_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10287_ input130/X input165/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10287_/X sky130_fd_sc_hd__mux2_8
XFILLER_3_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16903_ _16900_/Y _16902_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16903_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1520 _11987_/S vssd1 vssd1 vccd1 vccd1 _12124_/S sky130_fd_sc_hd__buf_6
X_12026_ _12103_/A1 _12025_/X _12024_/X vssd1 vssd1 vccd1 vccd1 _12026_/X sky130_fd_sc_hd__o21a_1
Xfanout1531 fanout1534/X vssd1 vssd1 vccd1 vccd1 _10425_/S sky130_fd_sc_hd__buf_4
X_17883_ _20656_/Q _17917_/A1 _17883_/S vssd1 vssd1 vccd1 vccd1 _20656_/D sky130_fd_sc_hd__mux2_1
XFILLER_266_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1542 _10137_/C vssd1 vssd1 vccd1 vccd1 _10983_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_211_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1553 _11090_/S vssd1 vssd1 vccd1 vccd1 _12397_/S sky130_fd_sc_hd__buf_6
XFILLER_254_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1564 _10842_/S vssd1 vssd1 vccd1 vccd1 _11161_/S sky130_fd_sc_hd__clkbuf_8
X_19622_ _20410_/CLK _19622_/D vssd1 vssd1 vccd1 vccd1 _19622_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1575 _12151_/A1 vssd1 vssd1 vccd1 vccd1 _12140_/C1 sky130_fd_sc_hd__buf_6
X_16834_ _20408_/Q _17004_/A2 _17004_/B1 vssd1 vssd1 vccd1 vccd1 _16834_/X sky130_fd_sc_hd__a21o_1
Xfanout1586 _12144_/A1 vssd1 vssd1 vccd1 vccd1 _12147_/C1 sky130_fd_sc_hd__buf_8
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1597 _11528_/S vssd1 vssd1 vccd1 vccd1 _11917_/S sky130_fd_sc_hd__buf_6
XFILLER_65_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19553_ _19617_/CLK _19553_/D vssd1 vssd1 vccd1 vccd1 _19553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16765_ _19088_/Q _16996_/B1 _16764_/X vssd1 vssd1 vccd1 vccd1 _16765_/X sky130_fd_sc_hd__o21a_1
XFILLER_65_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13977_ _19159_/Q _14004_/A2 _14004_/B1 _13976_/X _16087_/B1 vssd1 vssd1 vccd1 vccd1
+ _19159_/D sky130_fd_sc_hd__o221a_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18504_ _18856_/A _18504_/B vssd1 vssd1 vccd1 vccd1 _20894_/D sky130_fd_sc_hd__nor2_1
X_15716_ _20741_/Q _15934_/A2 _15934_/B1 _20773_/Q vssd1 vssd1 vccd1 vccd1 _15716_/X
+ sky130_fd_sc_hd__a22o_1
X_12928_ _12928_/A _12928_/B _12928_/C _13466_/A vssd1 vssd1 vccd1 vccd1 _14117_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19484_ _20451_/CLK _19484_/D vssd1 vssd1 vccd1 vccd1 _19484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16696_ _19951_/Q _17874_/A1 _16701_/S vssd1 vssd1 vccd1 vccd1 _19951_/D sky130_fd_sc_hd__mux2_1
XFILLER_207_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18435_ _20872_/Q _18270_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18436_/B sky130_fd_sc_hd__mux2_1
X_15647_ _15890_/B _15629_/Y _15646_/X _15976_/B2 vssd1 vssd1 vccd1 vccd1 _15647_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12859_ _15703_/B2 _12856_/X _12857_/X _12860_/A vssd1 vssd1 vccd1 vccd1 _13332_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18366_ _20838_/Q _18375_/B _18365_/Y _18748_/A vssd1 vssd1 vccd1 vccd1 _20838_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_221_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15578_ _15069_/X _15577_/X _15578_/S vssd1 vssd1 vccd1 vccd1 _15578_/X sky130_fd_sc_hd__mux2_4
XFILLER_159_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17317_ input4/X input270/X _17320_/S vssd1 vssd1 vccd1 vccd1 _17317_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14529_ _19094_/Q _19093_/Q _14668_/B vssd1 vssd1 vccd1 vccd1 _16672_/A sky130_fd_sc_hd__or3_2
X_18297_ _18730_/A _18297_/B vssd1 vssd1 vccd1 vccd1 _20813_/D sky130_fd_sc_hd__and2_1
XFILLER_179_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17248_ _17248_/A _17275_/B _17269_/C vssd1 vssd1 vccd1 vccd1 _17248_/X sky130_fd_sc_hd__and3_1
XFILLER_190_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17179_ _20145_/Q _17704_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20145_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20190_ _20428_/CLK _20190_/D vssd1 vssd1 vccd1 vccd1 _20190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _13192_/A vssd1 vssd1 vccd1 vccd1 _09504_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_65_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_40 _16750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_51 _16935_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_62 _18195_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20526_ _20659_/CLK _20526_/D vssd1 vssd1 vccd1 vccd1 _20526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_73 _09607_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 _11132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_95 _15988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20457_ _20645_/CLK _20457_/D vssd1 vssd1 vccd1 vccd1 _20457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_273_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10210_ _10208_/X _10209_/X _10235_/S vssd1 vssd1 vccd1 vccd1 _10210_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ _11391_/A _19898_/Q _11393_/S0 _20023_/Q vssd1 vssd1 vccd1 vccd1 _11190_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_284_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20388_ _20712_/CLK _20388_/D vssd1 vssd1 vccd1 vccd1 _20388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ _10131_/X _10132_/X _12376_/S vssd1 vssd1 vccd1 vccd1 _10141_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10072_ _19810_/Q _10502_/A2 _10070_/X _11684_/A1 _10071_/X vssd1 vssd1 vccd1 vccd1
+ _10072_/X sky130_fd_sc_hd__o221a_1
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13900_ _18048_/A _13900_/A2 _14522_/A _14112_/A vssd1 vssd1 vccd1 vccd1 _19116_/D
+ sky130_fd_sc_hd__o22a_1
X_21009_ _21009_/CLK _21009_/D vssd1 vssd1 vccd1 vccd1 _21009_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14880_ _14881_/A _14881_/B vssd1 vssd1 vccd1 vccd1 _14880_/Y sky130_fd_sc_hd__nor2_1
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13831_ _20001_/Q _13473_/X _13785_/X split2/X vssd1 vssd1 vccd1 vccd1 _13831_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16550_ _19841_/Q _16578_/A2 _16578_/B1 input11/X vssd1 vssd1 vccd1 vccd1 _16551_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_262_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10974_ input140/X input135/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10974_/X sky130_fd_sc_hd__mux2_8
XFILLER_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13762_ _13777_/A _13762_/B vssd1 vssd1 vccd1 vccd1 _13762_/X sky130_fd_sc_hd__or2_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _14878_/B _15500_/X _10113_/A vssd1 vssd1 vccd1 vccd1 _15501_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_189_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12713_ _12709_/X _12711_/Y _12706_/Y _12707_/X vssd1 vssd1 vccd1 vccd1 _12726_/B
+ sky130_fd_sc_hd__a211oi_2
X_16481_ _19790_/Q _17804_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19790_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ _13693_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13693_/X sky130_fd_sc_hd__or2_2
XFILLER_280_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18220_ _18502_/B vssd1 vssd1 vccd1 vccd1 _18220_/Y sky130_fd_sc_hd__inv_4
X_15432_ _19536_/Q _15492_/A _15431_/Y _16179_/A vssd1 vssd1 vccd1 vccd1 _19536_/D
+ sky130_fd_sc_hd__o211a_1
X_12644_ _12642_/Y _12643_/X _12513_/A _13589_/A1 vssd1 vssd1 vccd1 vccd1 _12698_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_203_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18151_ _18318_/B _18318_/C vssd1 vssd1 vccd1 vccd1 _18157_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15363_ _15612_/S _15362_/Y _15610_/B1 vssd1 vssd1 vccd1 vccd1 _15363_/X sky130_fd_sc_hd__a21bo_1
X_12575_ _12577_/B vssd1 vssd1 vccd1 vccd1 _12575_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17102_ _20072_/Q _17695_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20072_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14314_ _14314_/A _14314_/B vssd1 vssd1 vccd1 vccd1 _14323_/B sky130_fd_sc_hd__or2_1
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18082_ _20768_/Q _18085_/C _18086_/A vssd1 vssd1 vccd1 vccd1 _18082_/Y sky130_fd_sc_hd__a21oi_1
X_11526_ _20038_/Q _19913_/Q _11916_/S vssd1 vssd1 vccd1 vccd1 _11526_/X sky130_fd_sc_hd__mux2_1
X_15294_ _15290_/X _15293_/X _15578_/S vssd1 vssd1 vccd1 vccd1 _15294_/X sky130_fd_sc_hd__mux2_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17033_ _20011_/Q input197/X _17040_/S vssd1 vssd1 vccd1 vccd1 _20011_/D sky130_fd_sc_hd__mux2_1
X_11457_ _12850_/A1 _11649_/S _11456_/Y vssd1 vssd1 vccd1 vccd1 _11495_/A sky130_fd_sc_hd__o21a_1
X_14245_ _14255_/A _16068_/B _14245_/C vssd1 vssd1 vccd1 vccd1 _14245_/X sky130_fd_sc_hd__or3_1
XFILLER_194_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10408_ _10406_/X _10407_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _10409_/B sky130_fd_sc_hd__mux2_1
X_14176_ _19500_/Q _14177_/B vssd1 vssd1 vccd1 vccd1 _14176_/Y sky130_fd_sc_hd__nor2_2
X_11388_ _19631_/Q _19937_/Q _19275_/Q _20062_/Q _12344_/S _11391_/C vssd1 vssd1 vccd1
+ vccd1 _11388_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10339_ _10336_/X _10338_/X _12514_/C vssd1 vssd1 vccd1 vccd1 _10339_/X sky130_fd_sc_hd__a21o_1
X_13127_ _19243_/Q _13114_/B _19244_/Q vssd1 vssd1 vccd1 vccd1 _13127_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18984_ _21012_/Q _18997_/B vssd1 vssd1 vccd1 vccd1 _18984_/X sky130_fd_sc_hd__or2_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _20704_/Q _17935_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20704_/D sky130_fd_sc_hd__mux2_1
X_13058_ _20949_/Q _20883_/Q vssd1 vssd1 vccd1 vccd1 _13060_/C sky130_fd_sc_hd__nand2_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1350 _17038_/S vssd1 vssd1 vccd1 vccd1 _17849_/S sky130_fd_sc_hd__buf_6
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12009_ _19393_/Q _12009_/A2 _12007_/X _12190_/C1 _12008_/X vssd1 vssd1 vccd1 vccd1
+ _12009_/X sky130_fd_sc_hd__o221a_1
Xfanout1361 _14002_/B1 vssd1 vssd1 vccd1 vccd1 _14038_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17866_ _20639_/Q _17866_/A1 _17883_/S vssd1 vssd1 vccd1 vccd1 _20639_/D sky130_fd_sc_hd__mux2_1
XFILLER_239_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1372 _12455_/Y vssd1 vssd1 vccd1 vccd1 _12565_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1383 _11642_/S0 vssd1 vssd1 vccd1 vccd1 _11936_/S sky130_fd_sc_hd__buf_6
Xfanout1394 _11698_/B2 vssd1 vssd1 vccd1 vccd1 _12097_/S sky130_fd_sc_hd__clkbuf_8
X_19605_ _19606_/CLK _19605_/D vssd1 vssd1 vccd1 vccd1 _19605_/Q sky130_fd_sc_hd__dfxtp_1
X_16817_ _19224_/Q _17003_/B _16964_/B1 _19093_/Q _16816_/X vssd1 vssd1 vccd1 vccd1
+ _16817_/X sky130_fd_sc_hd__o221a_1
XFILLER_238_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17797_ _20574_/Q _17937_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20574_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19536_ _19603_/CLK _19536_/D vssd1 vssd1 vccd1 vccd1 _19536_/Q sky130_fd_sc_hd__dfxtp_1
X_16748_ _16746_/X _16747_/X _12930_/B vssd1 vssd1 vccd1 vccd1 _16748_/X sky130_fd_sc_hd__a21bo_1
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19467_ _20687_/CLK _19467_/D vssd1 vssd1 vccd1 vccd1 _19467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16679_ _19934_/Q _17751_/A1 _16704_/S vssd1 vssd1 vccd1 vccd1 _19934_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18418_ _18418_/A _18418_/B vssd1 vssd1 vccd1 vccd1 _20863_/D sky130_fd_sc_hd__and2_1
XFILLER_167_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19398_ _20704_/CLK _19398_/D vssd1 vssd1 vccd1 vccd1 _19398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18349_ _18502_/B _18349_/B vssd1 vssd1 vccd1 vccd1 _18349_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20311_ _21047_/A _20311_/D vssd1 vssd1 vccd1 vccd1 _20311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput60 dout0[25] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput71 dout0[35] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput82 dout0[45] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_2
Xinput93 dout0[55] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_2
X_20242_ _20296_/CLK _20242_/D vssd1 vssd1 vccd1 vccd1 _20242_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20173_ _20708_/CLK _20173_/D vssd1 vssd1 vccd1 vccd1 _20173_/Q sky130_fd_sc_hd__dfxtp_1
X_09984_ _12138_/A1 _16063_/B2 _09983_/X vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__a21oi_2
XFILLER_103_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10690_ _10688_/X _10689_/X _12414_/S vssd1 vssd1 vccd1 vccd1 _10690_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12360_ _12433_/A1 _17951_/A1 _12359_/X _09750_/Y vssd1 vssd1 vccd1 vccd1 _16037_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ _12342_/A _11294_/X _11310_/X vssd1 vssd1 vccd1 vccd1 _11311_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_153_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20509_ _20641_/CLK _20509_/D vssd1 vssd1 vccd1 vccd1 _20509_/Q sky130_fd_sc_hd__dfxtp_1
X_12291_ _19558_/Q _12365_/A2 _11225_/B _19622_/Q vssd1 vssd1 vccd1 vccd1 _12291_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14030_ _19209_/Q _14099_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _14030_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11242_ _11242_/A1 _14011_/A2 _11241_/X _11242_/B1 _19847_/Q vssd1 vssd1 vccd1 vccd1
+ _11242_/X sky130_fd_sc_hd__o32a_1
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11173_ _12311_/A1 _11168_/X _11172_/X vssd1 vssd1 vccd1 vccd1 _11173_/X sky130_fd_sc_hd__o21a_1
XFILLER_268_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10124_ _11236_/B _10124_/B vssd1 vssd1 vccd1 vccd1 _10124_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15981_ _15981_/A _15981_/B vssd1 vssd1 vccd1 vccd1 _15981_/X sky130_fd_sc_hd__or2_1
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ _20501_/Q _17894_/A1 _17742_/S vssd1 vssd1 vccd1 vccd1 _20501_/D sky130_fd_sc_hd__mux2_1
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932_ _15019_/B _15019_/C vssd1 vssd1 vccd1 vccd1 _15314_/C sky130_fd_sc_hd__nand2_8
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10055_ _19877_/Q _19778_/Q _10428_/S vssd1 vssd1 vccd1 vccd1 _10055_/X sky130_fd_sc_hd__mux2_1
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _20437_/Q _17928_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20437_/D sky130_fd_sc_hd__mux2_1
XFILLER_236_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _14860_/X _14862_/Y _15061_/S vssd1 vssd1 vccd1 vccd1 _15114_/B sky130_fd_sc_hd__mux2_1
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ _16596_/X _16601_/X _16567_/A vssd1 vssd1 vccd1 vccd1 _16602_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13814_ _13816_/A1 _13738_/B _13816_/B1 input230/X vssd1 vssd1 vccd1 vccd1 _13814_/X
+ sky130_fd_sc_hd__a22o_1
X_17582_ _20340_/Q _17893_/A1 _17606_/S vssd1 vssd1 vccd1 vccd1 _20340_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14794_ _19144_/Q _14798_/A2 _14793_/X _14794_/C1 vssd1 vssd1 vccd1 vccd1 _19521_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19321_ _19956_/CLK _19321_/D vssd1 vssd1 vccd1 vccd1 _19321_/Q sky130_fd_sc_hd__dfxtp_1
X_16533_ _16551_/A _16533_/B vssd1 vssd1 vccd1 vccd1 _19832_/D sky130_fd_sc_hd__or2_1
XFILLER_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13745_ _13765_/A _13745_/B vssd1 vssd1 vccd1 vccd1 _13745_/X sky130_fd_sc_hd__and2_2
X_10957_ _12429_/A1 _10956_/X _10955_/X vssd1 vssd1 vccd1 vccd1 _10957_/X sky130_fd_sc_hd__o21a_1
XFILLER_250_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19252_ _20273_/CLK _19252_/D vssd1 vssd1 vccd1 vccd1 _19252_/Q sky130_fd_sc_hd__dfxtp_1
X_16464_ _19773_/Q _17684_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19773_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13676_ _13718_/A _13676_/B vssd1 vssd1 vccd1 vccd1 _13676_/Y sky130_fd_sc_hd__nor2_1
X_10888_ _10373_/A _10033_/Y _09659_/B vssd1 vssd1 vccd1 vccd1 _10888_/X sky130_fd_sc_hd__a21o_1
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18203_ _19536_/Q _18213_/B vssd1 vssd1 vccd1 vccd1 _18203_/Y sky130_fd_sc_hd__nand2b_4
X_15415_ _20731_/Q _15445_/A2 _15445_/B1 _20763_/Q vssd1 vssd1 vccd1 vccd1 _15415_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19183_ _19560_/CLK _19183_/D vssd1 vssd1 vccd1 vccd1 _19183_/Q sky130_fd_sc_hd__dfxtp_1
X_12627_ _12628_/A _12628_/B vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__nand2_1
X_16395_ _18064_/A _16395_/B _16396_/B vssd1 vssd1 vccd1 vccd1 _19743_/D sky130_fd_sc_hd__nor3_1
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18134_ _18134_/A _19107_/Q vssd1 vssd1 vccd1 vccd1 _18322_/C sky130_fd_sc_hd__and2_1
X_15346_ _15282_/A _16794_/B _15331_/Y vssd1 vssd1 vccd1 vccd1 _15346_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _13635_/A _13653_/A vssd1 vssd1 vccd1 vccd1 _12558_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18065_ _20761_/Q _18063_/B _18064_/Y vssd1 vssd1 vccd1 vccd1 _20761_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11509_ _19678_/Q _20166_/Q _11527_/S vssd1 vssd1 vccd1 vccd1 _11509_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15277_ _17287_/A _15482_/A2 _15270_/X _15276_/X vssd1 vssd1 vccd1 vccd1 _15277_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12489_ _13863_/A _12490_/B vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__and2_4
X_17016_ _19994_/Q _18985_/A _17015_/B _12927_/B _17849_/S vssd1 vssd1 vccd1 vccd1
+ _19994_/D sky130_fd_sc_hd__a41o_1
X_14228_ _19505_/Q _14229_/B vssd1 vssd1 vccd1 vccd1 _14240_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _14157_/Y _14159_/B vssd1 vssd1 vccd1 vccd1 _14162_/A sky130_fd_sc_hd__and2b_1
XFILLER_171_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout609 _14599_/S vssd1 vssd1 vccd1 vccd1 _14598_/S sky130_fd_sc_hd__buf_12
XFILLER_112_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18967_ _19114_/Q _18974_/A2 _18967_/B1 _13181_/A vssd1 vssd1 vccd1 vccd1 _18968_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_47_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20179_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17918_ _17918_/A _17918_/B vssd1 vssd1 vccd1 vccd1 _17919_/C sky130_fd_sc_hd__nor2_1
XFILLER_267_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18898_ _18980_/A _18898_/B vssd1 vssd1 vccd1 vccd1 _20999_/D sky130_fd_sc_hd__nor2_1
XFILLER_255_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1180 _12516_/Y vssd1 vssd1 vccd1 vccd1 _13602_/A1 sky130_fd_sc_hd__buf_8
XFILLER_254_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1191 _09643_/Y vssd1 vssd1 vccd1 vccd1 _10561_/A sky130_fd_sc_hd__buf_6
XFILLER_82_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17849_ _20624_/Q input250/X _17849_/S vssd1 vssd1 vccd1 vccd1 _20624_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20860_ _20860_/CLK _20860_/D vssd1 vssd1 vccd1 vccd1 _20860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19519_ _21009_/CLK _19519_/D vssd1 vssd1 vccd1 vccd1 _19519_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_263_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20791_ _21020_/CLK _20791_/D vssd1 vssd1 vccd1 vccd1 _20791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20225_ _20818_/CLK _20225_/D vssd1 vssd1 vccd1 vccd1 _20225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20156_ _20563_/CLK _20156_/D vssd1 vssd1 vccd1 vccd1 _20156_/Q sky130_fd_sc_hd__dfxtp_1
X_09967_ _12138_/A1 _20513_/Q _11988_/S _09949_/X vssd1 vssd1 vccd1 vccd1 _09967_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20087_ _20561_/CLK _20087_/D vssd1 vssd1 vccd1 vccd1 _20087_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _12134_/S _09897_/X _09896_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _09898_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_503 _20624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _11946_/A1 _19358_/Q _20713_/Q _11860_/B2 _11946_/C1 vssd1 vssd1 vccd1 vccd1
+ _11860_/X sky130_fd_sc_hd__a221o_1
XFILLER_73_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_514 input221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_525 _19494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_536 _17949_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_547 ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ _11061_/A _16079_/A vssd1 vssd1 vccd1 vccd1 _10811_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_558 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11791_ _11791_/A _11791_/B _13421_/A vssd1 vssd1 vccd1 vccd1 _11792_/B sky130_fd_sc_hd__nand3_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20989_ _21023_/CLK _20989_/D vssd1 vssd1 vccd1 vccd1 _20989_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_569 _13780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13530_ _20919_/Q _13598_/A2 _13575_/C _13529_/X _14110_/A vssd1 vssd1 vccd1 vccd1
+ _13530_/X sky130_fd_sc_hd__a221o_1
X_10742_ _20371_/Q _20435_/Q _12381_/S vssd1 vssd1 vccd1 vccd1 _10742_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10673_ _10671_/X _10672_/X _12391_/S vssd1 vssd1 vccd1 vccd1 _10673_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13461_ _16232_/B _13462_/B vssd1 vssd1 vccd1 vccd1 _16278_/B sky130_fd_sc_hd__nand2b_1
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15200_ _17248_/A _15199_/X _15452_/S vssd1 vssd1 vccd1 vccd1 _15200_/X sky130_fd_sc_hd__mux2_1
X_12412_ _19396_/Q _12412_/A2 _12410_/X _12412_/B2 _12411_/X vssd1 vssd1 vccd1 vccd1
+ _12412_/X sky130_fd_sc_hd__o221a_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16180_ _19614_/Q _15834_/X _16190_/S vssd1 vssd1 vccd1 vccd1 _16181_/B sky130_fd_sc_hd__mux2_1
XFILLER_127_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13392_ _13323_/C _13255_/B _13390_/X _13391_/X vssd1 vssd1 vccd1 vccd1 _13392_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_138_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15131_ _20724_/Q _15445_/A2 _15445_/B1 _20756_/Q vssd1 vssd1 vccd1 vccd1 _15131_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12343_ _20149_/Q _20117_/Q _12346_/S vssd1 vssd1 vccd1 vccd1 _12343_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12274_ _12265_/A _12269_/Y _12271_/Y _12273_/Y _12431_/A1 vssd1 vssd1 vccd1 vccd1
+ _12274_/X sky130_fd_sc_hd__a221o_1
X_15062_ _14818_/X _14822_/X _15062_/S vssd1 vssd1 vccd1 vccd1 _15062_/X sky130_fd_sc_hd__mux2_2
XFILLER_182_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14013_ _12584_/C _14031_/A2 _14040_/B1 _14012_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1
+ _19171_/D sky130_fd_sc_hd__o221a_1
X_11225_ _19591_/Q _11225_/B vssd1 vssd1 vccd1 vccd1 _11225_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19870_ _20630_/CLK _19870_/D vssd1 vssd1 vccd1 vccd1 _19870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11156_ _19624_/Q _19930_/Q _12296_/S vssd1 vssd1 vccd1 vccd1 _11156_/X sky130_fd_sc_hd__mux2_1
X_18821_ _18821_/A _18821_/B vssd1 vssd1 vccd1 vccd1 _20988_/D sky130_fd_sc_hd__nor2_1
XFILLER_268_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10107_ _12088_/S _10106_/X _11396_/S vssd1 vssd1 vccd1 vccd1 _10107_/X sky130_fd_sc_hd__o21a_1
X_18752_ _18752_/A _18752_/B vssd1 vssd1 vccd1 vccd1 _20976_/D sky130_fd_sc_hd__and2_1
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ _11085_/X _11086_/X _12317_/S vssd1 vssd1 vccd1 vccd1 _11087_/X sky130_fd_sc_hd__mux2_1
X_15964_ _20878_/Q _16018_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15964_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput250 localMemory_wb_sel_i[3] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_hd__clkbuf_2
Xinput261 manufacturerID[7] vssd1 vssd1 vccd1 vccd1 input261/X sky130_fd_sc_hd__buf_2
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17703_ _20487_/Q _17806_/A1 _17703_/S vssd1 vssd1 vccd1 vccd1 _20487_/D sky130_fd_sc_hd__mux2_1
Xinput272 partID[2] vssd1 vssd1 vccd1 vccd1 input272/X sky130_fd_sc_hd__clkbuf_2
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10038_ input127/X input163/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10038_/X sky130_fd_sc_hd__mux2_8
X_14915_ _18148_/S _14915_/B vssd1 vssd1 vccd1 vccd1 _14915_/X sky130_fd_sc_hd__and2b_1
XFILLER_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput283 versionID[3] vssd1 vssd1 vccd1 vccd1 input283/X sky130_fd_sc_hd__buf_2
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18683_ _19524_/Q _18683_/B vssd1 vssd1 vccd1 vccd1 _18683_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15895_ _13439_/C _15894_/X _15895_/S vssd1 vssd1 vccd1 vccd1 _15895_/X sky130_fd_sc_hd__mux2_1
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _20390_/Q _17805_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20390_/D sky130_fd_sc_hd__mux2_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14846_ _09861_/B _10636_/Y _14882_/B vssd1 vssd1 vccd1 vccd1 _14846_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17565_ _20325_/Q _17944_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20325_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14777_ _19513_/Q _14797_/B vssd1 vssd1 vccd1 vccd1 _14777_/X sky130_fd_sc_hd__or2_1
XFILLER_44_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11989_ _12144_/A1 _11988_/X _11985_/X _12144_/C1 vssd1 vssd1 vccd1 vccd1 _11989_/X
+ sky130_fd_sc_hd__o211a_1
X_19304_ _20463_/CLK _19304_/D vssd1 vssd1 vccd1 vccd1 _19304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16516_ _19823_/Q _17945_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19823_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13728_ _13798_/A1 _13767_/B _13727_/X vssd1 vssd1 vccd1 vccd1 _13729_/B sky130_fd_sc_hd__a21oi_4
XFILLER_56_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17496_ _20283_/Q _17502_/B vssd1 vssd1 vccd1 vccd1 _17496_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_165_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21006_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_231_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19235_ _19520_/CLK _19235_/D vssd1 vssd1 vccd1 vccd1 _19235_/Q sky130_fd_sc_hd__dfxtp_4
X_16447_ _19763_/Q _16450_/C _18801_/A vssd1 vssd1 vccd1 vccd1 _16447_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_220_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13659_ _13659_/A _13659_/B vssd1 vssd1 vccd1 vccd1 _13660_/B sky130_fd_sc_hd__nor2_8
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19166_ _20659_/CLK _19166_/D vssd1 vssd1 vccd1 vccd1 _19166_/Q sky130_fd_sc_hd__dfxtp_4
X_16378_ _19736_/Q _19737_/Q _16378_/C vssd1 vssd1 vccd1 vccd1 _16380_/B sky130_fd_sc_hd__and3_1
XFILLER_173_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18117_ _20781_/Q _20780_/Q _18117_/C vssd1 vssd1 vccd1 vccd1 _18122_/C sky130_fd_sc_hd__and3_4
X_15329_ _10766_/Y _15328_/X _15591_/A vssd1 vssd1 vccd1 vccd1 _15329_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19097_ _19621_/CLK _19097_/D vssd1 vssd1 vccd1 vccd1 _19097_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_184_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18048_ _18048_/A _18053_/C vssd1 vssd1 vccd1 vccd1 _18048_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20010_ _20751_/CLK _20010_/D vssd1 vssd1 vccd1 vccd1 _20010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09821_ _09819_/X _09820_/X _12071_/S vssd1 vssd1 vccd1 vccd1 _09821_/X sky130_fd_sc_hd__mux2_1
X_19999_ _20624_/CLK _19999_/D vssd1 vssd1 vccd1 vccd1 _19999_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_86_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09752_ _09752_/A _19325_/Q _12003_/C vssd1 vssd1 vccd1 vccd1 _09752_/X sky130_fd_sc_hd__or3_1
XFILLER_228_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09683_ _10020_/B _09678_/X _09682_/Y _09592_/A _09592_/C vssd1 vssd1 vccd1 vccd1
+ _09683_/X sky130_fd_sc_hd__o221a_4
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20912_ _21010_/CLK _20912_/D vssd1 vssd1 vccd1 vccd1 _20912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _21006_/CLK _20843_/D vssd1 vssd1 vccd1 vccd1 _20843_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20774_ _21029_/CLK _20774_/D vssd1 vssd1 vccd1 vccd1 _20774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_278_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11010_ _11275_/A _11006_/X _11009_/X _12311_/C1 vssd1 vssd1 vccd1 vccd1 _11010_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_132_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20208_ _20766_/CLK _20208_/D vssd1 vssd1 vccd1 vccd1 _20208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1905 _13887_/C1 vssd1 vssd1 vccd1 vccd1 fanout1905/X sky130_fd_sc_hd__clkbuf_8
Xfanout1916 _18726_/A vssd1 vssd1 vccd1 vccd1 _18720_/A sky130_fd_sc_hd__buf_4
Xfanout1927 _16193_/A vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__buf_4
XFILLER_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout940 _15292_/S vssd1 vssd1 vccd1 vccd1 _15215_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_132_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1938 _09515_/Y vssd1 vssd1 vccd1 vccd1 _14185_/C1 sky130_fd_sc_hd__buf_4
XFILLER_104_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1949 _16381_/B1 vssd1 vssd1 vccd1 vccd1 _17241_/C1 sky130_fd_sc_hd__buf_4
XFILLER_237_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout951 _14233_/S vssd1 vssd1 vccd1 vccd1 _14202_/S sky130_fd_sc_hd__buf_6
X_20139_ _20482_/CLK _20139_/D vssd1 vssd1 vccd1 vccd1 _20139_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout962 _17861_/A1 vssd1 vssd1 vccd1 vccd1 _17929_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout973 _10386_/X vssd1 vssd1 vccd1 vccd1 split4/A sky130_fd_sc_hd__buf_6
XFILLER_285_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout984 _10128_/X vssd1 vssd1 vccd1 vccd1 _17199_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 _17003_/B vssd1 vssd1 vccd1 vccd1 _16980_/A2 sky130_fd_sc_hd__buf_4
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12961_ _19248_/Q _19247_/Q vssd1 vssd1 vccd1 vccd1 _12961_/X sky130_fd_sc_hd__or2_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _19459_/Q _17706_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19459_/D sky130_fd_sc_hd__mux2_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _19648_/Q _11915_/S _11897_/X _11528_/S vssd1 vssd1 vccd1 vccd1 _11912_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15680_ _13427_/A _15982_/C _16056_/B1 vssd1 vssd1 vccd1 vccd1 _15680_/X sky130_fd_sc_hd__a21o_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12892_ _12911_/A _12893_/B vssd1 vssd1 vccd1 vccd1 _13209_/B sky130_fd_sc_hd__nand2_1
XANTENNA_300 input228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_311 input239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_322 _13510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _19395_/Q _17915_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19395_/D sky130_fd_sc_hd__mux2_1
XFILLER_233_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 _19494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11843_ _11922_/A1 _11842_/Y _12158_/B1 vssd1 vssd1 vccd1 vccd1 _11843_/X sky130_fd_sc_hd__o21a_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_344 _14732_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_355 _09936_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_366 _12513_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _20223_/Q _17356_/A2 _17362_/B1 _20272_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17350_/X sky130_fd_sc_hd__a221o_1
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_377 _15678_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14562_ _19332_/Q _17707_/A1 _14562_/S vssd1 vssd1 vccd1 vccd1 _19332_/D sky130_fd_sc_hd__mux2_1
XANTENNA_388 _16824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11774_ _11774_/A _11774_/B vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_399 _16719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _19708_/Q _16298_/B _18414_/A vssd1 vssd1 vccd1 vccd1 _16302_/B sky130_fd_sc_hd__o21ai_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _12664_/C _13512_/X _12982_/B vssd1 vssd1 vccd1 vccd1 _13513_/Y sky130_fd_sc_hd__a21oi_2
X_17281_ _17281_/A _17290_/B _17290_/C vssd1 vssd1 vccd1 vccd1 _17281_/X sky130_fd_sc_hd__and3_1
X_10725_ _09672_/A _13960_/A2 _10724_/X _11239_/B1 _19837_/Q vssd1 vssd1 vccd1 vccd1
+ _16081_/A sky130_fd_sc_hd__o32ai_4
XFILLER_202_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _19271_/Q _17890_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19271_/D sky130_fd_sc_hd__mux2_1
X_19020_ _18245_/Y _19048_/A2 _19017_/X _12552_/C _19048_/C1 vssd1 vssd1 vccd1 vccd1
+ _19020_/X sky130_fd_sc_hd__a221o_1
XFILLER_202_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16232_ _16241_/A _16232_/B vssd1 vssd1 vccd1 vccd1 _19695_/D sky130_fd_sc_hd__nor2_2
X_13444_ _16598_/B vssd1 vssd1 vccd1 vccd1 _13463_/C sky130_fd_sc_hd__inv_4
X_10656_ _20340_/Q _12295_/B vssd1 vssd1 vccd1 vccd1 _10656_/X sky130_fd_sc_hd__or2_1
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16163_ _19605_/Q _16164_/B _16162_/Y _16165_/C1 vssd1 vssd1 vccd1 vccd1 _19605_/D
+ sky130_fd_sc_hd__o211a_1
X_10587_ _19632_/Q _19938_/Q _11676_/S vssd1 vssd1 vccd1 vccd1 _10587_/X sky130_fd_sc_hd__mux2_1
X_13375_ _13281_/A _12748_/B _13281_/B _12749_/C vssd1 vssd1 vccd1 vccd1 _13377_/B
+ sky130_fd_sc_hd__a31o_1
X_15114_ _15155_/S _15114_/B vssd1 vssd1 vccd1 vccd1 _15114_/Y sky130_fd_sc_hd__nor2_1
X_12326_ _12400_/A1 _12318_/X _12325_/X _12311_/X vssd1 vssd1 vccd1 vccd1 _12326_/X
+ sky130_fd_sc_hd__o31a_4
XFILLER_155_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16094_ _10026_/X _16106_/A2 _16093_/X vssd1 vssd1 vccd1 vccd1 _19571_/D sky130_fd_sc_hd__o21a_1
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19922_ _20682_/CLK _19922_/D vssd1 vssd1 vccd1 vccd1 _19922_/Q sky130_fd_sc_hd__dfxtp_1
X_15045_ _15043_/X _15044_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _15045_/X sky130_fd_sc_hd__mux2_1
X_12257_ _12255_/X _12256_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _12257_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ _12430_/S _11208_/B vssd1 vssd1 vccd1 vccd1 _11208_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19853_ _20862_/CLK _19853_/D vssd1 vssd1 vccd1 vccd1 _19853_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_214_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12188_ _19893_/Q _19794_/Q _12188_/S vssd1 vssd1 vccd1 vccd1 _12189_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18804_ _19123_/Q _18949_/A2 _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18804_/Y sky130_fd_sc_hd__a21oi_1
X_11139_ _11140_/B vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__inv_2
XFILLER_68_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16996_ _19245_/Q _16996_/A2 _16996_/B1 _19114_/Q _16995_/X vssd1 vssd1 vccd1 vccd1
+ _16996_/X sky130_fd_sc_hd__o221a_1
X_19784_ _20081_/CLK _19784_/D vssd1 vssd1 vccd1 vccd1 _19784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18735_ _20968_/Q _18270_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18736_/B sky130_fd_sc_hd__mux2_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15947_ _15976_/B2 _15946_/X _15930_/X _15526_/B vssd1 vssd1 vccd1 vccd1 _15947_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18666_ _20940_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18666_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _20971_/Q _16045_/A2 _16016_/S _20843_/Q _15877_/X vssd1 vssd1 vccd1 vccd1
+ _15878_/X sky130_fd_sc_hd__a221o_1
XFILLER_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17617_ _20373_/Q _17928_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20373_/D sky130_fd_sc_hd__mux2_1
XFILLER_221_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14829_ _10802_/B _11958_/B _14882_/B vssd1 vssd1 vccd1 vccd1 _14829_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18597_ _18490_/X _18621_/A2 _18595_/Y _18596_/Y vssd1 vssd1 vccd1 vccd1 _18598_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17548_ _20308_/Q _17684_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20308_/D sky130_fd_sc_hd__mux2_1
XFILLER_233_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17479_ _17487_/A1 _17478_/Y _18048_/A vssd1 vssd1 vccd1 vccd1 _20274_/D sky130_fd_sc_hd__a21oi_1
XFILLER_221_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19218_ _19219_/CLK _19218_/D vssd1 vssd1 vccd1 vccd1 _19218_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20490_ _20491_/CLK _20490_/D vssd1 vssd1 vccd1 vccd1 _20490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19149_ _19228_/CLK _19149_/D vssd1 vssd1 vccd1 vccd1 _19149_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20655_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21042_ _21042_/CLK _21042_/D vssd1 vssd1 vccd1 vccd1 _21042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ _09802_/X _09803_/X _09806_/S vssd1 vssd1 vccd1 vccd1 _09804_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09735_ _12504_/A _10979_/C vssd1 vssd1 vccd1 vccd1 _09735_/Y sky130_fd_sc_hd__nand2_8
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09666_ _19574_/Q _09666_/B vssd1 vssd1 vccd1 vccd1 _09680_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09609_/A _19091_/Q vssd1 vssd1 vccd1 vccd1 _16454_/A sky130_fd_sc_hd__and2b_4
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ _20863_/CLK _20826_/D vssd1 vssd1 vccd1 vccd1 _20826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20757_ _20757_/CLK _20757_/D vssd1 vssd1 vccd1 vccd1 _20757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10510_ _19408_/Q _20567_/Q _10518_/S vssd1 vssd1 vccd1 vccd1 _10510_/X sky130_fd_sc_hd__mux2_1
X_11490_ _11851_/C _11489_/X _11486_/X _12191_/C1 vssd1 vssd1 vccd1 vccd1 _11490_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20688_ _20688_/CLK _20688_/D vssd1 vssd1 vccd1 vccd1 _20688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ _19940_/Q _12068_/C1 _12044_/B _12071_/S vssd1 vssd1 vccd1 vccd1 _10441_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10372_ _19570_/Q _10371_/X _11243_/S vssd1 vssd1 vccd1 vccd1 _10372_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13160_ _11415_/A _13422_/B _10276_/Y vssd1 vssd1 vccd1 vccd1 _13421_/B sky130_fd_sc_hd__a21oi_4
XFILLER_109_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12111_ _12109_/Y _12111_/B vssd1 vssd1 vccd1 vccd1 _13432_/A sky130_fd_sc_hd__nand2b_4
Xclkbuf_4_10__f_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_59_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_237_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13091_ _13091_/A _13091_/B _13091_/C vssd1 vssd1 vccd1 vccd1 _13091_/X sky130_fd_sc_hd__and3_1
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12042_ _20551_/Q _12064_/S vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__or2_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1702 _11191_/A vssd1 vssd1 vccd1 vccd1 _12254_/A sky130_fd_sc_hd__buf_8
Xfanout1713 _11537_/A1 vssd1 vssd1 vccd1 vccd1 _12270_/B1 sky130_fd_sc_hd__buf_4
Xfanout1724 _12752_/A vssd1 vssd1 vccd1 vccd1 _10581_/A1 sky130_fd_sc_hd__buf_6
XFILLER_104_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16850_ _19973_/Q _16849_/A _16849_/Y _16896_/C1 vssd1 vssd1 vccd1 vccd1 _19973_/D
+ sky130_fd_sc_hd__a211o_1
Xfanout1735 _12123_/C1 vssd1 vssd1 vccd1 vccd1 _11892_/C1 sky130_fd_sc_hd__buf_6
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1746 _09502_/Y vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__buf_12
XFILLER_66_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1757 _11243_/S vssd1 vssd1 vccd1 vccd1 _11229_/S sky130_fd_sc_hd__buf_8
XFILLER_120_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout770 _18902_/A vssd1 vssd1 vccd1 vccd1 _18683_/B sky130_fd_sc_hd__buf_6
X_15801_ _20904_/Q _16043_/A2 _16043_/B1 _15800_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _15801_/X sky130_fd_sc_hd__a221o_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1768 _13275_/A1 vssd1 vssd1 vccd1 vccd1 _13373_/A sky130_fd_sc_hd__buf_4
XFILLER_266_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout781 _14110_/A vssd1 vssd1 vccd1 vccd1 _18760_/B sky130_fd_sc_hd__buf_4
Xfanout1779 _20262_/Q vssd1 vssd1 vccd1 vccd1 _17442_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_59_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16781_ _16726_/X _16780_/Y _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16781_/X sky130_fd_sc_hd__a21o_2
XFILLER_1_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout792 _13350_/A vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__buf_6
X_13993_ _14041_/A1 _09664_/B _09664_/C _14041_/B1 _19846_/Q vssd1 vssd1 vccd1 vccd1
+ _14075_/C sky130_fd_sc_hd__o32a_1
XFILLER_280_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18520_ _18671_/B _18520_/B vssd1 vssd1 vccd1 vccd1 _18520_/X sky130_fd_sc_hd__or2_1
XFILLER_219_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15732_ _15732_/A _15732_/B _15814_/A vssd1 vssd1 vccd1 vccd1 _15732_/X sky130_fd_sc_hd__or3b_1
X_12944_ _12944_/A _14906_/B _12944_/C _14912_/B vssd1 vssd1 vccd1 vccd1 _12945_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _20880_/Q _18310_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18452_/B sky130_fd_sc_hd__mux2_1
XFILLER_234_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15663_ _20867_/Q _16042_/A2 fanout819/X vssd1 vssd1 vccd1 vccd1 _15663_/X sky130_fd_sc_hd__o21ba_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12875_ _19518_/Q _12916_/A2 _12874_/X _12916_/B2 vssd1 vssd1 vccd1 vccd1 _12877_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_130 _13669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_141 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17402_ _17402_/A _17438_/B vssd1 vssd1 vccd1 vccd1 _17402_/Y sky130_fd_sc_hd__nand2_2
XFILLER_60_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_152 _13770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14614_ _19378_/Q _17898_/A1 _14628_/S vssd1 vssd1 vccd1 vccd1 _19378_/D sky130_fd_sc_hd__mux2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_163 _13853_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ _11981_/C1 _11825_/X _11822_/X _12137_/C1 vssd1 vssd1 vccd1 vccd1 _11826_/X
+ sky130_fd_sc_hd__a211o_4
X_18382_ _20846_/Q _18385_/B _18381_/Y _18748_/A vssd1 vssd1 vccd1 vccd1 _20846_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _19111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15594_ _16002_/A1 _15593_/Y _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15594_/X sky130_fd_sc_hd__a21o_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_196 _19549_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17333_ _17402_/A _13844_/B _17336_/B _17236_/Y _17430_/A vssd1 vssd1 vccd1 vccd1
+ _17333_/X sky130_fd_sc_hd__a41o_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _19315_/Q _17097_/A1 _14562_/S vssd1 vssd1 vccd1 vccd1 _19315_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _13422_/A _11757_/B vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_53_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17264_ _20193_/Q _17330_/A2 _17279_/C1 vssd1 vssd1 vccd1 vccd1 _17264_/X sky130_fd_sc_hd__a21o_1
X_10708_ _10705_/X _10706_/X _10707_/X _12357_/A1 _12265_/A vssd1 vssd1 vccd1 vccd1
+ _10708_/X sky130_fd_sc_hd__a221o_1
XFILLER_187_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14476_ _18718_/A _14476_/B vssd1 vssd1 vccd1 vccd1 _19262_/D sky130_fd_sc_hd__and2_1
X_11688_ _19545_/Q _12365_/A2 _09607_/X _19609_/Q vssd1 vssd1 vccd1 vccd1 _11688_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19003_ _21021_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _19003_/X sky130_fd_sc_hd__or2_1
X_16215_ _19638_/Q _17099_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19638_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13427_ _13427_/A _13427_/B _13427_/C _13427_/D vssd1 vssd1 vccd1 vccd1 _13428_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_127_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17195_ _20159_/Q _17861_/A1 _17212_/S vssd1 vssd1 vccd1 vccd1 _20159_/D sky130_fd_sc_hd__mux2_1
X_10639_ _13459_/A _13611_/A _13596_/A vssd1 vssd1 vccd1 vccd1 _10645_/A sky130_fd_sc_hd__nor3_4
X_16146_ _16784_/B _16194_/S vssd1 vssd1 vccd1 vccd1 _16146_/Y sky130_fd_sc_hd__nand2_1
X_13358_ _14295_/C1 _09496_/Y _16241_/A _13357_/X vssd1 vssd1 vccd1 vccd1 _13359_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_170_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12309_ _12307_/X _12308_/X _12309_/S vssd1 vssd1 vccd1 vccd1 _12309_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ _16077_/A _16077_/B vssd1 vssd1 vccd1 vccd1 _16077_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13289_ split6/X _13283_/X _13288_/X vssd1 vssd1 vccd1 vccd1 _13289_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19905_ _20658_/CLK _19905_/D vssd1 vssd1 vccd1 vccd1 _19905_/Q sky130_fd_sc_hd__dfxtp_1
X_15028_ _15246_/A _15028_/B vssd1 vssd1 vccd1 vccd1 _15028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19836_ _20268_/CLK _19836_/D vssd1 vssd1 vccd1 vccd1 _19836_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_111_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19767_ _20638_/CLK _19767_/D vssd1 vssd1 vccd1 vccd1 _19767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput3 coreIndex[2] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_6
X_16979_ _20425_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16979_/X sky130_fd_sc_hd__a21o_2
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09520_ input65/X vssd1 vssd1 vccd1 vccd1 _09520_/Y sky130_fd_sc_hd__inv_2
X_18718_ _18718_/A _18718_/B vssd1 vssd1 vccd1 vccd1 _20959_/D sky130_fd_sc_hd__and2_1
XFILLER_65_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19698_ _19698_/CLK _19698_/D vssd1 vssd1 vccd1 vccd1 _19698_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_180_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20296_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_252_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18649_ _18973_/A _18649_/B vssd1 vssd1 vccd1 vccd1 _20935_/D sky130_fd_sc_hd__nor2_1
XFILLER_225_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20611_ _20647_/CLK _20611_/D vssd1 vssd1 vccd1 vccd1 _20611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20542_ _20646_/CLK _20542_/D vssd1 vssd1 vccd1 vccd1 _20542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20473_ _20701_/CLK _20473_/D vssd1 vssd1 vccd1 vccd1 _20473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput340 _13702_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[15] sky130_fd_sc_hd__buf_4
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput351 _13750_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[25] sky130_fd_sc_hd__buf_4
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput362 _13660_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[6] sky130_fd_sc_hd__buf_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput373 _13475_/X vssd1 vssd1 vccd1 vccd1 csb0[1] sky130_fd_sc_hd__buf_4
XFILLER_248_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput384 _13808_/X vssd1 vssd1 vccd1 vccd1 din0[17] sky130_fd_sc_hd__buf_4
Xfanout1009 _15259_/B vssd1 vssd1 vccd1 vccd1 _15982_/C sky130_fd_sc_hd__buf_4
Xoutput395 _13818_/X vssd1 vssd1 vccd1 vccd1 din0[27] sky130_fd_sc_hd__buf_4
XFILLER_99_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21025_ _21025_/CLK _21025_/D vssd1 vssd1 vccd1 vccd1 _21025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ _11980_/S _09717_/X _09716_/X _12144_/A1 vssd1 vssd1 vccd1 vccd1 _09718_/X
+ sky130_fd_sc_hd__a211o_1
X_10990_ _20153_/Q _12213_/B vssd1 vssd1 vccd1 vccd1 _10990_/X sky130_fd_sc_hd__or2_1
XFILLER_215_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09649_ _19862_/Q _19660_/Q _20019_/Q vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__or3b_4
XFILLER_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _19497_/Q _12758_/B vssd1 vssd1 vccd1 vccd1 _12662_/C sky130_fd_sc_hd__nand2_1
XFILLER_163_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _19546_/Q _12155_/A2 _12155_/B1 _19610_/Q vssd1 vssd1 vccd1 vccd1 _11611_/X
+ sky130_fd_sc_hd__a22o_1
X_20809_ _21029_/CLK _20809_/D vssd1 vssd1 vccd1 vccd1 _20809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12591_ _13657_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _12591_/X sky130_fd_sc_hd__or2_4
XFILLER_169_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14330_ _20287_/Q _14330_/A2 _14330_/B1 input228/X vssd1 vssd1 vccd1 vccd1 _14332_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11542_ _09986_/A _20381_/Q _20445_/Q _09928_/S vssd1 vssd1 vccd1 vccd1 _11542_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ _14260_/A _14260_/B _14260_/C vssd1 vssd1 vccd1 vccd1 _14271_/B sky130_fd_sc_hd__a21o_1
X_11473_ _11849_/S _11472_/X _11471_/X _12183_/C1 vssd1 vssd1 vccd1 vccd1 _11473_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16000_ _16000_/A1 _15989_/X _15990_/X _15999_/X vssd1 vssd1 vccd1 vccd1 _16000_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13212_ _13114_/B _13212_/B _13323_/C vssd1 vssd1 vccd1 vccd1 _13212_/X sky130_fd_sc_hd__and3b_1
XFILLER_136_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10424_ _10430_/S _10422_/X _10423_/X vssd1 vssd1 vccd1 vccd1 _10424_/X sky130_fd_sc_hd__o21a_1
X_14192_ _14188_/B _14191_/Y _14202_/S vssd1 vssd1 vccd1 vccd1 _14192_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13143_ _15071_/S _13143_/B vssd1 vssd1 vccd1 vccd1 _13482_/B sky130_fd_sc_hd__nor2_2
X_10355_ _10356_/A _19911_/Q _10518_/S _20036_/Q vssd1 vssd1 vccd1 vccd1 _10355_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ _20720_/Q _17951_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20720_/D sky130_fd_sc_hd__mux2_1
X_10286_ _10032_/Y _10285_/Y _09638_/Y vssd1 vssd1 vccd1 vccd1 _10286_/X sky130_fd_sc_hd__a21o_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13074_ _13033_/X _13073_/Y _13034_/Y vssd1 vssd1 vccd1 vccd1 _13354_/A sky130_fd_sc_hd__a21boi_4
XFILLER_285_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1510 _11599_/S vssd1 vssd1 vccd1 vccd1 _11979_/S sky130_fd_sc_hd__buf_6
X_16902_ _16885_/A _16901_/X _16866_/B2 vssd1 vssd1 vccd1 vccd1 _16902_/Y sky130_fd_sc_hd__o21bai_4
X_12025_ _19425_/Q _20584_/Q _12025_/S vssd1 vssd1 vccd1 vccd1 _12025_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17882_ _20655_/Q _17916_/A1 _17882_/S vssd1 vssd1 vccd1 vccd1 _20655_/D sky130_fd_sc_hd__mux2_1
Xfanout1521 fanout1522/X vssd1 vssd1 vccd1 vccd1 _11987_/S sky130_fd_sc_hd__buf_4
Xfanout1532 _12064_/S vssd1 vssd1 vccd1 vccd1 _11676_/S sky130_fd_sc_hd__buf_6
XFILLER_250_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1543 _10316_/S vssd1 vssd1 vccd1 vccd1 _10137_/C sky130_fd_sc_hd__clkbuf_8
Xfanout1554 _11090_/S vssd1 vssd1 vccd1 vccd1 _11093_/S sky130_fd_sc_hd__buf_6
XFILLER_265_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1565 fanout1566/X vssd1 vssd1 vccd1 vccd1 _10842_/S sky130_fd_sc_hd__buf_4
X_19621_ _19621_/CLK _19621_/D vssd1 vssd1 vccd1 vccd1 _19621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16833_ _16878_/A _16833_/B vssd1 vssd1 vccd1 vccd1 _16833_/Y sky130_fd_sc_hd__nand2_1
Xfanout1576 _11597_/C1 vssd1 vssd1 vccd1 vccd1 _12151_/A1 sky130_fd_sc_hd__buf_8
Xfanout1587 _11600_/C1 vssd1 vssd1 vccd1 vccd1 _12144_/A1 sky130_fd_sc_hd__buf_8
XFILLER_281_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1598 _11833_/C1 vssd1 vssd1 vccd1 vccd1 _11528_/S sky130_fd_sc_hd__buf_6
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16764_ _20401_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16764_/X sky130_fd_sc_hd__a21o_1
X_19552_ _19552_/CLK _19552_/D vssd1 vssd1 vccd1 vccd1 _19552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13976_ _19191_/Q _14063_/C _14003_/S vssd1 vssd1 vccd1 vccd1 _13976_/X sky130_fd_sc_hd__mux2_1
XFILLER_253_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15715_ _19721_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15715_/X sky130_fd_sc_hd__or2_1
X_18503_ _20894_/Q _18474_/S _18502_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18504_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12927_ _17015_/B _12927_/B vssd1 vssd1 vccd1 vccd1 _13466_/B sky130_fd_sc_hd__nand2_4
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19483_ _20710_/CLK _19483_/D vssd1 vssd1 vccd1 vccd1 _19483_/Q sky130_fd_sc_hd__dfxtp_1
X_16695_ _19950_/Q _17835_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19950_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18434_ _18734_/A _18434_/B vssd1 vssd1 vccd1 vccd1 _20871_/D sky130_fd_sc_hd__and2_1
X_15646_ _16052_/A1 _15644_/Y _15645_/X _13427_/C _15975_/B2 vssd1 vssd1 vccd1 vccd1
+ _15646_/X sky130_fd_sc_hd__a32o_1
X_12858_ _15703_/B2 _12856_/X _12857_/X vssd1 vssd1 vccd1 vccd1 _12860_/B sky130_fd_sc_hd__o21a_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ _20549_/Q _12139_/S vssd1 vssd1 vccd1 vccd1 _11809_/X sky130_fd_sc_hd__or2_1
X_18365_ _18526_/B _18375_/B vssd1 vssd1 vccd1 vccd1 _18365_/Y sky130_fd_sc_hd__nand2_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15577_ _15289_/X _15291_/X _15577_/S vssd1 vssd1 vccd1 vccd1 _15577_/X sky130_fd_sc_hd__mux2_1
X_12789_ _12790_/C _12790_/D vssd1 vssd1 vccd1 vccd1 _13586_/B sky130_fd_sc_hd__nor2_1
XFILLER_187_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _20211_/Q _17328_/A2 _17315_/X _18416_/A vssd1 vssd1 vccd1 vccd1 _20211_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14528_ _14528_/A _16454_/B vssd1 vssd1 vccd1 vccd1 _17918_/A sky130_fd_sc_hd__or2_4
XFILLER_30_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18296_ _20813_/Q _18295_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18297_/B sky130_fd_sc_hd__mux2_1
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17247_ _20188_/Q _17268_/A2 _17245_/X _17246_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1
+ _20188_/D sky130_fd_sc_hd__o221a_1
X_14459_ _20225_/Q _19254_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14460_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17178_ _20144_/Q _17178_/A1 _17178_/S vssd1 vssd1 vccd1 vccd1 _20144_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16129_ _19589_/Q _16131_/A2 _16129_/B1 vssd1 vssd1 vccd1 vccd1 _16129_/X sky130_fd_sc_hd__o21a_1
XFILLER_277_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19819_ _20645_/CLK _19819_/D vssd1 vssd1 vccd1 vccd1 _19819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ _09503_/A vssd1 vssd1 vccd1 vccd1 _09503_/Y sky130_fd_sc_hd__inv_6
XFILLER_225_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 _15861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 _16811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_52 _16953_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_63 _18195_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20525_ _20657_/CLK _20525_/D vssd1 vssd1 vccd1 vccd1 _20525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_74 _09618_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_85 _11452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_96 _12402_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20456_ _20580_/CLK _20456_/D vssd1 vssd1 vccd1 vccd1 _20456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20387_ _20451_/CLK _20387_/D vssd1 vssd1 vccd1 vccd1 _20387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ _11336_/A _10129_/X _10130_/X vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10071_ _12060_/A1 _19314_/Q _11680_/C1 _09806_/S vssd1 vssd1 vccd1 vccd1 _10071_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21008_ _21008_/CLK _21008_/D vssd1 vssd1 vccd1 vccd1 _21008_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13830_ _20000_/Q _13473_/X _13784_/X split2/X vssd1 vssd1 vccd1 vccd1 _13830_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_275_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13761_ _12157_/Y _13742_/B _13776_/B1 vssd1 vssd1 vccd1 vccd1 _13764_/A sky130_fd_sc_hd__o21a_2
X_10973_ _10553_/B _10382_/Y _10972_/X _10373_/X vssd1 vssd1 vccd1 vccd1 _10973_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15500_ _15500_/A0 _15264_/B _15500_/S vssd1 vssd1 vccd1 vccd1 _15500_/X sky130_fd_sc_hd__mux2_1
XFILLER_216_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12712_ _12706_/Y _12707_/X _12709_/X _12711_/Y vssd1 vssd1 vccd1 vccd1 _12726_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_280_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _19789_/Q _17666_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19789_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _16598_/C _13692_/B vssd1 vssd1 vccd1 vccd1 _13692_/Y sky130_fd_sc_hd__nor2_1
XFILLER_243_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15431_ _10600_/Y _15430_/X _15591_/A vssd1 vssd1 vccd1 vccd1 _15431_/Y sky130_fd_sc_hd__o21ai_4
X_12643_ _19500_/Q _12758_/B vssd1 vssd1 vccd1 vccd1 _12643_/X sky130_fd_sc_hd__and2_1
XFILLER_157_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18150_ _18149_/S _19114_/Q _14912_/X vssd1 vssd1 vccd1 vccd1 _18318_/C sky130_fd_sc_hd__a21o_1
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15362_ _14841_/S _14840_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _15362_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_169_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12574_ _12574_/A _12574_/B _12580_/B vssd1 vssd1 vccd1 vccd1 _12577_/B sky130_fd_sc_hd__nor3_2
XFILLER_157_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17101_ _20071_/Q _17903_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20071_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14313_ _14314_/A _14314_/B vssd1 vssd1 vccd1 vccd1 _14315_/B sky130_fd_sc_hd__and2_1
X_18081_ _20767_/Q _18079_/B _18080_/Y vssd1 vssd1 vccd1 vccd1 _20767_/D sky130_fd_sc_hd__o21a_1
XFILLER_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ _11902_/S _11524_/X _11523_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _11525_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15293_ _15291_/X _15292_/X _15577_/S vssd1 vssd1 vccd1 vccd1 _15293_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17032_ _20010_/Q input196/X _17040_/S vssd1 vssd1 vccd1 vccd1 _20010_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14244_ _14244_/A1 _14243_/X _13319_/Y vssd1 vssd1 vccd1 vccd1 _14245_/C sky130_fd_sc_hd__o21a_1
X_11456_ _11922_/A1 _13707_/A _12158_/B1 vssd1 vssd1 vccd1 vccd1 _11456_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ _20408_/Q _20344_/Q _20636_/Q _20600_/Q _12081_/S0 _10405_/C vssd1 vssd1
+ vccd1 vccd1 _10407_/X sky130_fd_sc_hd__mux4_1
X_14175_ _20272_/Q _14237_/A2 _14216_/B1 input243/X vssd1 vssd1 vccd1 vccd1 _14177_/B
+ sky130_fd_sc_hd__a22o_4
X_11387_ _19806_/Q _11392_/A2 _11385_/X _09738_/A _11386_/X vssd1 vssd1 vccd1 vccd1
+ _11387_/X sky130_fd_sc_hd__o221a_1
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ _17532_/A _13941_/A vssd1 vssd1 vccd1 vccd1 _13242_/A sky130_fd_sc_hd__nor2_1
X_10338_ _20315_/Q _11295_/S _10337_/X vssd1 vssd1 vccd1 vccd1 _10338_/X sky130_fd_sc_hd__a21o_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18983_ _18985_/B _18983_/B vssd1 vssd1 vccd1 vccd1 _18983_/Y sky130_fd_sc_hd__nand2_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21016_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _20950_/Q _20884_/Q vssd1 vssd1 vccd1 vccd1 _13517_/B sky130_fd_sc_hd__nand2_1
X_17934_ _20703_/Q _17934_/A1 _17934_/S vssd1 vssd1 vccd1 vccd1 _20703_/D sky130_fd_sc_hd__mux2_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _20412_/Q _20348_/Q _20640_/Q _20604_/Q _11035_/S _11021_/C vssd1 vssd1 vccd1
+ vccd1 _10269_/X sky130_fd_sc_hd__mux4_1
XFILLER_285_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1340 _09688_/Y vssd1 vssd1 vccd1 vccd1 _11009_/A2 sky130_fd_sc_hd__buf_2
XFILLER_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12008_ _12008_/A _20684_/Q _12008_/C vssd1 vssd1 vccd1 vccd1 _12008_/X sky130_fd_sc_hd__or3_1
Xfanout1351 _17038_/S vssd1 vssd1 vccd1 vccd1 _17026_/S sky130_fd_sc_hd__buf_2
XFILLER_39_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1362 _13853_/Y vssd1 vssd1 vccd1 vccd1 _14002_/B1 sky130_fd_sc_hd__clkbuf_8
X_17865_ _20638_/Q _17899_/A1 _17883_/S vssd1 vssd1 vccd1 vccd1 _20638_/D sky130_fd_sc_hd__mux2_1
XFILLER_266_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1373 _11213_/B vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__buf_6
XFILLER_282_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1384 _11642_/S0 vssd1 vssd1 vccd1 vccd1 _12013_/S sky130_fd_sc_hd__clkbuf_8
X_19604_ _19606_/CLK _19604_/D vssd1 vssd1 vccd1 vccd1 _19604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1395 _11698_/B2 vssd1 vssd1 vccd1 vccd1 _12025_/S sky130_fd_sc_hd__clkbuf_8
X_16816_ _20406_/Q _16963_/A2 _16963_/B1 vssd1 vssd1 vccd1 vccd1 _16816_/X sky130_fd_sc_hd__a21o_1
X_17796_ _20573_/Q _17936_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20573_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19535_ _19606_/CLK _19535_/D vssd1 vssd1 vccd1 vccd1 _19535_/Q sky130_fd_sc_hd__dfxtp_2
X_13959_ _19153_/Q _19050_/S _14043_/B1 _13958_/X _16097_/B1 vssd1 vssd1 vccd1 vccd1
+ _19153_/D sky130_fd_sc_hd__o221a_1
X_16747_ _17219_/B _16743_/Y _16745_/X _12952_/X vssd1 vssd1 vccd1 vccd1 _16747_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19466_ _20561_/CLK _19466_/D vssd1 vssd1 vccd1 vccd1 _19466_/Q sky130_fd_sc_hd__dfxtp_1
X_16678_ _19933_/Q _17750_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19933_/D sky130_fd_sc_hd__mux2_1
XFILLER_222_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18417_ _20863_/Q _18225_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18418_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15629_ _15626_/Y _15628_/X _15625_/Y vssd1 vssd1 vccd1 vccd1 _15629_/Y sky130_fd_sc_hd__a21oi_1
X_19397_ _20688_/CLK _19397_/D vssd1 vssd1 vccd1 vccd1 _19397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18348_ _20829_/Q _18349_/B _18347_/Y _18714_/A vssd1 vssd1 vccd1 vccd1 _20829_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18279_ _18299_/A1 _14364_/B _18278_/Y vssd1 vssd1 vccd1 vccd1 _18538_/B sky130_fd_sc_hd__o21ai_4
XFILLER_174_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20310_ _20679_/CLK _20310_/D vssd1 vssd1 vccd1 vccd1 _20310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput50 dout0[16] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_2
XFILLER_238_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput61 dout0[26] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput72 dout0[36] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput83 dout0[46] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_2
X_20241_ _21010_/CLK _20241_/D vssd1 vssd1 vccd1 vccd1 _20241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput94 dout0[56] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_2
XFILLER_254_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20172_ _20568_/CLK _20172_/D vssd1 vssd1 vccd1 vccd1 _20172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09983_ _11922_/A1 _13722_/A _12158_/B1 vssd1 vssd1 vccd1 vccd1 _09983_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11310_ _12504_/A _11301_/X _11309_/X _11396_/S vssd1 vssd1 vccd1 vccd1 _11310_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_5_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20508_ _20672_/CLK _20508_/D vssd1 vssd1 vccd1 vccd1 _20508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12290_ _12290_/A _15955_/A _12290_/C _12290_/D vssd1 vssd1 vccd1 vccd1 _12454_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11241_ input114/X input149/X _11241_/S vssd1 vssd1 vccd1 vccd1 _11241_/X sky130_fd_sc_hd__mux2_8
X_20439_ _21047_/A _20439_/D vssd1 vssd1 vccd1 vccd1 _20439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11172_ _11169_/X _11170_/X _11171_/X _10152_/S _09621_/A vssd1 vssd1 vccd1 vccd1
+ _11172_/X sky130_fd_sc_hd__a221o_1
XFILLER_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_212_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20047_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10123_ _19588_/Q _10122_/X _11229_/S vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__mux2_2
X_15980_ _19555_/Q _15980_/A2 _15979_/X _16191_/A vssd1 vssd1 vccd1 vccd1 _19555_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14931_ _14955_/B _15133_/B vssd1 vssd1 vccd1 vccd1 _15019_/C sky130_fd_sc_hd__nor2_4
X_10054_ _10052_/X _10053_/X _10585_/S vssd1 vssd1 vccd1 vccd1 _10054_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17650_ _20436_/Q _17684_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20436_/D sky130_fd_sc_hd__mux2_1
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14862_ _14862_/A vssd1 vssd1 vccd1 vccd1 _14862_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ _13463_/C _13765_/A _16598_/A vssd1 vssd1 vccd1 vccd1 _16601_/X sky130_fd_sc_hd__a21o_1
X_13813_ _13816_/A1 _13733_/B _13816_/B1 input229/X vssd1 vssd1 vccd1 vccd1 _13813_/X
+ sky130_fd_sc_hd__a22o_1
X_17581_ _20339_/Q _17892_/A1 _17606_/S vssd1 vssd1 vccd1 vccd1 _20339_/D sky130_fd_sc_hd__mux2_1
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14793_ _19521_/Q _14797_/B vssd1 vssd1 vccd1 vccd1 _14793_/X sky130_fd_sc_hd__or2_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16532_ _19832_/Q _16566_/A2 _16566_/B1 input21/X vssd1 vssd1 vccd1 vccd1 _16533_/B
+ sky130_fd_sc_hd__o22a_1
X_19320_ _20081_/CLK _19320_/D vssd1 vssd1 vccd1 vccd1 _19320_/Q sky130_fd_sc_hd__dfxtp_1
X_13744_ _13744_/A _13744_/B vssd1 vssd1 vccd1 vccd1 _13745_/B sky130_fd_sc_hd__nor2_8
X_10956_ _19402_/Q _20561_/Q _12346_/S vssd1 vssd1 vccd1 vccd1 _10956_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16463_ _19772_/Q _17683_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19772_/D sky130_fd_sc_hd__mux2_1
X_19251_ _20184_/CLK _19251_/D vssd1 vssd1 vccd1 vccd1 _19251_/Q sky130_fd_sc_hd__dfxtp_1
X_13675_ _13675_/A _13675_/B _13675_/C _13684_/B vssd1 vssd1 vccd1 vccd1 _13675_/Y
+ sky130_fd_sc_hd__nand4_4
X_10887_ _19531_/Q _09613_/A _18152_/C _19595_/Q vssd1 vssd1 vccd1 vccd1 _10887_/X
+ sky130_fd_sc_hd__a22o_1
X_15414_ _19711_/Q _15595_/A2 _15595_/B1 _19743_/Q vssd1 vssd1 vccd1 vccd1 _15414_/X
+ sky130_fd_sc_hd__a22o_1
X_18202_ _19051_/A _18202_/B vssd1 vssd1 vccd1 vccd1 _20794_/D sky130_fd_sc_hd__nor2_1
XFILLER_176_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19182_ _19560_/CLK _19182_/D vssd1 vssd1 vccd1 vccd1 _19182_/Q sky130_fd_sc_hd__dfxtp_1
X_12626_ _19523_/Q _12916_/A2 _12625_/X _12916_/B2 vssd1 vssd1 vccd1 vccd1 _12628_/B
+ sky130_fd_sc_hd__o22a_1
X_16394_ _19742_/Q _19743_/Q _16394_/C vssd1 vssd1 vccd1 vccd1 _16396_/B sky130_fd_sc_hd__and3_1
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18133_ _12959_/B _19106_/Q _18134_/A vssd1 vssd1 vccd1 vccd1 _18323_/B sky130_fd_sc_hd__mux2_2
X_15345_ _15396_/A1 _15332_/X _15344_/X vssd1 vssd1 vccd1 vccd1 _16794_/B sky130_fd_sc_hd__a21oi_4
XFILLER_156_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _12587_/A _18462_/B vssd1 vssd1 vccd1 vccd1 _12557_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18064_ _18064_/A _18069_/C vssd1 vssd1 vccd1 vccd1 _18064_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11508_ _11983_/A1 _19478_/Q _19446_/Q _11916_/S _11892_/C1 vssd1 vssd1 vccd1 vccd1
+ _11508_/X sky130_fd_sc_hd__a221o_1
X_15276_ _20791_/Q _15016_/A _15021_/X _15275_/X vssd1 vssd1 vccd1 vccd1 _15276_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_89_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12488_ split8/A _12847_/A2 _15948_/A1 vssd1 vssd1 vccd1 vccd1 _12488_/X sky130_fd_sc_hd__a21o_4
XFILLER_176_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17015_ _18821_/A _17015_/B _17015_/C vssd1 vssd1 vccd1 vccd1 _17015_/Y sky130_fd_sc_hd__nor3_1
X_14227_ _20277_/Q _14237_/A2 _14267_/B1 input217/X vssd1 vssd1 vccd1 vccd1 _14229_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_7_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11439_ _12150_/S _11438_/X _11437_/X _12140_/C1 vssd1 vssd1 vccd1 vccd1 _11439_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_160_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14158_ _19498_/Q _14158_/B vssd1 vssd1 vccd1 vccd1 _14159_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13109_ _20944_/Q _13363_/B _18667_/B vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__a21o_1
XFILLER_112_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14089_ _14105_/A _14107_/B _14089_/C vssd1 vssd1 vccd1 vccd1 _14089_/X sky130_fd_sc_hd__or3_1
XFILLER_26_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18966_ _18966_/A _18966_/B vssd1 vssd1 vccd1 vccd1 _21009_/D sky130_fd_sc_hd__nor2_1
XFILLER_86_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17917_ _20688_/Q _17917_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20688_/D sky130_fd_sc_hd__mux2_1
XFILLER_255_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18897_ _18523_/X _18978_/B _18895_/X _18896_/Y vssd1 vssd1 vccd1 vccd1 _18898_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_239_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1170 _14897_/Y vssd1 vssd1 vccd1 vccd1 _15282_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1181 _12516_/Y vssd1 vssd1 vccd1 vccd1 _13598_/A2 sky130_fd_sc_hd__clkbuf_4
X_17848_ _20623_/Q input249/X _17849_/S vssd1 vssd1 vccd1 vccd1 _20623_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1192 _12403_/A1 vssd1 vssd1 vccd1 vccd1 _11922_/A1 sky130_fd_sc_hd__buf_4
XFILLER_226_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _21044_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_17779_ _17919_/A _17919_/B _17779_/C vssd1 vssd1 vccd1 vccd1 _17779_/X sky130_fd_sc_hd__and3_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19518_ _20291_/CLK _19518_/D vssd1 vssd1 vccd1 vccd1 _19518_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20790_ _20863_/CLK _20790_/D vssd1 vssd1 vccd1 vccd1 _20790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_wb_clk_i _20408_/CLK vssd1 vssd1 vccd1 vccd1 _20669_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_241_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19449_ _20081_/CLK _19449_/D vssd1 vssd1 vccd1 vccd1 _19449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20224_ _20818_/CLK _20224_/D vssd1 vssd1 vccd1 vccd1 _20224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20155_ _20155_/CLK _20155_/D vssd1 vssd1 vccd1 vccd1 _20155_/Q sky130_fd_sc_hd__dfxtp_1
X_09966_ _11981_/C1 _09965_/X _09962_/X _12137_/C1 vssd1 vssd1 vccd1 vccd1 _09966_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_134_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20086_ _20557_/CLK _20086_/D vssd1 vssd1 vccd1 vccd1 _20086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _19819_/Q _19323_/Q _12149_/S vssd1 vssd1 vccd1 vccd1 _09897_/X sky130_fd_sc_hd__mux2_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_504 _20624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_515 input240/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_526 _19504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _09672_/A _13960_/A2 _10809_/X _11228_/B1 _19836_/Q vssd1 vssd1 vccd1 vccd1
+ _16079_/A sky130_fd_sc_hd__o32ai_4
XANTENNA_537 _13473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_548 ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11790_ _13424_/A _11790_/B vssd1 vssd1 vccd1 vccd1 _15551_/A sky130_fd_sc_hd__xnor2_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_559 _15365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20988_ _21022_/CLK _20988_/D vssd1 vssd1 vccd1 vccd1 _20988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ _20467_/Q _20307_/Q _12219_/S vssd1 vssd1 vccd1 vccd1 _10741_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13460_ _13612_/A split3/A _13459_/Y _13458_/Y _13244_/X vssd1 vssd1 vccd1 vccd1
+ _13462_/B sky130_fd_sc_hd__a32o_4
X_10672_ _19805_/Q _19309_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10672_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12411_ _12411_/A _20687_/Q _12411_/C vssd1 vssd1 vccd1 vccd1 _12411_/X sky130_fd_sc_hd__or3_1
XFILLER_199_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13391_ _20936_/Q _13363_/B _18683_/B vssd1 vssd1 vccd1 vccd1 _13391_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15130_ _19704_/Q _15475_/A2 _15475_/B1 _19736_/Q vssd1 vssd1 vccd1 vccd1 _15130_/X
+ sky130_fd_sc_hd__a22o_1
X_12342_ _12342_/A _12342_/B vssd1 vssd1 vccd1 vccd1 _12342_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15061_ _14819_/X _14829_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _15061_/X sky130_fd_sc_hd__mux2_1
X_12273_ _12420_/B1 _12272_/X _12265_/A vssd1 vssd1 vccd1 vccd1 _12273_/Y sky130_fd_sc_hd__a21oi_1
X_14012_ _19203_/Q _14087_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _14012_/X sky130_fd_sc_hd__mux2_1
X_11224_ _15071_/S _11224_/B vssd1 vssd1 vccd1 vccd1 _13636_/A sky130_fd_sc_hd__or2_4
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18820_ _18490_/X _18819_/B _18818_/X _18819_/Y vssd1 vssd1 vccd1 vccd1 _18821_/B
+ sky130_fd_sc_hd__o211a_1
X_11155_ _12301_/S _11155_/B _11155_/C vssd1 vssd1 vccd1 vccd1 _11155_/X sky130_fd_sc_hd__or3_1
XFILLER_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10106_ _10104_/X _10105_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _10106_/X sky130_fd_sc_hd__mux2_1
XFILLER_249_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18751_ _20976_/Q _18310_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18752_/B sky130_fd_sc_hd__mux2_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11086_ _19368_/Q _20659_/Q _11161_/S vssd1 vssd1 vccd1 vccd1 _11086_/X sky130_fd_sc_hd__mux2_1
X_15963_ _20750_/Q _16011_/A2 _16011_/B1 _20782_/Q vssd1 vssd1 vccd1 vccd1 _15963_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput240 localMemory_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_hd__buf_12
XFILLER_48_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput251 localMemory_wb_stb_i vssd1 vssd1 vccd1 vccd1 _17014_/B sky130_fd_sc_hd__clkbuf_2
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ _20486_/Q _17805_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20486_/D sky130_fd_sc_hd__mux2_1
Xinput262 manufacturerID[8] vssd1 vssd1 vccd1 vccd1 _17263_/A sky130_fd_sc_hd__buf_2
X_14914_ _14951_/A _14951_/B vssd1 vssd1 vccd1 vccd1 _15022_/A sky130_fd_sc_hd__nand2_4
X_10037_ _11236_/B _10037_/B vssd1 vssd1 vccd1 vccd1 _10037_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_49_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput273 partID[3] vssd1 vssd1 vccd1 vccd1 _17281_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18682_ _20944_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18682_/Y sky130_fd_sc_hd__nand2_1
X_15894_ _15948_/A1 _12884_/Y _15893_/X _15921_/B2 vssd1 vssd1 vccd1 vccd1 _15894_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput284 wb_rst_i vssd1 vssd1 vccd1 vccd1 _16278_/A sky130_fd_sc_hd__buf_12
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _20389_/Q _17804_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20389_/D sky130_fd_sc_hd__mux2_1
XFILLER_236_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14845_ _11799_/B _11404_/B _14882_/B vssd1 vssd1 vccd1 vccd1 _14845_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17564_ _20324_/Q _17943_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20324_/D sky130_fd_sc_hd__mux2_1
X_14776_ _19135_/Q _14798_/A2 _14775_/X _14776_/C1 vssd1 vssd1 vccd1 vccd1 _19512_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_251_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11988_ _11986_/X _11987_/X _11988_/S vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19303_ _20670_/CLK _19303_/D vssd1 vssd1 vccd1 vccd1 _19303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16515_ _19822_/Q _17876_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19822_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13727_ _13659_/A _13688_/X _13655_/B _13714_/S vssd1 vssd1 vccd1 vccd1 _13727_/X
+ sky130_fd_sc_hd__o211a_1
X_10939_ _19627_/Q _19933_/Q _19271_/Q _20058_/Q _11211_/S _11021_/C vssd1 vssd1 vccd1
+ vccd1 _10939_/X sky130_fd_sc_hd__mux4_1
XFILLER_260_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17495_ _17495_/A1 _17494_/Y _18863_/A vssd1 vssd1 vccd1 vccd1 _20282_/D sky130_fd_sc_hd__a21oi_1
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19234_ _19523_/CLK _19234_/D vssd1 vssd1 vccd1 vccd1 _19234_/Q sky130_fd_sc_hd__dfxtp_2
X_13658_ _13658_/A _13694_/C vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__or2_4
X_16446_ _19762_/Q _16444_/B _16445_/Y vssd1 vssd1 vccd1 vccd1 _19762_/D sky130_fd_sc_hd__o21a_1
XFILLER_231_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _19515_/Q _12811_/A vssd1 vssd1 vccd1 vccd1 _12804_/B sky130_fd_sc_hd__and2_2
X_16377_ _19736_/Q _16378_/C _19737_/Q vssd1 vssd1 vccd1 vccd1 _16379_/B sky130_fd_sc_hd__a21oi_1
X_19165_ _19704_/CLK _19165_/D vssd1 vssd1 vccd1 vccd1 _19165_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13589_ _13589_/A1 _13585_/Y _13586_/X _13588_/X vssd1 vssd1 vccd1 vccd1 _13589_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15328_ _12578_/B _12639_/X _15327_/X _10935_/B vssd1 vssd1 vccd1 vccd1 _15328_/X
+ sky130_fd_sc_hd__o211a_1
X_18116_ _20780_/Q _18117_/C _20781_/Q vssd1 vssd1 vccd1 vccd1 _18118_/B sky130_fd_sc_hd__a21oi_1
XFILLER_129_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19096_ _20721_/CLK _19096_/D vssd1 vssd1 vccd1 vccd1 _19096_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_134_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _20184_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18047_ _20755_/Q _18047_/B vssd1 vssd1 vccd1 vccd1 _18053_/C sky130_fd_sc_hd__and2_2
X_15259_ _15259_/A _15259_/B vssd1 vssd1 vccd1 vccd1 _15259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09820_ _19289_/Q _20076_/Q _11682_/S vssd1 vssd1 vccd1 vccd1 _09820_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19998_ _20624_/CLK _19998_/D vssd1 vssd1 vccd1 vccd1 _19998_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09751_ _09752_/A _19920_/Q _11932_/S0 _20045_/Q vssd1 vssd1 vccd1 vccd1 _09751_/X
+ sky130_fd_sc_hd__o22a_1
X_18949_ _19144_/Q _18949_/A2 _18949_/B1 vssd1 vssd1 vccd1 vccd1 _18949_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09682_ _09659_/B _09679_/X _09680_/X _09681_/X vssd1 vssd1 vccd1 vccd1 _09682_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_239_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20911_ _21009_/CLK _20911_/D vssd1 vssd1 vccd1 vccd1 _20911_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20842_ _21000_/CLK _20842_/D vssd1 vssd1 vccd1 vccd1 _20842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20773_ _21029_/CLK _20773_/D vssd1 vssd1 vccd1 vccd1 _20773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20207_ _20766_/CLK _20207_/D vssd1 vssd1 vccd1 vccd1 _20207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1906 _16167_/C1 vssd1 vssd1 vccd1 vccd1 _16189_/A sky130_fd_sc_hd__buf_4
XFILLER_278_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1917 _18726_/A vssd1 vssd1 vccd1 vccd1 _18718_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout930 _14933_/Y vssd1 vssd1 vccd1 vccd1 _15595_/A2 sky130_fd_sc_hd__buf_4
Xfanout1928 _14070_/C1 vssd1 vssd1 vccd1 vccd1 _16193_/A sky130_fd_sc_hd__buf_4
Xfanout1939 _16131_/B1 vssd1 vssd1 vccd1 vccd1 _16127_/B1 sky130_fd_sc_hd__buf_4
Xfanout941 _11137_/A vssd1 vssd1 vccd1 vccd1 _15292_/S sky130_fd_sc_hd__clkbuf_8
Xfanout952 _14121_/X vssd1 vssd1 vccd1 vccd1 _14233_/S sky130_fd_sc_hd__buf_4
X_20138_ _20481_/CLK _20138_/D vssd1 vssd1 vccd1 vccd1 _20138_/Q sky130_fd_sc_hd__dfxtp_1
X_09949_ _20545_/Q _12124_/S vssd1 vssd1 vccd1 vccd1 _09949_/X sky130_fd_sc_hd__or2_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout963 _17861_/A1 vssd1 vssd1 vccd1 vccd1 _17686_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_237_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout974 _17691_/A1 vssd1 vssd1 vccd1 vccd1 _17934_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_258_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout985 _10128_/X vssd1 vssd1 vccd1 vccd1 _17899_/A1 sky130_fd_sc_hd__buf_6
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20069_ _20692_/CLK _20069_/D vssd1 vssd1 vccd1 vccd1 _20069_/Q sky130_fd_sc_hd__dfxtp_1
X_12960_ _19995_/Q _19996_/Q _12930_/B vssd1 vssd1 vccd1 vccd1 _12960_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout996 _16709_/X vssd1 vssd1 vccd1 vccd1 _17003_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_218_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _11513_/S _11910_/X _11909_/X _12144_/A1 vssd1 vssd1 vccd1 vccd1 _11911_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_273_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _19520_/Q _12857_/B _12890_/X _15921_/B2 vssd1 vssd1 vccd1 vccd1 _12893_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_301 input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 input240/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _19394_/Q _17914_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19394_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _12157_/A1 _17876_/A1 _11841_/X _12153_/B1 vssd1 vssd1 vccd1 vccd1 _11842_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA_323 _13540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 _19494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 _14099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_356 _11033_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _19331_/Q _17915_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19331_/D sky130_fd_sc_hd__mux2_1
XFILLER_242_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_367 _12513_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11773_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _11773_/X sky130_fd_sc_hd__and2_1
XANTENNA_378 _15678_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_389 _16860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _19707_/Q _19708_/Q _16300_/C vssd1 vssd1 vccd1 vccd1 _16306_/C sky130_fd_sc_hd__and3_2
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ _13526_/B _13512_/B vssd1 vssd1 vccd1 vccd1 _13512_/X sky130_fd_sc_hd__or2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _20199_/Q _17280_/A2 _17279_/X _17331_/C1 vssd1 vssd1 vccd1 vccd1 _20199_/D
+ sky130_fd_sc_hd__o211a_1
X_10724_ input167/X input138/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10724_/X sky130_fd_sc_hd__mux2_8
XFILLER_159_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _19270_/Q _17855_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19270_/D sky130_fd_sc_hd__mux2_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16231_ _19654_/Q _17674_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19654_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13443_ _16066_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _16598_/B sky130_fd_sc_hd__nand2_8
X_10655_ _10651_/X _10654_/X _12377_/S vssd1 vssd1 vccd1 vccd1 _10655_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16162_ _16860_/B _16164_/B vssd1 vssd1 vccd1 vccd1 _16162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13374_ _13373_/A _19235_/Q _14780_/C1 _13373_/Y vssd1 vssd1 vccd1 vccd1 _13388_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_70_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10586_ _11684_/A1 _10585_/X _10582_/X _12073_/A1 vssd1 vssd1 vccd1 vccd1 _10586_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15113_ _14847_/X _14859_/X _15170_/A vssd1 vssd1 vccd1 vccd1 _15113_/X sky130_fd_sc_hd__mux2_1
X_12325_ _12398_/C1 _12324_/X _12321_/X _12399_/C1 vssd1 vssd1 vccd1 vccd1 _12325_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16093_ _19571_/Q _16081_/B _16107_/B1 vssd1 vssd1 vccd1 vccd1 _16093_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19921_ _20681_/CLK _19921_/D vssd1 vssd1 vccd1 vccd1 _19921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15044_ _14849_/X _14853_/X _15062_/S vssd1 vssd1 vccd1 vccd1 _15044_/X sky130_fd_sc_hd__mux2_1
X_12256_ _20426_/Q _20362_/Q _20654_/Q _20618_/Q _12339_/S0 _12337_/C vssd1 vssd1
+ vccd1 vccd1 _12256_/X sky130_fd_sc_hd__mux4_1
XFILLER_269_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11207_ _09507_/A _11205_/X _11206_/X vssd1 vssd1 vccd1 vccd1 _11208_/B sky130_fd_sc_hd__o21ai_1
X_19852_ _20017_/CLK _19852_/D vssd1 vssd1 vccd1 vccd1 _19852_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_141_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12187_ _19490_/Q _19458_/Q _12188_/S vssd1 vssd1 vccd1 vccd1 _12187_/X sky130_fd_sc_hd__mux2_1
XFILLER_256_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18803_ _18830_/A _18803_/B vssd1 vssd1 vccd1 vccd1 _18803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11138_ _15254_/S _11138_/B vssd1 vssd1 vccd1 vccd1 _11140_/B sky130_fd_sc_hd__and2_1
XFILLER_228_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19783_ _20574_/CLK _19783_/D vssd1 vssd1 vccd1 vccd1 _19783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16995_ _20427_/Q _17004_/A2 _17004_/B1 vssd1 vssd1 vccd1 vccd1 _16995_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18734_ _18734_/A _18734_/B vssd1 vssd1 vccd1 vccd1 _20967_/D sky130_fd_sc_hd__and2_1
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ _19400_/Q _11074_/S _11068_/X _12371_/C1 vssd1 vssd1 vccd1 vccd1 _11069_/X
+ sky130_fd_sc_hd__o211a_1
X_15946_ _16024_/A1 _15944_/X _15945_/Y _15949_/B _15975_/B2 vssd1 vssd1 vccd1 vccd1
+ _15946_/X sky130_fd_sc_hd__a32o_1
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18665_ _18966_/A _18665_/B vssd1 vssd1 vccd1 vccd1 _20939_/D sky130_fd_sc_hd__nor2_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ _20939_/Q _15995_/A2 _15876_/X vssd1 vssd1 vccd1 vccd1 _15877_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17616_ _20372_/Q _17684_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20372_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14828_ _14826_/X _14827_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _14828_/X sky130_fd_sc_hd__mux2_1
X_18596_ _19502_/Q _18604_/B vssd1 vssd1 vccd1 vccd1 _18596_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17547_ _20307_/Q _17683_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20307_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14759_ _19504_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14759_/X sky130_fd_sc_hd__or2_1
XFILLER_233_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17478_ _20274_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17478_/Y sky130_fd_sc_hd__nand2_1
X_19217_ _19219_/CLK _19217_/D vssd1 vssd1 vccd1 vccd1 _19217_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16429_ _18096_/A _16434_/C vssd1 vssd1 vccd1 vccd1 _16429_/Y sky130_fd_sc_hd__nor2_1
XFILLER_146_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19148_ _20300_/CLK _19148_/D vssd1 vssd1 vccd1 vccd1 _19148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19079_ _20424_/Q vssd1 vssd1 vccd1 vccd1 _20424_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21041_ _21041_/CLK _21041_/D vssd1 vssd1 vccd1 vccd1 _21041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09803_ _20140_/Q _20108_/Q _10428_/S vssd1 vssd1 vccd1 vccd1 _09803_/X sky130_fd_sc_hd__mux2_1
XFILLER_259_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09734_ _10260_/S _09734_/B vssd1 vssd1 vccd1 vccd1 _09734_/Y sky130_fd_sc_hd__nor2_8
XFILLER_228_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_31_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20672_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09665_ _19846_/Q _19660_/Q _20019_/Q vssd1 vssd1 vccd1 vccd1 _09665_/X sky130_fd_sc_hd__or3b_4
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09596_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09596_/X sky130_fd_sc_hd__or2_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ _21019_/CLK _20825_/D vssd1 vssd1 vccd1 vccd1 _20825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20756_ _20757_/CLK _20756_/D vssd1 vssd1 vccd1 vccd1 _20756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20687_ _20687_/CLK _20687_/D vssd1 vssd1 vccd1 vccd1 _20687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10440_ _19278_/Q _12044_/B _11684_/A1 vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__a21o_1
XFILLER_137_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371_ _11228_/A1 _09664_/B _10370_/X _11242_/B1 _19842_/Q vssd1 vssd1 vccd1 vccd1
+ _10371_/X sky130_fd_sc_hd__o32a_1
XFILLER_137_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12110_ _12110_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12111_/B sky130_fd_sc_hd__nand2_2
XFILLER_136_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13090_ _13007_/Y _13135_/A _13134_/B vssd1 vssd1 vccd1 vccd1 _13091_/C sky130_fd_sc_hd__o21ai_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12041_ _20359_/Q _12041_/B vssd1 vssd1 vccd1 vccd1 _12041_/X sky130_fd_sc_hd__or2_1
Xfanout1703 _09508_/Y vssd1 vssd1 vccd1 vccd1 _11191_/A sky130_fd_sc_hd__buf_12
XFILLER_172_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1714 _09507_/Y vssd1 vssd1 vccd1 vccd1 _11537_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_133_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1725 _09504_/Y vssd1 vssd1 vccd1 vccd1 _12752_/A sky130_fd_sc_hd__clkbuf_16
Xfanout1736 _11423_/C1 vssd1 vssd1 vccd1 vccd1 _12123_/C1 sky130_fd_sc_hd__buf_6
XFILLER_278_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1747 _09502_/Y vssd1 vssd1 vccd1 vccd1 _12310_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1758 _11240_/S vssd1 vssd1 vccd1 vccd1 _11243_/S sky130_fd_sc_hd__buf_8
Xfanout760 _18769_/Y vssd1 vssd1 vccd1 vccd1 _18840_/B sky130_fd_sc_hd__buf_6
X_15800_ _21034_/Q _21002_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _15800_/X sky130_fd_sc_hd__mux2_1
Xfanout771 _18560_/A vssd1 vssd1 vccd1 vccd1 _18667_/B sky130_fd_sc_hd__clkbuf_8
Xfanout1769 _13275_/A1 vssd1 vssd1 vccd1 vccd1 _14306_/A1 sky130_fd_sc_hd__buf_2
Xfanout782 _18490_/A vssd1 vssd1 vccd1 vccd1 _14110_/A sky130_fd_sc_hd__buf_4
X_13992_ _19164_/Q _14043_/A2 _14034_/B1 _13991_/X _16129_/B1 vssd1 vssd1 vccd1 vccd1
+ _19164_/D sky130_fd_sc_hd__o221a_1
X_16780_ _16780_/A vssd1 vssd1 vccd1 vccd1 _16780_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout793 _12488_/X vssd1 vssd1 vccd1 vccd1 _13350_/A sky130_fd_sc_hd__buf_8
XFILLER_120_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12943_ _14899_/B _14915_/B vssd1 vssd1 vccd1 vccd1 _16720_/B sky130_fd_sc_hd__or2_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15731_ _12828_/A _15978_/A2 _13428_/C _16063_/B2 vssd1 vssd1 vccd1 vccd1 _15732_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_280_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _18746_/A _18450_/B vssd1 vssd1 vccd1 vccd1 _20879_/D sky130_fd_sc_hd__and2_1
X_15662_ _20739_/Q _16011_/A2 _16011_/B1 _20771_/Q vssd1 vssd1 vccd1 vccd1 _15662_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 _16239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ _12483_/Y _12873_/X _15849_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12874_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_131 _13674_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _20249_/Q _17401_/A2 _17400_/X _17536_/D vssd1 vssd1 vccd1 vccd1 _20249_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_142 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _19377_/Q split4/X _14628_/S vssd1 vssd1 vccd1 vccd1 _19377_/D sky130_fd_sc_hd__mux2_1
X_11825_ _11823_/X _11824_/X _11904_/S vssd1 vssd1 vccd1 vccd1 _11825_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_153 _13770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18381_ _18550_/B _18385_/B vssd1 vssd1 vccd1 vccd1 _18381_/Y sky130_fd_sc_hd__nand2_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593_ _15593_/A _16009_/B vssd1 vssd1 vccd1 vccd1 _15593_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_164 _14522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _19111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_197 _19556_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17332_ _17402_/A _13844_/B _17231_/A _20217_/Q vssd1 vssd1 vccd1 vccd1 _17334_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _19314_/Q _17096_/A1 _14558_/S vssd1 vssd1 vccd1 vccd1 _19314_/D sky130_fd_sc_hd__mux2_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _10367_/Y _11796_/B _11415_/B vssd1 vssd1 vccd1 vccd1 _11757_/B sky130_fd_sc_hd__o21a_1
XFILLER_230_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10707_ _12427_/A1 _20125_/Q _20093_/Q _12417_/S vssd1 vssd1 vccd1 vccd1 _10707_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17263_ _17263_/A _17275_/B _17269_/C vssd1 vssd1 vccd1 vccd1 _17263_/X sky130_fd_sc_hd__and3_1
XFILLER_201_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14475_ _20233_/Q _19262_/Q _14477_/S vssd1 vssd1 vccd1 vccd1 _14476_/B sky130_fd_sc_hd__mux2_1
X_11687_ _12039_/A1 _10465_/B split7/A vssd1 vssd1 vccd1 vccd1 _11687_/X sky130_fd_sc_hd__a21o_4
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19002_ _18200_/Y _18983_/B _19002_/B1 _19001_/X vssd1 vssd1 vccd1 vccd1 _21020_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_220_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16214_ _19637_/Q _17900_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19637_/D sky130_fd_sc_hd__mux2_1
X_13426_ _13426_/A _13426_/B _13426_/C _15494_/A vssd1 vssd1 vccd1 vccd1 _13427_/D
+ sky130_fd_sc_hd__or4_1
X_17194_ _20158_/Q _17788_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20158_/D sky130_fd_sc_hd__mux2_1
X_10638_ _10642_/B _10638_/B vssd1 vssd1 vccd1 vccd1 _13596_/A sky130_fd_sc_hd__xor2_4
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16145_ _19596_/Q _16194_/S _16144_/Y _16195_/A vssd1 vssd1 vccd1 vccd1 _19596_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13357_ _13352_/X _13356_/X _14306_/A1 vssd1 vssd1 vccd1 vccd1 _13357_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10569_ _10057_/S _20095_/Q _11994_/S _10568_/X vssd1 vssd1 vccd1 vccd1 _10569_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12308_ _20396_/Q _20460_/Q _12389_/S vssd1 vssd1 vccd1 vccd1 _12308_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16076_ _19562_/Q _16079_/B _16075_/Y _16097_/B1 vssd1 vssd1 vccd1 vccd1 _19562_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_170_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13288_ _20927_/Q _13602_/A1 _13575_/C _13287_/Y _18612_/B vssd1 vssd1 vccd1 vccd1
+ _13288_/X sky130_fd_sc_hd__a221o_1
XFILLER_142_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19904_ _20467_/CLK _19904_/D vssd1 vssd1 vccd1 vccd1 _19904_/Q sky130_fd_sc_hd__dfxtp_1
X_15027_ _14896_/X _15283_/A _15096_/B vssd1 vssd1 vccd1 vccd1 _15028_/B sky130_fd_sc_hd__a21oi_1
X_12239_ _20051_/Q _19926_/Q _12316_/S vssd1 vssd1 vccd1 vccd1 _12239_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19835_ _20014_/CLK _19835_/D vssd1 vssd1 vccd1 vccd1 _19835_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19766_ _20704_/CLK _19766_/D vssd1 vssd1 vccd1 vccd1 _19766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16978_ _19988_/Q _17012_/A2 _16977_/Y _17012_/C1 vssd1 vssd1 vccd1 vccd1 _19988_/D
+ sky130_fd_sc_hd__a211o_1
Xinput4 coreIndex[3] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_6
XFILLER_237_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18717_ _20959_/Q _18225_/Y _18719_/S vssd1 vssd1 vccd1 vccd1 _18718_/B sky130_fd_sc_hd__mux2_1
X_15929_ _12034_/Y _12468_/X _15928_/X vssd1 vssd1 vccd1 vccd1 _15929_/X sky130_fd_sc_hd__o21a_1
X_19697_ _19697_/CLK _19697_/D vssd1 vssd1 vccd1 vccd1 _19697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18648_ _18529_/X _18684_/A2 _18646_/Y _18647_/Y vssd1 vssd1 vccd1 vccd1 _18649_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18579_ _18577_/Y _18578_/X _18598_/A vssd1 vssd1 vccd1 vccd1 _20917_/D sky130_fd_sc_hd__a21oi_1
XFILLER_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20610_ _20646_/CLK _20610_/D vssd1 vssd1 vccd1 vccd1 _20610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20541_ _20641_/CLK _20541_/D vssd1 vssd1 vccd1 vccd1 _20541_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20472_ _20472_/CLK _20472_/D vssd1 vssd1 vccd1 vccd1 _20472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput330 _13569_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[7] sky130_fd_sc_hd__buf_4
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput341 _13706_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[16] sky130_fd_sc_hd__buf_4
Xoutput352 _13755_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[26] sky130_fd_sc_hd__buf_4
XFILLER_273_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput363 _13663_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[7] sky130_fd_sc_hd__buf_4
Xoutput374 _13462_/X vssd1 vssd1 vccd1 vccd1 csb1[0] sky130_fd_sc_hd__buf_4
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput385 _13809_/X vssd1 vssd1 vccd1 vccd1 din0[18] sky130_fd_sc_hd__buf_4
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput396 _13819_/X vssd1 vssd1 vccd1 vccd1 din0[28] sky130_fd_sc_hd__buf_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21024_ _21024_/CLK _21024_/D vssd1 vssd1 vccd1 vccd1 _21024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09717_ _19821_/Q _19325_/Q _11915_/S vssd1 vssd1 vccd1 vccd1 _09717_/X sky130_fd_sc_hd__mux2_1
XFILLER_216_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09648_ _19660_/Q _20019_/Q vssd1 vssd1 vccd1 vccd1 _09648_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09579_ _19111_/Q _19110_/Q vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__or2_2
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _12039_/A1 _10377_/B _10037_/B vssd1 vssd1 vccd1 vccd1 _11610_/X sky130_fd_sc_hd__a21o_4
XFILLER_169_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20808_ _21029_/CLK _20808_/D vssd1 vssd1 vccd1 vccd1 _20808_/Q sky130_fd_sc_hd__dfxtp_1
X_12590_ _13657_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _12590_/Y sky130_fd_sc_hd__nor2_2
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11541_ _20477_/Q _11563_/S _11616_/B _11539_/X _11540_/X vssd1 vssd1 vccd1 vccd1
+ _11541_/X sky130_fd_sc_hd__a311o_1
XFILLER_51_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20739_ _20862_/CLK _20739_/D vssd1 vssd1 vccd1 vccd1 _20739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ _14260_/A _14260_/B _14260_/C vssd1 vssd1 vccd1 vccd1 _14262_/B sky130_fd_sc_hd__and3_1
XFILLER_167_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11472_ _19815_/Q _19319_/Q _12182_/S vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ _19241_/Q _19240_/Q _13231_/B _19242_/Q vssd1 vssd1 vccd1 vccd1 _13212_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10423_ _12060_/A1 _19345_/Q _20700_/Q _10426_/S _12051_/C1 vssd1 vssd1 vccd1 vccd1
+ _10423_/X sky130_fd_sc_hd__a221o_1
X_14191_ _14191_/A _14191_/B vssd1 vssd1 vccd1 vccd1 _14191_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ _13141_/X _13242_/B _13242_/A _13245_/A vssd1 vssd1 vccd1 vccd1 _13142_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_100_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10354_ _10409_/A _10354_/B vssd1 vssd1 vccd1 vccd1 _10354_/X sky130_fd_sc_hd__or2_1
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17950_ _20719_/Q _17950_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20719_/D sky130_fd_sc_hd__mux2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _13035_/Y _13383_/A _13382_/B vssd1 vssd1 vccd1 vccd1 _13073_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_279_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10285_ _10285_/A _10465_/A vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1500 _12041_/B vssd1 vssd1 vccd1 vccd1 _10897_/A3 sky130_fd_sc_hd__buf_2
X_16901_ input52/X input88/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16901_/X sky130_fd_sc_hd__mux2_8
X_12024_ _12102_/A1 _19361_/Q _20716_/Q _12025_/S _12100_/B1 vssd1 vssd1 vccd1 vccd1
+ _12024_/X sky130_fd_sc_hd__a221o_1
XFILLER_250_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1511 _11965_/B vssd1 vssd1 vccd1 vccd1 _11915_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17881_ _20654_/Q _17881_/A1 _17883_/S vssd1 vssd1 vccd1 vccd1 _20654_/D sky130_fd_sc_hd__mux2_1
Xfanout1522 fanout1534/X vssd1 vssd1 vccd1 vccd1 fanout1522/X sky130_fd_sc_hd__buf_4
Xfanout1533 fanout1534/X vssd1 vssd1 vccd1 vccd1 _12064_/S sky130_fd_sc_hd__buf_4
XFILLER_265_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19620_ _19620_/CLK _19620_/D vssd1 vssd1 vccd1 vccd1 _19620_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1544 _11174_/S vssd1 vssd1 vccd1 vccd1 _10924_/S sky130_fd_sc_hd__buf_6
Xfanout1555 fanout1556/X vssd1 vssd1 vccd1 vccd1 _11090_/S sky130_fd_sc_hd__clkbuf_4
X_16832_ _19971_/Q _16849_/A _16831_/Y _16896_/C1 vssd1 vssd1 vccd1 vccd1 _19971_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1566 _09627_/Y vssd1 vssd1 vccd1 vccd1 fanout1566/X sky130_fd_sc_hd__buf_6
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1577 _11597_/C1 vssd1 vssd1 vccd1 vccd1 _11684_/A1 sky130_fd_sc_hd__buf_6
XFILLER_93_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout590 _14738_/Y vssd1 vssd1 vccd1 vccd1 _14774_/A2 sky130_fd_sc_hd__buf_4
Xfanout1588 _11600_/C1 vssd1 vssd1 vccd1 vccd1 _11680_/C1 sky130_fd_sc_hd__buf_6
XFILLER_219_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19551_ _20425_/CLK _19551_/D vssd1 vssd1 vccd1 vccd1 _19551_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1599 _09901_/S vssd1 vssd1 vccd1 vccd1 _12150_/S sky130_fd_sc_hd__buf_6
X_16763_ _19964_/Q _16849_/A _16762_/Y _16451_/A vssd1 vssd1 vccd1 vccd1 _19964_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13975_ _14002_/A1 _13978_/A2 _10545_/X _14002_/B1 _19840_/Q vssd1 vssd1 vccd1 vccd1
+ _14063_/C sky130_fd_sc_hd__o32a_1
XFILLER_81_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18502_ _18612_/B _18502_/B vssd1 vssd1 vccd1 vccd1 _18502_/X sky130_fd_sc_hd__or2_2
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15714_ _19721_/Q _15961_/A2 _15961_/B1 _19753_/Q vssd1 vssd1 vccd1 vccd1 _15714_/X
+ sky130_fd_sc_hd__a22o_1
X_12926_ _20021_/Q _20020_/Q vssd1 vssd1 vccd1 vccd1 _12927_/B sky130_fd_sc_hd__nand2_2
X_19482_ _20712_/CLK _19482_/D vssd1 vssd1 vccd1 vccd1 _19482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16694_ _19949_/Q _17872_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19949_/D sky130_fd_sc_hd__mux2_1
XFILLER_234_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18433_ _20871_/Q _18265_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18434_/B sky130_fd_sc_hd__mux2_1
XFILLER_261_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15645_ _16002_/A1 _15630_/X _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15645_/X sky130_fd_sc_hd__a21o_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12857_ _19510_/Q _12857_/B vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__or2_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _20357_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__or2_1
XFILLER_61_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18364_ _20837_/Q _18363_/B _18363_/Y _18730_/A vssd1 vssd1 vccd1 vccd1 _20837_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15576_ _16052_/A1 _15562_/X _15575_/Y _13426_/B _16052_/B2 vssd1 vssd1 vccd1 vccd1
+ _15576_/X sky130_fd_sc_hd__a32o_1
X_12788_ _12785_/Y _12786_/X _19179_/Q _12652_/B vssd1 vssd1 vccd1 vccd1 _12790_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _20210_/Q _17321_/A2 _17305_/C _17314_/X _17330_/C1 vssd1 vssd1 vccd1 vccd1
+ _17315_/X sky130_fd_sc_hd__a221o_1
XFILLER_203_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14527_ _19301_/Q _14527_/A2 _14111_/B _17952_/A _14112_/C vssd1 vssd1 vccd1 vccd1
+ _19301_/D sky130_fd_sc_hd__a311oi_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ _13418_/A _11733_/Y _11737_/Y _11738_/X vssd1 vssd1 vccd1 vccd1 _11795_/B
+ sky130_fd_sc_hd__o211a_2
X_18295_ _18547_/B vssd1 vssd1 vccd1 vccd1 _18295_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17246_ _20187_/Q _17235_/Y _17279_/C1 vssd1 vssd1 vccd1 vccd1 _17246_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14458_ _14458_/A _14458_/B vssd1 vssd1 vccd1 vccd1 _19253_/D sky130_fd_sc_hd__and2_1
XFILLER_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13409_ _13405_/X _13408_/X _14295_/C1 vssd1 vssd1 vccd1 vccd1 _13409_/X sky130_fd_sc_hd__a21o_1
X_17177_ _20143_/Q _17805_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20143_/D sky130_fd_sc_hd__mux2_1
X_14389_ _14437_/A _14397_/B _14389_/C vssd1 vssd1 vccd1 vccd1 _14389_/X sky130_fd_sc_hd__or3_1
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16128_ _10122_/X _16132_/A2 _16127_/X vssd1 vssd1 vccd1 vccd1 _19588_/D sky130_fd_sc_hd__o21a_1
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16059_ _15983_/A _14877_/B _16057_/X _16058_/X _16054_/Y vssd1 vssd1 vccd1 vccd1
+ _16059_/X sky130_fd_sc_hd__a221o_1
XFILLER_97_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19818_ _20677_/CLK _19818_/D vssd1 vssd1 vccd1 vccd1 _19818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19749_ _20862_/CLK _19749_/D vssd1 vssd1 vccd1 vccd1 _19749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09502_ _09502_/A vssd1 vssd1 vccd1 vccd1 _09502_/Y sky130_fd_sc_hd__inv_6
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_20 _15600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 _15861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 _16840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20524_ _20688_/CLK _20524_/D vssd1 vssd1 vccd1 vccd1 _20524_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_53 _16961_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_64 _18225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_75 _09618_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_86 _11532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_97 _12402_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20455_ _20583_/CLK _20455_/D vssd1 vssd1 vccd1 vccd1 _20455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20386_ _20714_/CLK _20386_/D vssd1 vssd1 vccd1 vccd1 _20386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10070_ _12060_/A1 _19909_/Q _12070_/S _20034_/Q vssd1 vssd1 vccd1 vccd1 _10070_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21007_ _21011_/CLK _21007_/D vssd1 vssd1 vccd1 vccd1 _21007_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13760_ _13765_/A _13760_/B vssd1 vssd1 vccd1 vccd1 _13760_/X sky130_fd_sc_hd__and2_2
XFILLER_244_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10972_ _10373_/A _10377_/Y _09659_/B vssd1 vssd1 vccd1 vccd1 _10972_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12711_ _12711_/A _12716_/B vssd1 vssd1 vccd1 vccd1 _12711_/Y sky130_fd_sc_hd__nand2_1
X_13691_ _13692_/B vssd1 vssd1 vccd1 vccd1 _13691_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ _12640_/X _12641_/Y _12752_/B vssd1 vssd1 vccd1 vccd1 _12642_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15430_ _12578_/B _12782_/X _15429_/X _15589_/S vssd1 vssd1 vccd1 vccd1 _15430_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15361_ _10720_/A _15500_/A0 _15360_/X _10720_/B vssd1 vssd1 vccd1 vccd1 _15365_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_157_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12573_ _19156_/Q _11268_/C _12572_/Y vssd1 vssd1 vccd1 vccd1 _12580_/B sky130_fd_sc_hd__a21o_2
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17100_ _20070_/Q _17202_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20070_/D sky130_fd_sc_hd__mux2_1
X_11524_ _19814_/Q _19318_/Q _11527_/S vssd1 vssd1 vccd1 vccd1 _11524_/X sky130_fd_sc_hd__mux2_1
X_14312_ _19513_/Q _14312_/B vssd1 vssd1 vccd1 vccd1 _14314_/B sky130_fd_sc_hd__xnor2_1
X_18080_ _18080_/A _18085_/C vssd1 vssd1 vccd1 vccd1 _18080_/Y sky130_fd_sc_hd__nor2_1
X_15292_ _15110_/X _15113_/X _15292_/S vssd1 vssd1 vccd1 vccd1 _15292_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17031_ _20009_/Q input195/X _17040_/S vssd1 vssd1 vccd1 vccd1 _20009_/D sky130_fd_sc_hd__mux2_1
X_14243_ _14262_/A _14239_/B _14242_/X vssd1 vssd1 vccd1 vccd1 _14243_/X sky130_fd_sc_hd__a21bo_1
XFILLER_171_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11455_ _12157_/A1 _11454_/X _11451_/X _12153_/B1 vssd1 vssd1 vccd1 vccd1 _13707_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10406_ _19377_/Q _10603_/B _10404_/X _12085_/B2 _10405_/X vssd1 vssd1 vccd1 vccd1
+ _10406_/X sky130_fd_sc_hd__o221a_1
X_14174_ _19220_/Q _14205_/A2 _14172_/X _14173_/X _18476_/A vssd1 vssd1 vccd1 vccd1
+ _19220_/D sky130_fd_sc_hd__o221a_1
X_11386_ _11391_/A _19310_/Q _11391_/C vssd1 vssd1 vccd1 vccd1 _11386_/X sky130_fd_sc_hd__or3_1
XFILLER_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13125_ _13139_/A _19243_/Q _13119_/X _13124_/X vssd1 vssd1 vccd1 vccd1 _13941_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10337_ _20475_/Q _11305_/B _12504_/B vssd1 vssd1 vccd1 vccd1 _10337_/X sky130_fd_sc_hd__a21o_1
X_18982_ _18985_/B _18982_/B vssd1 vssd1 vccd1 vccd1 _18982_/X sky130_fd_sc_hd__and2_2
XFILLER_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17933_ _20702_/Q _17933_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20702_/D sky130_fd_sc_hd__mux2_1
X_13056_ _20950_/Q _20884_/Q vssd1 vssd1 vccd1 vccd1 _13056_/Y sky130_fd_sc_hd__nor2_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _19381_/Q _11291_/A2 _10266_/X _15129_/A0 _10267_/X vssd1 vssd1 vccd1 vccd1
+ _10268_/X sky130_fd_sc_hd__o221a_1
XFILLER_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12007_ _12007_/A1 _20520_/Q _12185_/S _20552_/Q vssd1 vssd1 vccd1 vccd1 _12007_/X
+ sky130_fd_sc_hd__o22a_1
Xfanout1330 _12458_/X vssd1 vssd1 vccd1 vccd1 _16030_/D1 sky130_fd_sc_hd__buf_6
XFILLER_267_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1341 _09688_/Y vssd1 vssd1 vccd1 vccd1 _10502_/A2 sky130_fd_sc_hd__buf_6
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1352 _17038_/S vssd1 vssd1 vccd1 vccd1 _17040_/S sky130_fd_sc_hd__buf_6
XFILLER_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17864_ _20637_/Q _17898_/A1 _17878_/S vssd1 vssd1 vccd1 vccd1 _20637_/D sky130_fd_sc_hd__mux2_1
X_10199_ _19542_/Q _09596_/A _11225_/B _19606_/Q _11246_/A1 vssd1 vssd1 vccd1 vccd1
+ _10199_/X sky130_fd_sc_hd__a221o_1
Xfanout1363 _17290_/B vssd1 vssd1 vccd1 vccd1 _17275_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_238_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_159_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21029_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_266_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19603_ _19603_/CLK _19603_/D vssd1 vssd1 vccd1 vccd1 _19603_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1374 _11693_/B vssd1 vssd1 vccd1 vccd1 _11708_/B sky130_fd_sc_hd__buf_6
X_16815_ _16878_/A _16815_/B vssd1 vssd1 vccd1 vccd1 _16815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1385 _11642_/S0 vssd1 vssd1 vccd1 vccd1 _11932_/S0 sky130_fd_sc_hd__buf_6
Xfanout1396 _11698_/B2 vssd1 vssd1 vccd1 vccd1 _10622_/S sky130_fd_sc_hd__buf_6
X_17795_ _20572_/Q _17935_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20572_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19534_ _19603_/CLK _19534_/D vssd1 vssd1 vccd1 vccd1 _19534_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_59_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16746_ _20182_/Q _17219_/B _16717_/X vssd1 vssd1 vccd1 vccd1 _16746_/X sky130_fd_sc_hd__a21o_1
XFILLER_35_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13958_ _19185_/Q _14051_/C _14003_/S vssd1 vssd1 vccd1 vccd1 _13958_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19465_ _20565_/CLK _19465_/D vssd1 vssd1 vccd1 vccd1 _19465_/Q sky130_fd_sc_hd__dfxtp_1
X_12909_ _13116_/A _13116_/B _13116_/C vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__a21o_1
XFILLER_262_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16677_ _19932_/Q _17855_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19932_/D sky130_fd_sc_hd__mux2_1
X_13889_ _19107_/Q _14738_/B _13889_/B1 _12513_/D _16189_/A vssd1 vssd1 vccd1 vccd1
+ _19107_/D sky130_fd_sc_hd__o221a_1
XFILLER_261_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18416_ _18416_/A _18416_/B vssd1 vssd1 vccd1 vccd1 _20862_/D sky130_fd_sc_hd__and2_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _11575_/A _12468_/X _15610_/Y _16053_/A _15627_/Y vssd1 vssd1 vccd1 vccd1
+ _15628_/X sky130_fd_sc_hd__o221a_1
X_19396_ _20687_/CLK _19396_/D vssd1 vssd1 vccd1 vccd1 _19396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18347_ _18499_/B _18349_/B vssd1 vssd1 vccd1 vccd1 _18347_/Y sky130_fd_sc_hd__nand2_1
X_15559_ _12464_/A _16063_/A2 _15591_/A vssd1 vssd1 vccd1 vccd1 _15559_/X sky130_fd_sc_hd__a21bo_1
XFILLER_159_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18278_ _19551_/Q _18308_/B vssd1 vssd1 vccd1 vccd1 _18278_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_257_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17229_ _17441_/A _17423_/D _17441_/C vssd1 vssd1 vccd1 vccd1 _17235_/B sky130_fd_sc_hd__and3_4
Xinput40 core_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_4
XFILLER_162_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput51 dout0[17] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput62 dout0[27] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_2
Xinput73 dout0[37] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_2
Xinput84 dout0[47] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_2
X_20240_ _21010_/CLK _20240_/D vssd1 vssd1 vccd1 vccd1 _20240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput95 dout0[57] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20171_ _20482_/CLK _20171_/D vssd1 vssd1 vccd1 vccd1 _20171_/Q sky130_fd_sc_hd__dfxtp_1
X_09982_ _12157_/A1 _17872_/A1 _09981_/X _12153_/B1 vssd1 vssd1 vccd1 vccd1 _13722_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_116_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20507_ _20539_/CLK _20507_/D vssd1 vssd1 vccd1 vccd1 _20507_/Q sky130_fd_sc_hd__dfxtp_1
X_11240_ _19559_/Q _11239_/X _11240_/S vssd1 vssd1 vccd1 vccd1 _11240_/X sky130_fd_sc_hd__mux2_1
X_20438_ _20438_/CLK _20438_/D vssd1 vssd1 vccd1 vccd1 _20438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11171_ _11258_/A1 _20119_/Q _20087_/Q _10924_/S vssd1 vssd1 vccd1 vccd1 _11171_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_268_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20369_ _20465_/CLK _20369_/D vssd1 vssd1 vccd1 vccd1 _20369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10122_ _11228_/A1 _14041_/A2 _10121_/X _11242_/B1 _19860_/Q vssd1 vssd1 vccd1 vccd1
+ _10122_/X sky130_fd_sc_hd__o32a_1
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14930_ _14119_/B _13192_/A _18148_/S vssd1 vssd1 vccd1 vccd1 _14930_/X sky130_fd_sc_hd__mux2_4
X_10053_ _20377_/Q _20441_/Q _10428_/S vssd1 vssd1 vccd1 vccd1 _10053_/X sky130_fd_sc_hd__mux2_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ _11322_/B _12114_/B _14870_/S vssd1 vssd1 vccd1 vccd1 _14862_/A sky130_fd_sc_hd__mux2_2
XFILLER_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16600_ _19863_/Q _16597_/X _16599_/Y vssd1 vssd1 vccd1 vccd1 _19863_/D sky130_fd_sc_hd__o21a_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _13816_/A1 _13729_/B _13816_/B1 input228/X vssd1 vssd1 vccd1 vccd1 _13812_/X
+ sky130_fd_sc_hd__a22o_1
X_17580_ _20338_/Q _17857_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20338_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14792_ _19143_/Q _14798_/A2 _14791_/X _14794_/C1 vssd1 vssd1 vccd1 vccd1 _19520_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_235_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16531_ _16557_/A _16531_/B vssd1 vssd1 vccd1 vccd1 _19831_/D sky130_fd_sc_hd__or2_1
XFILLER_44_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10955_ _12347_/A1 _19338_/Q _20693_/Q _11377_/S _11212_/S vssd1 vssd1 vccd1 vccd1
+ _10955_/X sky130_fd_sc_hd__a221o_1
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13743_ _13665_/Y _13741_/B _13741_/Y _13666_/Y _13742_/X vssd1 vssd1 vccd1 vccd1
+ _13744_/B sky130_fd_sc_hd__o221a_4
XFILLER_250_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19250_ _21013_/CLK _19250_/D vssd1 vssd1 vccd1 vccd1 _19250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16462_ _19771_/Q _17857_/A1 _16471_/S vssd1 vssd1 vccd1 vccd1 _19771_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10886_ _15264_/A vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__inv_2
X_13674_ _16598_/C _13674_/B vssd1 vssd1 vccd1 vccd1 _13674_/Y sky130_fd_sc_hd__nor2_1
XFILLER_73_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18201_ _09482_/Y _18490_/B _18236_/S vssd1 vssd1 vccd1 vccd1 _18202_/B sky130_fd_sc_hd__mux2_1
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15413_ _15413_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _15413_/Y sky130_fd_sc_hd__nand2_1
X_19181_ _21044_/CLK _19181_/D vssd1 vssd1 vccd1 vccd1 _19181_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12625_ _12483_/Y _12624_/X _15988_/A _15527_/A vssd1 vssd1 vccd1 vccd1 _12625_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16393_ _19742_/Q _16394_/C _19743_/Q vssd1 vssd1 vccd1 vccd1 _16395_/B sky130_fd_sc_hd__a21oi_1
XFILLER_231_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18132_ _18457_/B _18320_/A vssd1 vssd1 vccd1 vccd1 _18563_/A sky130_fd_sc_hd__nand2b_1
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15344_ _19709_/Q _15343_/X _15454_/S vssd1 vssd1 vccd1 vccd1 _15344_/X sky130_fd_sc_hd__mux2_2
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12556_ _13479_/A _13478_/A _18472_/B vssd1 vssd1 vccd1 vccd1 _18462_/B sky130_fd_sc_hd__or3b_1
XFILLER_40_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ _19881_/Q _19782_/Q _11916_/S vssd1 vssd1 vccd1 vccd1 _11507_/X sky130_fd_sc_hd__mux2_1
X_18063_ _20761_/Q _18063_/B vssd1 vssd1 vccd1 vccd1 _18069_/C sky130_fd_sc_hd__and2_2
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15275_ _20855_/Q _15274_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15275_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12487_ split8/A _12847_/A2 _16005_/A1 vssd1 vssd1 vccd1 vccd1 _12487_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17014_ _17014_/A _17014_/B vssd1 vssd1 vccd1 vccd1 _17015_/C sky130_fd_sc_hd__nand2_1
X_11438_ _20642_/Q _20606_/Q _12146_/S vssd1 vssd1 vccd1 vccd1 _11438_/X sky130_fd_sc_hd__mux2_1
X_14226_ _14219_/B _14221_/B _14219_/A vssd1 vssd1 vccd1 vccd1 _14232_/A sky130_fd_sc_hd__a21bo_1
X_14157_ _19498_/Q _14158_/B vssd1 vssd1 vccd1 vccd1 _14157_/Y sky130_fd_sc_hd__nor2_1
X_11369_ _19406_/Q _20565_/Q _11377_/S vssd1 vssd1 vccd1 vccd1 _11369_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13108_ _12913_/X _13106_/Y _13107_/Y _13323_/C vssd1 vssd1 vccd1 vccd1 _13108_/X
+ sky130_fd_sc_hd__a31o_1
X_14088_ _19203_/Q _14104_/A2 _14087_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1 _19203_/D
+ sky130_fd_sc_hd__o211a_1
X_18965_ _18553_/X _18964_/B _18963_/X _18964_/Y vssd1 vssd1 vccd1 vccd1 _18966_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17916_ _20687_/Q _17916_/A1 _17916_/S vssd1 vssd1 vccd1 vccd1 _20687_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _20958_/Q _20892_/Q vssd1 vssd1 vccd1 vccd1 _13039_/Y sky130_fd_sc_hd__nor2_2
XFILLER_224_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18896_ _20999_/Q _18978_/B vssd1 vssd1 vccd1 vccd1 _18896_/Y sky130_fd_sc_hd__nand2_1
Xfanout1160 _09631_/X vssd1 vssd1 vccd1 vccd1 _12401_/A1 sky130_fd_sc_hd__buf_4
Xfanout1171 _16009_/B vssd1 vssd1 vccd1 vccd1 _15988_/B sky130_fd_sc_hd__buf_4
XFILLER_254_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17847_ _20622_/Q input248/X _17849_/S vssd1 vssd1 vccd1 vccd1 _20622_/D sky130_fd_sc_hd__mux2_1
Xfanout1182 _16005_/A1 vssd1 vssd1 vccd1 vccd1 _15948_/A1 sky130_fd_sc_hd__buf_4
XFILLER_239_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1193 _11368_/A1 vssd1 vssd1 vccd1 vccd1 _12403_/A1 sky130_fd_sc_hd__buf_4
XFILLER_282_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17778_ _17918_/B _17812_/A vssd1 vssd1 vccd1 vccd1 _17779_/C sky130_fd_sc_hd__nor2_1
XFILLER_214_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19517_ _20291_/CLK _19517_/D vssd1 vssd1 vccd1 vccd1 _19517_/Q sky130_fd_sc_hd__dfxtp_4
X_16729_ _13468_/B _16725_/X _16728_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16730_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_34_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19448_ _20081_/CLK _19448_/D vssd1 vssd1 vccd1 vccd1 _19448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19379_ _20670_/CLK _19379_/D vssd1 vssd1 vccd1 vccd1 _19379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20084_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20223_ _20818_/CLK _20223_/D vssd1 vssd1 vccd1 vccd1 _20223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20154_ _20561_/CLK _20154_/D vssd1 vssd1 vccd1 vccd1 _20154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09965_ _09963_/X _09964_/X _11904_/S vssd1 vssd1 vccd1 vccd1 _09965_/X sky130_fd_sc_hd__mux2_1
XFILLER_277_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20085_ _20085_/CLK _20085_/D vssd1 vssd1 vccd1 vccd1 _20085_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _19644_/Q _12149_/S _09873_/X _09901_/S vssd1 vssd1 vccd1 vccd1 _09896_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_505 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_516 input242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_527 _19495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_538 _13473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_549 _16774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20987_ _21019_/CLK _20987_/D vssd1 vssd1 vccd1 vccd1 _20987_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_129_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10740_ _20028_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10740_/X sky130_fd_sc_hd__or2_1
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10671_ _19630_/Q _19936_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12410_ _12411_/A _20523_/Q _11116_/S _20555_/Q vssd1 vssd1 vccd1 vccd1 _12410_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ _19237_/Q _13390_/B vssd1 vssd1 vccd1 vccd1 _13390_/X sky130_fd_sc_hd__or2_1
XFILLER_223_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12341_ _12335_/X _12340_/X _12415_/S vssd1 vssd1 vccd1 vccd1 _12342_/B sky130_fd_sc_hd__mux2_2
XFILLER_182_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15060_ _15158_/B _15059_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _15060_/X sky130_fd_sc_hd__mux2_1
X_12272_ _10692_/A _20394_/Q _20458_/Q _12272_/B2 vssd1 vssd1 vccd1 vccd1 _12272_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14011_ _14035_/A1 _14011_/A2 _09866_/X _14035_/B1 _19852_/Q vssd1 vssd1 vccd1 vccd1
+ _14087_/C sky130_fd_sc_hd__o32a_1
XFILLER_5_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11223_ _11223_/A _11223_/B vssd1 vssd1 vccd1 vccd1 _15075_/A sky130_fd_sc_hd__xnor2_4
XFILLER_5_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11154_ _12230_/A1 _19898_/Q _11358_/S _20023_/Q _11363_/A1 vssd1 vssd1 vccd1 vccd1
+ _11155_/C sky130_fd_sc_hd__o221a_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10105_ _19635_/Q _19941_/Q _19279_/Q _20066_/Q _10092_/S _12084_/C vssd1 vssd1 vccd1
+ vccd1 _10105_/X sky130_fd_sc_hd__mux4_1
X_18750_ _18754_/A _18750_/B vssd1 vssd1 vccd1 vccd1 _20975_/D sky130_fd_sc_hd__and2_1
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11085_ _20399_/Q _20335_/Q _11161_/S vssd1 vssd1 vccd1 vccd1 _11085_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15962_ _19730_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15962_/X sky130_fd_sc_hd__or2_1
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput230 localMemory_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_hd__buf_12
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput241 localMemory_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_hd__buf_12
X_17701_ _20485_/Q _17944_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20485_/D sky130_fd_sc_hd__mux2_1
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14913_ _18149_/S _12512_/B _14912_/X vssd1 vssd1 vccd1 vccd1 _14951_/B sky130_fd_sc_hd__a21o_1
XFILLER_208_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10036_ _09684_/A _10021_/Y _10284_/A vssd1 vssd1 vccd1 vccd1 _11230_/A sky130_fd_sc_hd__mux2_2
Xinput252 localMemory_wb_we_i vssd1 vssd1 vccd1 vccd1 input252/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput263 manufacturerID[9] vssd1 vssd1 vccd1 vccd1 _17266_/A sky130_fd_sc_hd__buf_2
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18681_ _18966_/A _18681_/B vssd1 vssd1 vccd1 vccd1 _20943_/D sky130_fd_sc_hd__nor2_1
Xinput274 partID[4] vssd1 vssd1 vccd1 vccd1 _17284_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _15893_/A _15893_/B _15893_/C vssd1 vssd1 vccd1 vccd1 _15893_/X sky130_fd_sc_hd__and3_1
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _20388_/Q _17666_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20388_/D sky130_fd_sc_hd__mux2_1
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14844_ _14842_/X _14843_/X _15058_/S vssd1 vssd1 vccd1 vccd1 _14844_/X sky130_fd_sc_hd__mux2_1
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17563_ _20323_/Q _17802_/A1 _17567_/S vssd1 vssd1 vccd1 vccd1 _20323_/D sky130_fd_sc_hd__mux2_1
X_14775_ _19512_/Q _14797_/B vssd1 vssd1 vccd1 vccd1 _14775_/X sky130_fd_sc_hd__or2_1
X_11987_ _19393_/Q _20684_/Q _11987_/S vssd1 vssd1 vccd1 vccd1 _11987_/X sky130_fd_sc_hd__mux2_1
X_19302_ _20379_/CLK _19302_/D vssd1 vssd1 vccd1 vccd1 _19302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16514_ _19821_/Q _17107_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19821_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13726_ _13726_/A _13742_/B vssd1 vssd1 vccd1 vccd1 _13767_/B sky130_fd_sc_hd__or2_4
X_10938_ _19802_/Q _11291_/A2 _10936_/X _11291_/B2 _10937_/X vssd1 vssd1 vccd1 vccd1
+ _10938_/X sky130_fd_sc_hd__o221a_1
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17494_ _20282_/Q _17494_/B vssd1 vssd1 vccd1 vccd1 _17494_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19233_ _19511_/CLK _19233_/D vssd1 vssd1 vccd1 vccd1 _19233_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_232_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16445_ _18835_/A _16450_/C vssd1 vssd1 vccd1 vccd1 _16445_/Y sky130_fd_sc_hd__nor2_1
X_10869_ _09731_/A _10867_/X _10868_/X vssd1 vssd1 vccd1 vccd1 _10869_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_220_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13657_ _13657_/A _13657_/B vssd1 vssd1 vccd1 vccd1 _13694_/C sky130_fd_sc_hd__or2_4
XFILLER_143_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19164_ _19704_/CLK _19164_/D vssd1 vssd1 vccd1 vccd1 _19164_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _19514_/Q _19513_/Q _12835_/A vssd1 vssd1 vccd1 vccd1 _12811_/A sky130_fd_sc_hd__and3_1
X_16376_ _19736_/Q _16378_/C _16375_/Y vssd1 vssd1 vccd1 vccd1 _19736_/D sky130_fd_sc_hd__o21a_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13588_ _20923_/Q _13602_/A1 _13575_/C _13587_/X _18604_/B vssd1 vssd1 vccd1 vccd1
+ _13588_/X sky130_fd_sc_hd__a221o_1
XFILLER_8_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18115_ _20780_/Q _18117_/C _18114_/Y vssd1 vssd1 vccd1 vccd1 _20780_/D sky130_fd_sc_hd__o21a_1
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15327_ _15246_/A _15324_/X _15325_/Y _15326_/X _15303_/Y vssd1 vssd1 vccd1 vccd1
+ _15327_/X sky130_fd_sc_hd__o311a_1
XFILLER_145_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19095_ _19620_/CLK _19095_/D vssd1 vssd1 vccd1 vccd1 _19095_/Q sky130_fd_sc_hd__dfxtp_4
X_12539_ _20877_/Q _12549_/B _12539_/C vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__and3_1
XFILLER_118_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18046_ _18048_/A _18046_/B _18047_/B vssd1 vssd1 vccd1 vccd1 _20754_/D sky130_fd_sc_hd__nor3_1
X_15258_ _15258_/A _15258_/B vssd1 vssd1 vccd1 vccd1 _15258_/X sky130_fd_sc_hd__or2_1
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14209_ _14209_/A _14209_/B vssd1 vssd1 vccd1 vccd1 _14211_/A sky130_fd_sc_hd__nand2_1
XFILLER_125_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ _19705_/Q _15475_/A2 _15475_/B1 _19737_/Q vssd1 vssd1 vccd1 vccd1 _15189_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_174_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21004_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19997_ _20624_/CLK _19997_/D vssd1 vssd1 vccd1 vccd1 _19997_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_103_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20818_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09750_ _09748_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09750_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18948_ _18975_/A _18948_/B vssd1 vssd1 vccd1 vccd1 _18948_/Y sky130_fd_sc_hd__nand2_1
XFILLER_274_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09681_ _10284_/A _09681_/B _09681_/C vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__and3_1
X_18879_ _18975_/A _18879_/B vssd1 vssd1 vccd1 vccd1 _18879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_251_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20910_ _21008_/CLK _20910_/D vssd1 vssd1 vccd1 vccd1 _20910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20841_ _20969_/CLK _20841_/D vssd1 vssd1 vccd1 vccd1 _20841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20772_ _20862_/CLK _20772_/D vssd1 vssd1 vccd1 vccd1 _20772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20206_ _20763_/CLK _20206_/D vssd1 vssd1 vccd1 vccd1 _20206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_277_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1907 _16167_/C1 vssd1 vssd1 vccd1 vccd1 _16171_/A sky130_fd_sc_hd__clkbuf_2
Xfanout920 _15934_/A2 vssd1 vssd1 vccd1 vccd1 _16011_/A2 sky130_fd_sc_hd__buf_6
Xfanout1918 _13887_/C1 vssd1 vssd1 vccd1 vccd1 _18726_/A sky130_fd_sc_hd__buf_6
Xfanout931 _15035_/S vssd1 vssd1 vccd1 vccd1 _15062_/S sky130_fd_sc_hd__buf_6
Xfanout1929 _09515_/Y vssd1 vssd1 vccd1 vccd1 _14070_/C1 sky130_fd_sc_hd__buf_4
X_20137_ _20708_/CLK _20137_/D vssd1 vssd1 vccd1 vccd1 _20137_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout942 _11137_/A vssd1 vssd1 vccd1 vccd1 _15254_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_38_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09948_ _20353_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _09948_/X sky130_fd_sc_hd__or2_1
XFILLER_219_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout953 _14121_/X vssd1 vssd1 vccd1 vccd1 _14417_/S sky130_fd_sc_hd__buf_6
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout964 _17895_/A1 vssd1 vssd1 vccd1 vccd1 _17861_/A1 sky130_fd_sc_hd__buf_4
XFILLER_246_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout975 _17691_/A1 vssd1 vssd1 vccd1 vccd1 _17900_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout986 _10128_/X vssd1 vssd1 vccd1 vccd1 _17097_/A1 sky130_fd_sc_hd__buf_2
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20068_ _20315_/CLK _20068_/D vssd1 vssd1 vccd1 vccd1 _20068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout997 _16862_/A2 vssd1 vssd1 vccd1 vccd1 _16996_/A2 sky130_fd_sc_hd__buf_4
X_09879_ _20386_/Q _20450_/Q _11527_/S vssd1 vssd1 vccd1 vccd1 _09879_/X sky130_fd_sc_hd__mux2_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _19391_/Q _20682_/Q _11915_/S vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _12483_/Y _12889_/X _15904_/A _15527_/A vssd1 vssd1 vccd1 vccd1 _12890_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_79_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_302 input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 input243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11826_/X _11840_/X _12153_/A1 vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__a21o_2
XANTENNA_324 _13555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 _19494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_346 _13663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_357 _12426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14560_ _19330_/Q _17705_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19330_/D sky130_fd_sc_hd__mux2_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11772_/A _11772_/B _13596_/A vssd1 vssd1 vccd1 vccd1 _11773_/B sky130_fd_sc_hd__or3b_1
XANTENNA_368 _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_379 _15649_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _10553_/B _10290_/Y _10722_/X _10284_/X vssd1 vssd1 vccd1 vccd1 _10723_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_186_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13511_ _13511_/A _13511_/B vssd1 vssd1 vccd1 vccd1 _13512_/B sky130_fd_sc_hd__nor2_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14491_ _19269_/Q _17679_/A1 _14519_/S vssd1 vssd1 vccd1 vccd1 _19269_/D sky130_fd_sc_hd__mux2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _19653_/Q _17114_/A1 _16230_/S vssd1 vssd1 vccd1 vccd1 _19653_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10654_ _10652_/X _10653_/X _12376_/S vssd1 vssd1 vccd1 vccd1 _10654_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13442_ _16241_/B _13412_/X _13430_/Y split3/A vssd1 vssd1 vccd1 vccd1 _13463_/B
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_186_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16161_ _19604_/Q _16164_/B _16160_/Y _16165_/C1 vssd1 vssd1 vccd1 vccd1 _19604_/D
+ sky130_fd_sc_hd__o211a_1
X_13373_ _13373_/A _13373_/B vssd1 vssd1 vccd1 vccd1 _13373_/Y sky130_fd_sc_hd__nand2_1
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10585_ _10583_/X _10584_/X _10585_/S vssd1 vssd1 vccd1 vccd1 _10585_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ _15111_/X _15110_/X _15292_/S vssd1 vssd1 vccd1 vccd1 _15112_/X sky130_fd_sc_hd__mux2_1
X_12324_ _12322_/X _12323_/X _12324_/S vssd1 vssd1 vccd1 vccd1 _12324_/X sky130_fd_sc_hd__mux2_1
X_16092_ _10371_/X _16126_/A2 _16091_/X vssd1 vssd1 vccd1 vccd1 _19570_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20712_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12255_ _19395_/Q _12255_/A2 _12253_/X _12412_/B2 _12254_/X vssd1 vssd1 vccd1 vccd1
+ _12255_/X sky130_fd_sc_hd__o221a_1
XFILLER_182_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19920_ _20077_/CLK _19920_/D vssd1 vssd1 vccd1 vccd1 _19920_/Q sky130_fd_sc_hd__dfxtp_1
X_15043_ _14814_/X _14850_/X _15062_/S vssd1 vssd1 vccd1 vccd1 _15043_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11206_ _10937_/A _19335_/Q _20690_/Q _11211_/S _09730_/A vssd1 vssd1 vccd1 vccd1
+ _11206_/X sky130_fd_sc_hd__a221o_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19851_ _20017_/CLK _19851_/D vssd1 vssd1 vccd1 vccd1 _19851_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12186_ _12184_/X _12185_/X _12186_/S vssd1 vssd1 vccd1 vccd1 _12186_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18802_ _19090_/Q _12589_/B _12592_/C _15303_/B vssd1 vssd1 vccd1 vccd1 _18803_/B
+ sky130_fd_sc_hd__a22o_1
X_11137_ _11137_/A _11138_/B vssd1 vssd1 vccd1 vccd1 _11140_/A sky130_fd_sc_hd__nor2_1
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19782_ _20677_/CLK _19782_/D vssd1 vssd1 vccd1 vccd1 _19782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16994_ _19990_/Q _17012_/A2 _16993_/Y _17998_/A vssd1 vssd1 vccd1 vccd1 _19990_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18733_ _20967_/Q _18265_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18734_/B sky130_fd_sc_hd__mux2_1
XFILLER_283_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11068_ _20559_/Q _12213_/B vssd1 vssd1 vccd1 vccd1 _11068_/X sky130_fd_sc_hd__or2_1
X_15945_ _16051_/A1 _15931_/Y _16051_/B1 vssd1 vssd1 vccd1 vccd1 _15945_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ _19539_/Q _09596_/A _09613_/B _19603_/Q _11246_/A1 vssd1 vssd1 vccd1 vccd1
+ _10019_/X sky130_fd_sc_hd__a221o_1
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18664_ _18541_/X _18688_/A2 _18662_/Y _18663_/Y vssd1 vssd1 vccd1 vccd1 _18665_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_236_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _20907_/Q _16043_/A2 _15994_/B1 _15875_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _15876_/X sky130_fd_sc_hd__a221o_1
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17615_ _20371_/Q _17649_/A1 _17623_/S vssd1 vssd1 vccd1 vccd1 _20371_/D sky130_fd_sc_hd__mux2_1
XFILLER_225_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14827_ _11320_/B _12035_/B _14837_/S vssd1 vssd1 vccd1 vccd1 _14827_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18595_ _20922_/Q _18619_/B vssd1 vssd1 vccd1 vccd1 _18595_/Y sky130_fd_sc_hd__nand2_1
XFILLER_252_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17546_ _20306_/Q _17857_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20306_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14758_ _19126_/Q _14774_/A2 _14757_/X _14758_/C1 vssd1 vssd1 vccd1 vccd1 _19503_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_211_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13709_ _13655_/A _13670_/Y _13708_/Y _13714_/S vssd1 vssd1 vccd1 vccd1 _13709_/X
+ sky130_fd_sc_hd__o211a_1
X_17477_ _17487_/A1 _17476_/Y _18048_/A vssd1 vssd1 vccd1 vccd1 _20273_/D sky130_fd_sc_hd__a21oi_1
X_14689_ _19448_/Q _17938_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19448_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19216_ _19219_/CLK _19216_/D vssd1 vssd1 vccd1 vccd1 _19216_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_177_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16428_ _19756_/Q _16428_/B vssd1 vssd1 vccd1 vccd1 _16434_/C sky130_fd_sc_hd__and2_2
XFILLER_177_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19147_ _20300_/CLK _19147_/D vssd1 vssd1 vccd1 vccd1 _19147_/Q sky130_fd_sc_hd__dfxtp_1
X_16359_ _19730_/Q _16362_/C _18835_/A vssd1 vssd1 vccd1 vccd1 _16359_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19078_ _20423_/Q vssd1 vssd1 vccd1 vccd1 _20423_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18029_ _20748_/Q _18030_/C _18028_/Y vssd1 vssd1 vccd1 vccd1 _20748_/D sky130_fd_sc_hd__o21a_1
XFILLER_133_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21040_ _21040_/CLK _21040_/D vssd1 vssd1 vccd1 vccd1 _21040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09802_ _19684_/Q _20172_/Q _10428_/S vssd1 vssd1 vccd1 vccd1 _09802_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09733_ _10866_/A _10979_/C vssd1 vssd1 vccd1 vccd1 _09733_/Y sky130_fd_sc_hd__nand2_8
XFILLER_189_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09664_ _09672_/A _09664_/B _09664_/C vssd1 vssd1 vccd1 vccd1 _09664_/X sky130_fd_sc_hd__or3_1
XFILLER_255_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09595_ _09596_/B vssd1 vssd1 vccd1 vccd1 _09595_/Y sky130_fd_sc_hd__inv_2
XFILLER_270_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20341_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20824_ _21018_/CLK _20824_/D vssd1 vssd1 vccd1 vccd1 _20824_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20755_ _20794_/CLK _20755_/D vssd1 vssd1 vccd1 vccd1 _20755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20686_ _20686_/CLK _20686_/D vssd1 vssd1 vccd1 vccd1 _20686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ input109/X input144/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10370_/X sky130_fd_sc_hd__mux2_8
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _12156_/A1 _12039_/X _12038_/X vssd1 vssd1 vccd1 vccd1 _12040_/X sky130_fd_sc_hd__a21o_2
XFILLER_49_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1704 _12016_/C1 vssd1 vssd1 vccd1 vccd1 _11946_/C1 sky130_fd_sc_hd__buf_6
Xfanout1715 _10525_/S vssd1 vssd1 vccd1 vccd1 _10260_/S sky130_fd_sc_hd__buf_12
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1726 _11273_/A1 vssd1 vssd1 vccd1 vccd1 _11266_/A1 sky130_fd_sc_hd__buf_6
XFILLER_78_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1737 _11423_/C1 vssd1 vssd1 vccd1 vccd1 _12051_/C1 sky130_fd_sc_hd__buf_8
XFILLER_238_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout750 _18458_/X vssd1 vssd1 vccd1 vccd1 fanout750/X sky130_fd_sc_hd__buf_4
XFILLER_277_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1748 _12046_/B1 vssd1 vssd1 vccd1 vccd1 _12129_/S sky130_fd_sc_hd__buf_8
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1759 _09495_/Y vssd1 vssd1 vccd1 vccd1 _11240_/S sky130_fd_sc_hd__buf_6
XFILLER_219_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout761 _18686_/B vssd1 vssd1 vccd1 vccd1 _18682_/B sky130_fd_sc_hd__buf_6
XFILLER_265_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout772 _18560_/A vssd1 vssd1 vccd1 vccd1 _18687_/B sky130_fd_sc_hd__buf_2
X_13991_ _19196_/Q _14073_/C _14039_/S vssd1 vssd1 vccd1 vccd1 _13991_/X sky130_fd_sc_hd__mux2_1
Xfanout783 _18490_/A vssd1 vssd1 vccd1 vccd1 _18570_/B sky130_fd_sc_hd__buf_8
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout794 _12652_/B vssd1 vssd1 vccd1 vccd1 split6/A sky130_fd_sc_hd__buf_8
XFILLER_74_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _15977_/A1 _12824_/X _15729_/X _16062_/B2 vssd1 vssd1 vccd1 vccd1 _15732_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_218_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12942_ _19259_/Q _12950_/B2 _12930_/X _20007_/Q vssd1 vssd1 vccd1 vccd1 _14912_/B
+ sky130_fd_sc_hd__a22o_2
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15661_ _19719_/Q _15933_/B vssd1 vssd1 vccd1 vccd1 _15661_/X sky130_fd_sc_hd__or2_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_110 _13507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ _12884_/B _12873_/B vssd1 vssd1 vccd1 vccd1 _12873_/X sky130_fd_sc_hd__or2_1
XFILLER_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_121 _13708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _20248_/Q _17337_/B _17530_/A2 _20297_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17400_/X sky130_fd_sc_hd__a221o_1
XANTENNA_132 _13683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _19376_/Q _17896_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19376_/D sky130_fd_sc_hd__mux2_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _11903_/A1 _11817_/X _11818_/X vssd1 vssd1 vccd1 vccd1 _11824_/X sky130_fd_sc_hd__o21a_1
X_18380_ _20845_/Q _18387_/B _18379_/Y _18730_/A vssd1 vssd1 vccd1 vccd1 _20845_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _19541_/Q _15591_/A _15591_/Y _16167_/C1 vssd1 vssd1 vccd1 vccd1 _19541_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_154 _13775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _14522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_176 _19114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _20216_/Q _17331_/A2 _17330_/X _17331_/C1 vssd1 vssd1 vccd1 vccd1 _20216_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_187 _19165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _19557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14543_ _19313_/Q _17095_/A1 _14558_/S vssd1 vssd1 vccd1 vccd1 _19313_/D sky130_fd_sc_hd__mux2_1
XFILLER_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11755_ _13424_/A _11754_/B _11413_/Y vssd1 vssd1 vccd1 vccd1 _11796_/B sky130_fd_sc_hd__a21boi_4
XFILLER_201_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17262_ _20193_/Q _17280_/A2 _17261_/X _17331_/C1 vssd1 vssd1 vccd1 vccd1 _20193_/D
+ sky130_fd_sc_hd__o211a_1
X_10706_ _19669_/Q _12417_/S _12419_/C1 vssd1 vssd1 vccd1 vccd1 _10706_/X sky130_fd_sc_hd__o21a_1
XFILLER_202_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14474_ _18985_/A _14474_/B vssd1 vssd1 vccd1 vccd1 _19261_/D sky130_fd_sc_hd__and2_1
XFILLER_230_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ _11671_/X _11685_/X _12074_/B1 vssd1 vssd1 vccd1 vccd1 _11686_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19001_ _21020_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _19001_/X sky130_fd_sc_hd__or2_1
X_16213_ _19636_/Q _17097_/A1 _16230_/S vssd1 vssd1 vccd1 vccd1 _19636_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13425_ _13425_/A _13425_/B vssd1 vssd1 vccd1 vccd1 _15494_/A sky130_fd_sc_hd__xnor2_4
X_17193_ _20157_/Q _17927_/A1 _17215_/S vssd1 vssd1 vccd1 vccd1 _20157_/D sky130_fd_sc_hd__mux2_1
X_10637_ _10642_/B _10638_/B vssd1 vssd1 vccd1 vccd1 _15410_/S sky130_fd_sc_hd__nor2_2
XFILLER_127_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16144_ _16774_/B _16196_/S vssd1 vssd1 vccd1 vccd1 _16144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10568_ _10057_/S _10581_/A1 _20127_/Q _12059_/A1 vssd1 vssd1 vccd1 vccd1 _10568_/X
+ sky130_fd_sc_hd__a31o_1
X_13356_ _13355_/B _13354_/Y _13355_/Y _18628_/B vssd1 vssd1 vccd1 vccd1 _13356_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12307_ _20492_/Q _20332_/Q _12389_/S vssd1 vssd1 vccd1 vccd1 _12307_/X sky130_fd_sc_hd__mux2_1
X_16075_ _16075_/A _16079_/B vssd1 vssd1 vccd1 vccd1 _16075_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10499_ _19633_/Q _09689_/D _10496_/X _10497_/X _10498_/X vssd1 vssd1 vccd1 vccd1
+ _10499_/X sky130_fd_sc_hd__o221a_1
X_13287_ _13287_/A _13378_/B vssd1 vssd1 vccd1 vccd1 _13287_/Y sky130_fd_sc_hd__nor2_1
X_19903_ _20061_/CLK _19903_/D vssd1 vssd1 vccd1 vccd1 _19903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _15026_/A _15095_/B vssd1 vssd1 vccd1 vccd1 _15026_/Y sky130_fd_sc_hd__nand2_4
X_12238_ _12317_/S _12237_/X _12236_/X _12318_/A1 vssd1 vssd1 vccd1 vccd1 _12238_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19834_ _20004_/CLK _19834_/D vssd1 vssd1 vccd1 vccd1 _19834_/Q sky130_fd_sc_hd__dfxtp_4
X_12169_ _20393_/Q _20457_/Q _12174_/S vssd1 vssd1 vccd1 vccd1 _12169_/X sky130_fd_sc_hd__mux2_1
XFILLER_268_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19765_ _19978_/CLK _19765_/D vssd1 vssd1 vccd1 vccd1 _19765_/Q sky130_fd_sc_hd__dfxtp_1
X_16977_ _16974_/Y _16976_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16977_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput5 coreIndex[4] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
XFILLER_49_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15928_ _14815_/S _15218_/B _15224_/Y _16053_/A _15927_/X vssd1 vssd1 vccd1 vccd1
+ _15928_/X sky130_fd_sc_hd__o221a_1
X_18716_ _18720_/A _18716_/B vssd1 vssd1 vccd1 vccd1 _20958_/D sky130_fd_sc_hd__and2_1
XFILLER_283_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19696_ _19696_/CLK _19696_/D vssd1 vssd1 vccd1 vccd1 _19696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18647_ _19515_/Q _18683_/B vssd1 vssd1 vccd1 vccd1 _18647_/Y sky130_fd_sc_hd__nand2_1
X_15859_ _20810_/Q _15941_/A2 _15852_/X _15941_/B2 _15858_/X vssd1 vssd1 vccd1 vccd1
+ _15859_/X sky130_fd_sc_hd__a221o_2
XFILLER_80_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18578_ _19497_/Q _18589_/B _18473_/A _18564_/A vssd1 vssd1 vccd1 vccd1 _18578_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_212_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17529_ _20300_/Q _20298_/Q _17528_/X vssd1 vssd1 vccd1 vccd1 _17529_/X sky130_fd_sc_hd__or3b_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20540_ _20672_/CLK _20540_/D vssd1 vssd1 vccd1 vccd1 _20540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20471_ _21047_/A _20471_/D vssd1 vssd1 vccd1 vccd1 _20471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput320 _13626_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[23] sky130_fd_sc_hd__buf_4
XFILLER_273_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput331 _13584_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[8] sky130_fd_sc_hd__buf_4
Xoutput342 _13711_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[17] sky130_fd_sc_hd__buf_4
Xoutput353 _13760_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[27] sky130_fd_sc_hd__buf_4
XFILLER_0_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput364 _13669_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[8] sky130_fd_sc_hd__buf_4
Xoutput375 _16278_/B vssd1 vssd1 vccd1 vccd1 csb1[1] sky130_fd_sc_hd__buf_4
XFILLER_160_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput386 _13810_/X vssd1 vssd1 vccd1 vccd1 din0[19] sky130_fd_sc_hd__buf_4
X_21023_ _21023_/CLK _21023_/D vssd1 vssd1 vccd1 vccd1 _21023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput397 _13820_/X vssd1 vssd1 vccd1 vccd1 din0[29] sky130_fd_sc_hd__buf_4
XFILLER_87_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09716_ _19646_/Q _11915_/S _09692_/X _11917_/S vssd1 vssd1 vccd1 vccd1 _09716_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09647_ input131/X input166/X _11241_/S vssd1 vssd1 vccd1 vccd1 _09647_/X sky130_fd_sc_hd__mux2_8
XFILLER_216_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09578_ _19098_/Q _10020_/B _09576_/X _19114_/Q vssd1 vssd1 vccd1 vccd1 _09578_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20807_ _21029_/CLK _20807_/D vssd1 vssd1 vccd1 vccd1 _20807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_169_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11540_ _20317_/Q _11563_/S _09928_/S _11945_/S vssd1 vssd1 vccd1 vccd1 _11540_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20738_ _20862_/CLK _20738_/D vssd1 vssd1 vccd1 vccd1 _20738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_206_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20673_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11471_ _12189_/A _11471_/B vssd1 vssd1 vccd1 vccd1 _11471_/X sky130_fd_sc_hd__or2_1
X_20669_ _20669_/CLK _20669_/D vssd1 vssd1 vccd1 vccd1 _20669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13210_ _13209_/B _13209_/C _13209_/A vssd1 vssd1 vccd1 vccd1 _13210_/X sky130_fd_sc_hd__a21o_1
X_10422_ _19409_/Q _20568_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _10422_/X sky130_fd_sc_hd__mux2_1
X_14190_ _14176_/Y _14181_/B _14178_/B vssd1 vssd1 vccd1 vccd1 _14191_/B sky130_fd_sc_hd__o21ai_4
XFILLER_136_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10353_ _10351_/X _10352_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _10354_/B sky130_fd_sc_hd__mux2_1
X_13141_ _13138_/X _13139_/X _16187_/A vssd1 vssd1 vccd1 vccd1 _13141_/X sky130_fd_sc_hd__o21a_2
XFILLER_164_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13072_ _13290_/A _13290_/C _13290_/B vssd1 vssd1 vccd1 vccd1 _13383_/A sky130_fd_sc_hd__a21boi_4
X_10284_ _10284_/A _11234_/B _10283_/X vssd1 vssd1 vccd1 vccd1 _10284_/X sky130_fd_sc_hd__or3b_2
XFILLER_183_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16900_ _16932_/A1 _16899_/X _16932_/B1 vssd1 vssd1 vccd1 vccd1 _16900_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12023_ _12021_/X _12022_/X _12023_/S vssd1 vssd1 vccd1 vccd1 _12023_/X sky130_fd_sc_hd__mux2_1
Xfanout1501 _12213_/B vssd1 vssd1 vccd1 vccd1 _12295_/B sky130_fd_sc_hd__buf_8
XFILLER_151_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17880_ _20653_/Q _17914_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20653_/D sky130_fd_sc_hd__mux2_1
Xfanout1512 _11599_/S vssd1 vssd1 vccd1 vccd1 _11965_/B sky130_fd_sc_hd__buf_6
XFILLER_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_250_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1523 _11665_/S vssd1 vssd1 vccd1 vccd1 _12053_/S sky130_fd_sc_hd__buf_6
XFILLER_278_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1534 fanout1566/X vssd1 vssd1 vccd1 vccd1 fanout1534/X sky130_fd_sc_hd__buf_6
XFILLER_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1545 _10316_/S vssd1 vssd1 vccd1 vccd1 _11174_/S sky130_fd_sc_hd__buf_4
X_16831_ _16849_/A _16831_/B vssd1 vssd1 vccd1 vccd1 _16831_/Y sky130_fd_sc_hd__nor2_1
Xfanout1556 fanout1566/X vssd1 vssd1 vccd1 vccd1 fanout1556/X sky130_fd_sc_hd__clkbuf_8
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1567 _09625_/Y vssd1 vssd1 vccd1 vccd1 _12144_/C1 sky130_fd_sc_hd__buf_8
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1578 _11597_/C1 vssd1 vssd1 vccd1 vccd1 _12072_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout580 _16199_/X vssd1 vssd1 vccd1 vccd1 _16228_/S sky130_fd_sc_hd__buf_12
XFILLER_281_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1589 _11600_/C1 vssd1 vssd1 vccd1 vccd1 _12068_/C1 sky130_fd_sc_hd__clkbuf_4
X_19550_ _20425_/CLK _19550_/D vssd1 vssd1 vccd1 vccd1 _19550_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout591 _14733_/S vssd1 vssd1 vccd1 vccd1 _14732_/S sky130_fd_sc_hd__buf_12
XFILLER_265_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16762_ _16758_/Y _16761_/X _17011_/B1 vssd1 vssd1 vccd1 vccd1 _16762_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13974_ _19158_/Q _13986_/A2 _14004_/B1 _13973_/X _16143_/A vssd1 vssd1 vccd1 vccd1
+ _19158_/D sky130_fd_sc_hd__o221a_1
XFILLER_253_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18501_ _18856_/A _18501_/B vssd1 vssd1 vccd1 vccd1 _20893_/D sky130_fd_sc_hd__nor2_1
XFILLER_207_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15713_ _15713_/A _16037_/B vssd1 vssd1 vccd1 vccd1 _15713_/Y sky130_fd_sc_hd__nor2_1
X_12925_ _20021_/Q _20020_/Q vssd1 vssd1 vccd1 vccd1 _17015_/B sky130_fd_sc_hd__or2_4
X_19481_ _20081_/CLK _19481_/D vssd1 vssd1 vccd1 vccd1 _19481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16693_ _19948_/Q _17939_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19948_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18432_ _18736_/A _18432_/B vssd1 vssd1 vccd1 vccd1 _20870_/D sky130_fd_sc_hd__and2_1
XFILLER_61_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15644_ _15644_/A1 _16878_/B _15630_/X vssd1 vssd1 vccd1 vccd1 _15644_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_234_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12856_ _11570_/Y _15527_/A _12484_/X _12855_/X vssd1 vssd1 vccd1 vccd1 _12856_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_33_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _12156_/A1 _11806_/X _11805_/X vssd1 vssd1 vccd1 vccd1 _11807_/X sky130_fd_sc_hd__a21o_4
X_18363_ _18523_/B _18363_/B vssd1 vssd1 vccd1 vccd1 _18363_/Y sky130_fd_sc_hd__nand2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _15644_/A1 _16860_/B _15561_/Y vssd1 vssd1 vccd1 vccd1 _15575_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_187_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12787_ _19179_/Q _12652_/B _12785_/Y _12786_/X vssd1 vssd1 vccd1 vccd1 _12790_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17314_ input3/X input269/X _17320_/S vssd1 vssd1 vccd1 vccd1 _17314_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14524_/X _14525_/X _16167_/C1 vssd1 vssd1 vccd1 vccd1 _19300_/D sky130_fd_sc_hd__o21a_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18294_ _18313_/B _14392_/B _18293_/Y vssd1 vssd1 vccd1 vccd1 _18547_/B sky130_fd_sc_hd__o21ai_4
X_11738_ _13418_/A _13419_/A _11736_/Y vssd1 vssd1 vccd1 vccd1 _11738_/X sky130_fd_sc_hd__or3b_1
XFILLER_202_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17245_ _17245_/A _17290_/B _17269_/C vssd1 vssd1 vccd1 vccd1 _17245_/X sky130_fd_sc_hd__and3_1
X_14457_ _20224_/Q _19253_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14458_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11669_ _10430_/S _11662_/X _11663_/X vssd1 vssd1 vccd1 vccd1 _11669_/X sky130_fd_sc_hd__o21a_1
X_13408_ _20961_/Q _13355_/B _13407_/Y _18767_/A vssd1 vssd1 vccd1 vccd1 _13408_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_259_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17176_ _20142_/Q _17804_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20142_/D sky130_fd_sc_hd__mux2_1
X_14388_ _13139_/A _14387_/X _13229_/X vssd1 vssd1 vccd1 vccd1 _14389_/C sky130_fd_sc_hd__a21o_1
XFILLER_127_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16127_ _19588_/Q _16127_/A2 _16127_/B1 vssd1 vssd1 vccd1 vccd1 _16127_/X sky130_fd_sc_hd__o21a_1
XFILLER_128_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13339_ _20963_/Q _20897_/Q vssd1 vssd1 vccd1 vccd1 _13340_/B sky130_fd_sc_hd__xor2_1
XFILLER_116_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16058_ _14882_/A _16058_/A2 _12467_/Y vssd1 vssd1 vccd1 vccd1 _16058_/X sky130_fd_sc_hd__a21o_1
XFILLER_170_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15009_ _14903_/Y _14936_/Y _15008_/Y vssd1 vssd1 vccd1 vccd1 _16708_/B sky130_fd_sc_hd__o21a_4
XFILLER_116_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19817_ _19956_/CLK _19817_/D vssd1 vssd1 vccd1 vccd1 _19817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19748_ _20863_/CLK _19748_/D vssd1 vssd1 vccd1 vccd1 _19748_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_238_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09501_ _10831_/S vssd1 vssd1 vccd1 vccd1 _09501_/Y sky130_fd_sc_hd__inv_12
XFILLER_271_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19679_ _20641_/CLK _19679_/D vssd1 vssd1 vccd1 vccd1 _19679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_10 _15419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _15600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 _15861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20523_ _20655_/CLK _20523_/D vssd1 vssd1 vccd1 vccd1 _20523_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_43 _16849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_54 _16969_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 _18225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_76 _09625_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_87 _11568_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20454_ _20481_/CLK _20454_/D vssd1 vssd1 vccd1 vccd1 _20454_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_98 _16009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20385_ _20481_/CLK _20385_/D vssd1 vssd1 vccd1 vccd1 _20385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21006_ _21006_/CLK _21006_/D vssd1 vssd1 vccd1 vccd1 _21006_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10971_ _19530_/Q _09613_/A _18152_/C _19594_/Q vssd1 vssd1 vccd1 vccd1 _10971_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12710_ _13350_/A _12710_/B vssd1 vssd1 vccd1 vccd1 _12839_/A sky130_fd_sc_hd__nand2_4
XFILLER_271_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13690_ _13735_/A _13688_/X _13689_/X _13659_/A vssd1 vssd1 vccd1 vccd1 _13692_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_253_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12641_ _15304_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _12641_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15360_ _10720_/A _12471_/X _12468_/X vssd1 vssd1 vccd1 vccd1 _15360_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12572_ _19155_/Q _19154_/Q vssd1 vssd1 vccd1 vccd1 _12572_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14311_ _19513_/Q _14312_/B vssd1 vssd1 vccd1 vccd1 _14323_/A sky130_fd_sc_hd__nand2_1
XFILLER_200_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11523_ _19639_/Q _11527_/S _11500_/X _11528_/S vssd1 vssd1 vccd1 vccd1 _11523_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15291_ _15106_/X _15111_/X _15292_/S vssd1 vssd1 vccd1 vccd1 _15291_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17030_ _20008_/Q input194/X _17040_/S vssd1 vssd1 vccd1 vccd1 _20008_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14242_ _14262_/A _14242_/B _14250_/B vssd1 vssd1 vccd1 vccd1 _14242_/X sky130_fd_sc_hd__or3b_1
X_11454_ _12156_/A1 _11452_/X _11453_/X vssd1 vssd1 vccd1 vccd1 _11454_/X sky130_fd_sc_hd__a21o_2
XFILLER_183_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10405_ _12084_/A _20668_/Q _10405_/C vssd1 vssd1 vccd1 vccd1 _10405_/X sky130_fd_sc_hd__or3_1
X_11385_ _11391_/A _19905_/Q _11393_/S0 _20030_/Q vssd1 vssd1 vccd1 vccd1 _11385_/X
+ sky130_fd_sc_hd__o22a_1
X_14173_ _14173_/A _14255_/A _16068_/B vssd1 vssd1 vccd1 vccd1 _14173_/X sky130_fd_sc_hd__or3_1
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ _13205_/A _13124_/B vssd1 vssd1 vccd1 vccd1 _13124_/X sky130_fd_sc_hd__and2_1
X_10336_ _10356_/A _20379_/Q _20443_/Q _11295_/S _09730_/A vssd1 vssd1 vccd1 vccd1
+ _10336_/X sky130_fd_sc_hd__a221o_1
X_18981_ _18981_/A _18981_/B _18981_/C vssd1 vssd1 vccd1 vccd1 _18981_/X sky130_fd_sc_hd__or3_4
XFILLER_113_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10267_ _11021_/A _20672_/Q _11021_/C vssd1 vssd1 vccd1 vccd1 _10267_/X sky130_fd_sc_hd__or3_1
X_13055_ _20951_/Q _20885_/Q vssd1 vssd1 vccd1 vccd1 _13055_/Y sky130_fd_sc_hd__nand2_1
X_17932_ _20701_/Q _17932_/A1 _17934_/S vssd1 vssd1 vccd1 vccd1 _20701_/D sky130_fd_sc_hd__mux2_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1320 _15500_/A0 vssd1 vssd1 vccd1 vccd1 _15984_/A2 sky130_fd_sc_hd__buf_6
XFILLER_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12006_ _12004_/X _12005_/X _12006_/S vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__mux2_1
Xfanout1331 _12085_/A2 vssd1 vssd1 vccd1 vccd1 _12009_/A2 sky130_fd_sc_hd__clkbuf_16
X_17863_ _20636_/Q split4/X _17878_/S vssd1 vssd1 vccd1 vccd1 _20636_/D sky130_fd_sc_hd__mux2_1
XFILLER_266_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1342 _17390_/A2 vssd1 vssd1 vccd1 vccd1 _17337_/B sky130_fd_sc_hd__buf_6
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10198_ _10198_/A _15549_/S vssd1 vssd1 vccd1 vccd1 _13424_/A sky130_fd_sc_hd__nand2_8
XFILLER_121_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1353 _17015_/Y vssd1 vssd1 vccd1 vccd1 _17038_/S sky130_fd_sc_hd__buf_6
Xfanout1364 _17320_/S vssd1 vssd1 vccd1 vccd1 _17290_/B sky130_fd_sc_hd__buf_2
XFILLER_239_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19602_ _19603_/CLK _19602_/D vssd1 vssd1 vccd1 vccd1 _19602_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1375 _11213_/B vssd1 vssd1 vccd1 vccd1 _11693_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_282_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16814_ _19969_/Q _16887_/A _16813_/Y _16896_/C1 vssd1 vssd1 vccd1 vccd1 _19969_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_93_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17794_ _20571_/Q _17934_/A1 _17794_/S vssd1 vssd1 vccd1 vccd1 _20571_/D sky130_fd_sc_hd__mux2_1
Xfanout1386 _11860_/B2 vssd1 vssd1 vccd1 vccd1 _11642_/S0 sky130_fd_sc_hd__buf_4
XFILLER_19_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1397 _11698_/B2 vssd1 vssd1 vccd1 vccd1 _10621_/S sky130_fd_sc_hd__buf_4
XFILLER_219_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16745_ _19217_/Q _16996_/A2 _16996_/B1 _19086_/Q _16744_/X vssd1 vssd1 vccd1 vccd1
+ _16745_/X sky130_fd_sc_hd__o221a_1
X_19533_ _19620_/CLK _19533_/D vssd1 vssd1 vccd1 vccd1 _19533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13957_ _14041_/A1 _13969_/A2 _10974_/X _14041_/B1 _19834_/Q vssd1 vssd1 vccd1 vccd1
+ _14051_/C sky130_fd_sc_hd__o32a_1
XFILLER_207_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_199_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20681_/CLK sky130_fd_sc_hd__clkbuf_16
X_19464_ _20563_/CLK _19464_/D vssd1 vssd1 vccd1 vccd1 _19464_/Q sky130_fd_sc_hd__dfxtp_1
X_12908_ _12908_/A vssd1 vssd1 vccd1 vccd1 _13116_/C sky130_fd_sc_hd__inv_2
X_16676_ _19931_/Q _17679_/A1 _16704_/S vssd1 vssd1 vccd1 vccd1 _19931_/D sky130_fd_sc_hd__mux2_1
XFILLER_207_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13888_ _19106_/Q _14527_/A2 _13896_/B1 _12584_/B _16193_/A vssd1 vssd1 vccd1 vccd1
+ _19106_/D sky130_fd_sc_hd__o221a_1
XFILLER_146_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_128_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21017_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18415_ _20862_/Q _18220_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18416_/B sky130_fd_sc_hd__mux2_1
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15627_ _11575_/B _16058_/A2 _15264_/B _13421_/A _16030_/D1 vssd1 vssd1 vccd1 vccd1
+ _15627_/Y sky130_fd_sc_hd__a221oi_1
X_19395_ _20663_/CLK _19395_/D vssd1 vssd1 vccd1 vccd1 _19395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12839_ _12839_/A _12839_/B _12839_/C _12839_/D vssd1 vssd1 vccd1 vccd1 _13300_/B
+ sky130_fd_sc_hd__or4_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18346_ _20828_/Q _18349_/B _18345_/Y _18985_/A vssd1 vssd1 vccd1 vccd1 _20828_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _13426_/C _15557_/X _15589_/S vssd1 vssd1 vccd1 vccd1 _15558_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14509_ _19287_/Q _17872_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19287_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18277_ _18724_/A _18277_/B vssd1 vssd1 vccd1 vccd1 _20809_/D sky130_fd_sc_hd__and2_1
X_15489_ _16052_/A1 _15474_/X _15487_/Y _15488_/Y vssd1 vssd1 vccd1 vccd1 _15489_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17228_ _20265_/Q _20264_/Q vssd1 vssd1 vccd1 vccd1 _17421_/B sky130_fd_sc_hd__or2_1
Xinput30 core_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_4
Xinput41 core_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
Xinput52 dout0[18] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput63 dout0[28] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
X_17159_ _20125_/Q _17927_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20125_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput74 dout0[38] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_2
Xinput85 dout0[48] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_2
Xinput96 dout0[58] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20170_ _20481_/CLK _20170_/D vssd1 vssd1 vccd1 vccd1 _20170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09981_ _09966_/X _09980_/X _12153_/A1 vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__a21o_2
XFILLER_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20506_ _20638_/CLK _20506_/D vssd1 vssd1 vccd1 vccd1 _20506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20437_ _20718_/CLK _20437_/D vssd1 vssd1 vccd1 vccd1 _20437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ _19663_/Q _10924_/S _11170_/B1 vssd1 vssd1 vccd1 vccd1 _11170_/X sky130_fd_sc_hd__o21a_1
X_20368_ _20565_/CLK _20368_/D vssd1 vssd1 vccd1 vccd1 _20368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10121_ input128/X input164/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10121_/X sky130_fd_sc_hd__mux2_8
XFILLER_106_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20299_ _20300_/CLK _20299_/D vssd1 vssd1 vccd1 vccd1 _20299_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10052_ _20473_/Q _20313_/Q _10485_/S vssd1 vssd1 vccd1 vccd1 _10052_/X sky130_fd_sc_hd__mux2_1
XFILLER_276_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ _10969_/B _12033_/Y _14870_/S vssd1 vssd1 vccd1 vccd1 _14860_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _13816_/A1 _13725_/B _13816_/B1 input227/X vssd1 vssd1 vccd1 vccd1 _13811_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14791_ _19520_/Q _14797_/B vssd1 vssd1 vccd1 vccd1 _14791_/X sky130_fd_sc_hd__or2_1
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16530_ _19831_/Q _16578_/A2 _16578_/B1 input10/X vssd1 vssd1 vccd1 vccd1 _16531_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13742_ _13742_/A _13742_/B _13777_/A vssd1 vssd1 vccd1 vccd1 _13742_/X sky130_fd_sc_hd__or3_1
XFILLER_232_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10954_ _12514_/C _10953_/Y _10950_/Y _12504_/A vssd1 vssd1 vccd1 vccd1 _10954_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16461_ _19770_/Q _17647_/A1 _16471_/S vssd1 vssd1 vccd1 vccd1 _19770_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13673_ _13674_/B vssd1 vssd1 vccd1 vccd1 _13673_/Y sky130_fd_sc_hd__inv_2
X_10885_ _10885_/A _10885_/B vssd1 vssd1 vccd1 vccd1 _15264_/A sky130_fd_sc_hd__nor2_8
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18200_ _18490_/B vssd1 vssd1 vccd1 vccd1 _18200_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15412_ _14882_/B _15406_/Y _15409_/Y _15411_/X _15526_/B vssd1 vssd1 vccd1 vccd1
+ _15412_/X sky130_fd_sc_hd__o2111a_1
X_19180_ _20426_/CLK _19180_/D vssd1 vssd1 vccd1 vccd1 _19180_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12624_ _12624_/A _12624_/B vssd1 vssd1 vccd1 vccd1 _12624_/X sky130_fd_sc_hd__or2_2
X_16392_ _19742_/Q _16394_/C _16391_/Y vssd1 vssd1 vccd1 vccd1 _19742_/D sky130_fd_sc_hd__o21a_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18131_ _14119_/A _19105_/Q _18134_/A vssd1 vssd1 vccd1 vccd1 _18457_/B sky130_fd_sc_hd__mux2_4
X_15343_ _19741_/Q _15453_/A2 _15333_/X _15396_/A1 _15342_/X vssd1 vssd1 vccd1 vccd1
+ _15343_/X sky130_fd_sc_hd__a221o_1
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _12555_/A _12555_/B vssd1 vssd1 vccd1 vccd1 _18472_/B sky130_fd_sc_hd__nor2_8
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18062_ _18064_/A _18062_/B _18063_/B vssd1 vssd1 vccd1 vccd1 _20760_/D sky130_fd_sc_hd__nor3_1
XFILLER_200_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11506_ _20381_/Q _20445_/Q _11527_/S vssd1 vssd1 vccd1 vccd1 _11506_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15274_ _20951_/Q _15322_/C _15568_/B1 _20823_/Q _15273_/X vssd1 vssd1 vccd1 vccd1
+ _15274_/X sky130_fd_sc_hd__a221o_2
X_12486_ _12832_/B _12486_/B vssd1 vssd1 vccd1 vccd1 _12486_/Y sky130_fd_sc_hd__nand2_8
XFILLER_156_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17013_ _09486_/Y _16706_/X _13466_/B _18821_/A vssd1 vssd1 vccd1 vccd1 _19993_/D
+ sky130_fd_sc_hd__a211oi_1
X_14225_ _19225_/Q _14256_/A2 _14224_/X _14758_/C1 vssd1 vssd1 vccd1 vccd1 _19225_/D
+ sky130_fd_sc_hd__o211a_1
X_11437_ _12138_/A1 _20510_/Q _12134_/S _11427_/X vssd1 vssd1 vccd1 vccd1 _11437_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14156_ _20270_/Q _14117_/A _14267_/B1 input241/X vssd1 vssd1 vccd1 vccd1 _14158_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11368_ _11368_/A1 _13664_/A _11367_/X _11398_/S vssd1 vssd1 vccd1 vccd1 _11400_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13107_ _13107_/A _13107_/B vssd1 vssd1 vccd1 vccd1 _13107_/Y sky130_fd_sc_hd__nor2_2
X_10319_ _11270_/A2 _10318_/X _10315_/X _11275_/A vssd1 vssd1 vccd1 vccd1 _10319_/X
+ sky130_fd_sc_hd__o211a_1
X_14087_ _14099_/A _14099_/B _14087_/C vssd1 vssd1 vccd1 vccd1 _14087_/X sky130_fd_sc_hd__or3_1
X_18964_ _21009_/Q _18964_/B vssd1 vssd1 vccd1 vccd1 _18964_/Y sky130_fd_sc_hd__nand2_1
X_11299_ _10262_/A _19334_/Q _20689_/Q _11303_/S _11304_/S vssd1 vssd1 vccd1 vccd1
+ _11299_/X sky130_fd_sc_hd__a221o_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17915_ _20686_/Q _17915_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20686_/D sky130_fd_sc_hd__mux2_1
XFILLER_85_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13038_ _20959_/Q _20893_/Q vssd1 vssd1 vccd1 vccd1 _13290_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18895_ _18640_/Y _18977_/A2 _18893_/Y _18894_/Y vssd1 vssd1 vccd1 vccd1 _18895_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1150 _17107_/A1 vssd1 vssd1 vccd1 vccd1 _17943_/A1 sky130_fd_sc_hd__buf_2
XFILLER_227_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1161 _12403_/B1 vssd1 vssd1 vccd1 vccd1 _12158_/B1 sky130_fd_sc_hd__buf_4
X_17846_ _20621_/Q input247/X _17849_/S vssd1 vssd1 vccd1 vccd1 _20621_/D sky130_fd_sc_hd__mux2_1
Xfanout1172 _16009_/B vssd1 vssd1 vccd1 vccd1 _15528_/B sky130_fd_sc_hd__buf_6
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1183 _12486_/Y vssd1 vssd1 vccd1 vccd1 _16005_/A1 sky130_fd_sc_hd__clkbuf_16
Xfanout1194 _09572_/X vssd1 vssd1 vccd1 vccd1 _11368_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17777_ _20556_/Q _17917_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20556_/D sky130_fd_sc_hd__mux2_1
XFILLER_270_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14989_ input1/X _15021_/B _14986_/C _14988_/Y vssd1 vssd1 vccd1 vccd1 _14989_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_242_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19516_ _20300_/CLK _19516_/D vssd1 vssd1 vccd1 vccd1 _19516_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16728_ _09518_/Y _16799_/S _16726_/X _16727_/Y vssd1 vssd1 vccd1 vccd1 _16728_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_34_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19447_ _20574_/CLK _19447_/D vssd1 vssd1 vccd1 vccd1 _19447_/Q sky130_fd_sc_hd__dfxtp_1
X_16659_ _19916_/Q _17871_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19916_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19378_ _20669_/CLK _19378_/D vssd1 vssd1 vccd1 vccd1 _19378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18329_ _18466_/B _18341_/B vssd1 vssd1 vccd1 vccd1 _18329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_96_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20759_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20222_ _21018_/CLK _20222_/D vssd1 vssd1 vccd1 vccd1 _20222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20153_ _20692_/CLK _20153_/D vssd1 vssd1 vccd1 vccd1 _20153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09964_ _11903_/A1 _09957_/X _09958_/X vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__o21a_1
XFILLER_281_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20084_ _20084_/CLK _20084_/D vssd1 vssd1 vccd1 vccd1 _20084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _12143_/S _09894_/X _09893_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _09895_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_506 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_517 input246/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_528 _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _21013_/CLK _20986_/D vssd1 vssd1 vccd1 vccd1 _20986_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_539 _11192_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10670_ _12391_/S _10669_/X _10668_/X _12399_/A1 vssd1 vssd1 vccd1 vccd1 _10670_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_201_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12340_ _12338_/X _12339_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _12340_/X sky130_fd_sc_hd__mux2_2
XFILLER_127_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12271_ _20330_/Q _11379_/B _12270_/X vssd1 vssd1 vccd1 vccd1 _12271_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14010_ _13192_/A _14043_/A2 _14034_/B1 _14009_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1
+ _19170_/D sky130_fd_sc_hd__o221a_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ _15067_/S _11223_/B vssd1 vssd1 vccd1 vccd1 _11224_/B sky130_fd_sc_hd__nor2_1
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11153_ _18765_/A _19303_/Q _11174_/S _19799_/Q _11353_/C1 vssd1 vssd1 vccd1 vccd1
+ _11155_/B sky130_fd_sc_hd__o221a_1
XFILLER_134_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10104_ _19810_/Q _12085_/A2 _10102_/X _12085_/B2 _10103_/X vssd1 vssd1 vccd1 vccd1
+ _10104_/X sky130_fd_sc_hd__o221a_1
X_11084_ _12324_/S _11083_/X _11082_/X _12314_/C1 vssd1 vssd1 vccd1 vccd1 _11084_/X
+ sky130_fd_sc_hd__a211o_1
X_15961_ _19730_/Q _15961_/A2 _15961_/B1 _19762_/Q vssd1 vssd1 vccd1 vccd1 _15961_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput220 localMemory_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_hd__buf_12
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput231 localMemory_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_hd__buf_12
XFILLER_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14912_ _18149_/S _14912_/B vssd1 vssd1 vccd1 vccd1 _14912_/X sky130_fd_sc_hd__and2b_1
X_10035_ _11236_/A split7/A _11326_/A vssd1 vssd1 vccd1 vccd1 _10035_/Y sky130_fd_sc_hd__a21oi_4
Xinput242 localMemory_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_hd__buf_12
X_17700_ _20484_/Q _17943_/A1 _17705_/S vssd1 vssd1 vccd1 vccd1 _20484_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput253 manufacturerID[0] vssd1 vssd1 vccd1 vccd1 _17239_/A sky130_fd_sc_hd__buf_4
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18680_ _18553_/X _18684_/A2 _18678_/Y _18679_/Y vssd1 vssd1 vccd1 vccd1 _18681_/B
+ sky130_fd_sc_hd__o211a_1
X_15892_ _12290_/A _16028_/C _15891_/X _15890_/B vssd1 vssd1 vccd1 vccd1 _15893_/C
+ sky130_fd_sc_hd__a211o_1
Xinput264 partID[0] vssd1 vssd1 vccd1 vccd1 _17272_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput275 partID[5] vssd1 vssd1 vccd1 vccd1 _17287_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17631_ _20387_/Q _17802_/A1 _17635_/S vssd1 vssd1 vccd1 vccd1 _20387_/D sky130_fd_sc_hd__mux2_1
X_14843_ _11742_/B _10640_/B _14843_/S vssd1 vssd1 vccd1 vccd1 _14843_/X sky130_fd_sc_hd__mux2_1
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17562_ _20322_/Q _17801_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20322_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14774_ _19134_/Q _14774_/A2 _14773_/X _14776_/C1 vssd1 vssd1 vccd1 vccd1 _19511_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11986_ _20424_/Q _20360_/Q _11987_/S vssd1 vssd1 vccd1 vccd1 _11986_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19301_ _20721_/CLK _19301_/D vssd1 vssd1 vccd1 vccd1 _19301_/Q sky130_fd_sc_hd__dfxtp_1
X_16513_ _19820_/Q _17874_/A1 _16517_/S vssd1 vssd1 vccd1 vccd1 _19820_/D sky130_fd_sc_hd__mux2_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13725_ _13780_/A _13725_/B vssd1 vssd1 vccd1 vccd1 _13725_/X sky130_fd_sc_hd__and2_1
X_10937_ _10937_/A _19306_/Q _11021_/C vssd1 vssd1 vccd1 vccd1 _10937_/X sky130_fd_sc_hd__or3_1
XFILLER_16_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17493_ _17495_/A1 _17492_/Y _18863_/A vssd1 vssd1 vccd1 vccd1 _20281_/D sky130_fd_sc_hd__a21oi_1
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19232_ _19232_/CLK _19232_/D vssd1 vssd1 vccd1 vccd1 _19232_/Q sky130_fd_sc_hd__dfxtp_2
X_16444_ _19762_/Q _16444_/B vssd1 vssd1 vccd1 vccd1 _16450_/C sky130_fd_sc_hd__and2_4
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _13775_/A _13656_/B vssd1 vssd1 vccd1 vccd1 _13656_/X sky130_fd_sc_hd__and2_1
X_10868_ _12332_/A _19467_/Q _19435_/Q _12352_/S _12347_/C1 vssd1 vssd1 vccd1 vccd1
+ _10868_/X sky130_fd_sc_hd__a221o_1
X_19163_ _20659_/CLK _19163_/D vssd1 vssd1 vccd1 vccd1 _19163_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_220_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12607_ _19512_/Q _12845_/A vssd1 vssd1 vccd1 vccd1 _12835_/A sky130_fd_sc_hd__and2_4
X_16375_ _19736_/Q _16378_/C _18054_/A vssd1 vssd1 vccd1 vccd1 _16375_/Y sky130_fd_sc_hd__a21oi_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _19224_/Q _13587_/B vssd1 vssd1 vccd1 vccd1 _13587_/X sky130_fd_sc_hd__xor2_1
XFILLER_185_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10799_ _10799_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__or2_4
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18114_ _20780_/Q _18117_/C _18112_/A vssd1 vssd1 vccd1 vccd1 _18114_/Y sky130_fd_sc_hd__a21oi_1
X_15326_ _15326_/A _15326_/B _15326_/C vssd1 vssd1 vccd1 vccd1 _15326_/X sky130_fd_sc_hd__or3_1
XFILLER_118_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19094_ _19620_/CLK _19094_/D vssd1 vssd1 vccd1 vccd1 _19094_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_145_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12538_ _20880_/Q _12549_/B _12538_/C vssd1 vssd1 vccd1 vccd1 _12551_/B sky130_fd_sc_hd__and3_1
XFILLER_173_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18045_ _20754_/Q _20753_/Q _18045_/C vssd1 vssd1 vccd1 vccd1 _18047_/B sky130_fd_sc_hd__and3_1
XFILLER_144_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15257_ _15066_/S _15255_/X _15256_/X vssd1 vssd1 vccd1 vccd1 _15258_/B sky130_fd_sc_hd__a21oi_2
X_12469_ _16058_/A2 _16057_/A2 _12469_/S vssd1 vssd1 vccd1 vccd1 _12469_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14208_ _19503_/Q _14208_/B vssd1 vssd1 vccd1 vccd1 _14209_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15188_ _12342_/A _12658_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _15188_/X sky130_fd_sc_hd__mux2_1
XFILLER_259_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14139_ _19496_/Q _14139_/B vssd1 vssd1 vccd1 vccd1 _14140_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19996_ _20621_/CLK _19996_/D vssd1 vssd1 vccd1 vccd1 _19996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18947_ _19111_/Q _18974_/A2 _18967_/B1 _15949_/B vssd1 vssd1 vccd1 vccd1 _18948_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09680_ _11326_/A _09680_/B _09680_/C vssd1 vssd1 vccd1 vccd1 _09680_/X sky130_fd_sc_hd__and3_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18878_ _19101_/Q _18954_/A2 _18967_/B1 _13427_/B vssd1 vssd1 vccd1 vccd1 _18879_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_143_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19228_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_251_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17829_ _20604_/Q _17901_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20604_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20840_ _20969_/CLK _20840_/D vssd1 vssd1 vccd1 vccd1 _20840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20771_ _20862_/CLK _20771_/D vssd1 vssd1 vccd1 vccd1 _20771_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_251_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20205_ _20760_/CLK _20205_/D vssd1 vssd1 vccd1 vccd1 _20205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout910 _14996_/X vssd1 vssd1 vccd1 vccd1 _15601_/S sky130_fd_sc_hd__clkbuf_4
Xfanout1908 _13887_/C1 vssd1 vssd1 vccd1 vccd1 _16167_/C1 sky130_fd_sc_hd__buf_6
XFILLER_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout921 _14945_/Y vssd1 vssd1 vccd1 vccd1 _15934_/A2 sky130_fd_sc_hd__buf_12
Xfanout1919 _09515_/Y vssd1 vssd1 vccd1 vccd1 _13887_/C1 sky130_fd_sc_hd__buf_12
X_20136_ _20715_/CLK _20136_/D vssd1 vssd1 vccd1 vccd1 _20136_/Q sky130_fd_sc_hd__dfxtp_1
X_09947_ _12156_/A1 _09946_/X _09942_/X vssd1 vssd1 vccd1 vccd1 _09947_/X sky130_fd_sc_hd__a21o_4
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout932 _15039_/A vssd1 vssd1 vccd1 vccd1 _15058_/S sky130_fd_sc_hd__buf_8
XFILLER_131_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout943 _11102_/X vssd1 vssd1 vccd1 vccd1 _11137_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout954 _14262_/A vssd1 vssd1 vccd1 vccd1 _14427_/A sky130_fd_sc_hd__buf_4
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout965 _10562_/X vssd1 vssd1 vccd1 vccd1 _17895_/A1 sky130_fd_sc_hd__clkbuf_8
X_20067_ _20694_/CLK _20067_/D vssd1 vssd1 vccd1 vccd1 _20067_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout976 _17691_/A1 vssd1 vssd1 vccd1 vccd1 _17657_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_218_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout987 _17096_/A1 vssd1 vssd1 vccd1 vccd1 _17689_/A1 sky130_fd_sc_hd__clkbuf_4
X_09878_ _20482_/Q _20322_/Q _11527_/S vssd1 vssd1 vccd1 vccd1 _09878_/X sky130_fd_sc_hd__mux2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 _16709_/X vssd1 vssd1 vccd1 vccd1 _16862_/A2 sky130_fd_sc_hd__buf_4
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _12144_/C1 _11829_/X _11832_/X _11839_/X _12152_/A1 vssd1 vssd1 vccd1 vccd1
+ _11840_/X sky130_fd_sc_hd__a311o_1
XANTENNA_303 input230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_314 input246/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_325 _13643_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_336 _19507_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 _11397_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11771_ _13567_/A _11771_/B vssd1 vssd1 vccd1 vccd1 _11788_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_358 _12131_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _20969_/CLK _20969_/D vssd1 vssd1 vccd1 vccd1 _20969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_369 _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _13624_/B2 _13497_/Y _13509_/Y _19661_/D vssd1 vssd1 vccd1 vccd1 _13510_/X
+ sky130_fd_sc_hd__a22o_4
X_10722_ _10373_/A _10285_/Y _09659_/B vssd1 vssd1 vccd1 vccd1 _10722_/X sky130_fd_sc_hd__a21o_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _19268_/Q _17678_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19268_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13441_ _14525_/B _13440_/X _15843_/A _13437_/A _16066_/B vssd1 vssd1 vccd1 vccd1
+ _13441_/X sky130_fd_sc_hd__a2111o_1
X_10653_ _20125_/Q _20093_/Q _12368_/S vssd1 vssd1 vccd1 vccd1 _10653_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16160_ _16851_/B _16164_/B vssd1 vssd1 vccd1 vccd1 _16160_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13372_ _18767_/A _13363_/Y _13366_/X _13371_/X vssd1 vssd1 vccd1 vccd1 _13373_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10584_ _20534_/Q _20502_/Q _12064_/S vssd1 vssd1 vccd1 vccd1 _10584_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15111_ _14816_/X _14851_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _15111_/X sky130_fd_sc_hd__mux2_1
X_12323_ _19298_/Q _20085_/Q _12323_/S vssd1 vssd1 vccd1 vccd1 _12323_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16091_ _19570_/Q _16079_/B _16107_/B1 vssd1 vssd1 vccd1 vccd1 _16091_/X sky130_fd_sc_hd__o21a_1
XFILLER_182_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15042_ _15037_/X _15041_/Y _15254_/S vssd1 vssd1 vccd1 vccd1 _15042_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12254_ _12254_/A _20686_/Q _12254_/C vssd1 vssd1 vccd1 vccd1 _12254_/X sky130_fd_sc_hd__or3_1
XFILLER_253_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11205_ _19399_/Q _20558_/Q _11211_/S vssd1 vssd1 vccd1 vccd1 _11205_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19850_ _20014_/CLK _19850_/D vssd1 vssd1 vccd1 vccd1 _19850_/Q sky130_fd_sc_hd__dfxtp_4
X_12185_ _19362_/Q _20717_/Q _12185_/S vssd1 vssd1 vccd1 vccd1 _12185_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18801_ _18801_/A _18801_/B vssd1 vssd1 vccd1 vccd1 _20985_/D sky130_fd_sc_hd__nor2_1
XFILLER_123_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11136_ _11137_/A _11136_/B vssd1 vssd1 vccd1 vccd1 _11136_/X sky130_fd_sc_hd__and2_1
X_19781_ _20702_/CLK _19781_/D vssd1 vssd1 vccd1 vccd1 _19781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16993_ _16990_/Y _16992_/Y _17011_/B1 vssd1 vssd1 vccd1 vccd1 _16993_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_62_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18732_ _18748_/A _18732_/B vssd1 vssd1 vccd1 vccd1 _20966_/D sky130_fd_sc_hd__and2_1
XFILLER_49_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ _12396_/A1 _19464_/Q _19432_/Q _11090_/S _12371_/C1 vssd1 vssd1 vccd1 vccd1
+ _11067_/X sky130_fd_sc_hd__a221o_1
X_15944_ _15973_/A1 _15943_/X _15931_/Y vssd1 vssd1 vccd1 vccd1 _15944_/X sky130_fd_sc_hd__a21o_1
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10018_ _11761_/B vssd1 vssd1 vccd1 vccd1 _10018_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15875_ _21037_/Q _21005_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _15875_/X sky130_fd_sc_hd__mux2_1
X_18663_ _19519_/Q _18667_/B vssd1 vssd1 vccd1 vccd1 _18663_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17614_ _20370_/Q _17751_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20370_/D sky130_fd_sc_hd__mux2_1
XFILLER_252_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _11322_/B _12114_/B _14836_/S vssd1 vssd1 vccd1 vccd1 _14826_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18594_ _18592_/Y _18593_/X _18598_/A vssd1 vssd1 vccd1 vccd1 _20921_/D sky130_fd_sc_hd__a21oi_1
XFILLER_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17545_ _20305_/Q _17750_/A1 _17570_/S vssd1 vssd1 vccd1 vccd1 _20305_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14757_ _19503_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14757_/X sky130_fd_sc_hd__or2_1
XFILLER_189_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11969_ _11977_/A1 _11967_/X _11968_/X vssd1 vssd1 vccd1 vccd1 _11969_/X sky130_fd_sc_hd__o21a_1
XFILLER_251_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13708_ _13718_/A _13708_/B vssd1 vssd1 vccd1 vccd1 _13708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_260_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17476_ _20273_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17476_/Y sky130_fd_sc_hd__nand2_1
X_14688_ _19447_/Q _17937_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19447_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19215_ _19219_/CLK _19215_/D vssd1 vssd1 vccd1 vccd1 _19215_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16427_ _18096_/A _16427_/B _16428_/B vssd1 vssd1 vccd1 vccd1 _19755_/D sky130_fd_sc_hd__nor3_1
X_13639_ _13658_/A _16054_/B _15076_/A _14525_/B _13637_/C vssd1 vssd1 vccd1 vccd1
+ _16239_/B sky130_fd_sc_hd__o311a_4
XFILLER_177_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16358_ _16362_/C _16358_/B vssd1 vssd1 vccd1 vccd1 _19729_/D sky130_fd_sc_hd__nor2_1
X_19146_ _19523_/CLK _19146_/D vssd1 vssd1 vccd1 vccd1 _19146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15309_ _21018_/Q _20986_/Q _15309_/S vssd1 vssd1 vccd1 vccd1 _15309_/X sky130_fd_sc_hd__mux2_1
X_16289_ _19702_/Q _19703_/Q _19704_/Q vssd1 vssd1 vccd1 vccd1 _16294_/C sky130_fd_sc_hd__and3_2
XFILLER_145_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19077_ _20422_/Q vssd1 vssd1 vccd1 vccd1 _20422_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18028_ _18112_/A _18028_/B vssd1 vssd1 vccd1 vccd1 _18028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09801_ _19951_/Q _12043_/B vssd1 vssd1 vccd1 vccd1 _09801_/X sky130_fd_sc_hd__or2_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19979_ _20014_/CLK _19979_/D vssd1 vssd1 vccd1 vccd1 _19979_/Q sky130_fd_sc_hd__dfxtp_1
X_09732_ _10516_/S _09734_/B vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__nor2_8
XFILLER_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09663_ input113/X input148/X _11241_/S vssd1 vssd1 vccd1 vccd1 _09664_/C sky130_fd_sc_hd__mux2_8
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09594_ _09583_/A _19086_/Q _09588_/C _09593_/X _09588_/X vssd1 vssd1 vccd1 vccd1
+ _09594_/X sky130_fd_sc_hd__a41o_2
XFILLER_270_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _21017_/CLK _20823_/D vssd1 vssd1 vccd1 vccd1 _20823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20754_ _20794_/CLK _20754_/D vssd1 vssd1 vccd1 vccd1 _20754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20685_ _20685_/CLK _20685_/D vssd1 vssd1 vccd1 vccd1 _20685_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_40_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20557_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1705 _11537_/A1 vssd1 vssd1 vccd1 vccd1 _12016_/C1 sky130_fd_sc_hd__buf_6
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1716 _11309_/A1 vssd1 vssd1 vccd1 vccd1 _10516_/S sky130_fd_sc_hd__buf_12
XFILLER_278_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1727 _18765_/A vssd1 vssd1 vccd1 vccd1 _11273_/A1 sky130_fd_sc_hd__buf_6
XFILLER_265_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout740 _14204_/A vssd1 vssd1 vccd1 vccd1 _14255_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_120_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1738 _09503_/Y vssd1 vssd1 vccd1 vccd1 _11423_/C1 sky130_fd_sc_hd__buf_8
Xfanout751 _18458_/X vssd1 vssd1 vccd1 vccd1 _18559_/B sky130_fd_sc_hd__clkbuf_4
Xfanout1749 _09501_/Y vssd1 vssd1 vccd1 vccd1 _12046_/B1 sky130_fd_sc_hd__buf_6
XFILLER_131_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20119_ _20561_/CLK _20119_/D vssd1 vssd1 vccd1 vccd1 _20119_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout762 _18565_/Y vssd1 vssd1 vccd1 vccd1 _18686_/B sky130_fd_sc_hd__buf_4
X_13990_ _14041_/A1 _09664_/B _10281_/X _14041_/B1 _19845_/Q vssd1 vssd1 vccd1 vccd1
+ _14073_/C sky130_fd_sc_hd__o32a_1
Xfanout773 _18902_/A vssd1 vssd1 vccd1 vccd1 _18560_/A sky130_fd_sc_hd__buf_4
XFILLER_59_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout784 _12592_/X vssd1 vssd1 vccd1 vccd1 _18490_/A sky130_fd_sc_hd__buf_4
Xfanout795 _12652_/B vssd1 vssd1 vccd1 vccd1 _13589_/A1 sky130_fd_sc_hd__clkbuf_8
X_12941_ _19254_/Q _12964_/A2 _16945_/B _20002_/Q vssd1 vssd1 vccd1 vccd1 _14915_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15660_ _19719_/Q _15989_/A2 _15989_/B1 _19751_/Q vssd1 vssd1 vccd1 vccd1 _15660_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _19518_/Q _12872_/B vssd1 vssd1 vccd1 vccd1 _12873_/B sky130_fd_sc_hd__nor2_1
XANTENNA_100 _16009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 _13909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_122 _13708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _19375_/Q _17895_/A1 _14628_/S vssd1 vssd1 vccd1 vccd1 _19375_/D sky130_fd_sc_hd__mux2_1
X_11823_ _11815_/X _11816_/X _11902_/S vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__mux2_1
XANTENNA_133 _13683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 _13725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15591_/A _15591_/B vssd1 vssd1 vccd1 vccd1 _15591_/Y sky130_fd_sc_hd__nand2_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 _13780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 _14737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _20215_/Q _17330_/A2 _17305_/C _17329_/X _17330_/C1 vssd1 vssd1 vccd1 vccd1
+ _17330_/X sky130_fd_sc_hd__a221o_1
XFILLER_26_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14542_ _19312_/Q _17060_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19312_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _19114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 _19166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11754_ _11754_/A _11754_/B vssd1 vssd1 vccd1 vccd1 _11790_/B sky130_fd_sc_hd__nor2_1
XANTENNA_199 _20420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _20192_/Q _17330_/A2 _17269_/C _17260_/Y _17279_/C1 vssd1 vssd1 vccd1 vccd1
+ _17261_/X sky130_fd_sc_hd__a221o_1
X_10705_ _20157_/Q _11379_/B vssd1 vssd1 vccd1 vccd1 _10705_/X sky130_fd_sc_hd__or2_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14473_ _20232_/Q _19261_/Q _14477_/S vssd1 vssd1 vccd1 vccd1 _14474_/B sky130_fd_sc_hd__mux2_1
X_11685_ _12073_/A1 _11674_/X _11677_/X _11684_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1
+ _11685_/X sky130_fd_sc_hd__a311o_1
X_19000_ _18195_/Y _18982_/B _19016_/B1 _18999_/X vssd1 vssd1 vccd1 vccd1 _21019_/D
+ sky130_fd_sc_hd__o211a_1
X_16212_ _19635_/Q _17096_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19635_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13424_ _13424_/A _13424_/B vssd1 vssd1 vccd1 vccd1 _13426_/C sky130_fd_sc_hd__xnor2_4
X_17192_ _20156_/Q _17926_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20156_/D sky130_fd_sc_hd__mux2_1
X_10636_ _10638_/B vssd1 vssd1 vccd1 vccd1 _10636_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _16143_/A _16143_/B vssd1 vssd1 vccd1 vccd1 _19595_/D sky130_fd_sc_hd__and2_1
XFILLER_128_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13355_ _20962_/Q _13355_/B vssd1 vssd1 vccd1 vccd1 _13355_/Y sky130_fd_sc_hd__nand2_1
X_10567_ _19671_/Q _11682_/S _10566_/X _12051_/C1 vssd1 vssd1 vccd1 vccd1 _10567_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ _12306_/A1 _19461_/Q _12300_/S _12305_/X vssd1 vssd1 vccd1 vccd1 _12306_/X
+ sky130_fd_sc_hd__a31o_1
X_16074_ _19561_/Q _16081_/B _16073_/Y _16195_/A vssd1 vssd1 vccd1 vccd1 _19561_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ _19228_/Q _19227_/Q _13450_/A vssd1 vssd1 vccd1 vccd1 _13378_/B sky130_fd_sc_hd__and3_1
X_10498_ _19939_/Q _11270_/A2 _10897_/A3 _11250_/S vssd1 vssd1 vccd1 vccd1 _10498_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_170_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19902_ _20085_/CLK _19902_/D vssd1 vssd1 vccd1 vccd1 _19902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15025_ _15026_/A _15095_/B vssd1 vssd1 vccd1 vccd1 _15025_/X sky130_fd_sc_hd__and2_1
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ _19827_/Q _19331_/Q _12316_/S vssd1 vssd1 vccd1 vccd1 _12237_/X sky130_fd_sc_hd__mux2_1
XFILLER_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19833_ _20004_/CLK _19833_/D vssd1 vssd1 vccd1 vccd1 _19833_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12168_ _11846_/C _12163_/X _12167_/X _09839_/A vssd1 vssd1 vccd1 vccd1 _12168_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11119_ _19867_/Q _19768_/Q _11126_/B vssd1 vssd1 vccd1 vccd1 _11119_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19764_ _20268_/CLK _19764_/D vssd1 vssd1 vccd1 vccd1 _19764_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_96_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16976_ _16950_/Y _16975_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16976_/Y sky130_fd_sc_hd__o21bai_4
X_12099_ _12103_/A1 _12097_/X _12098_/X vssd1 vssd1 vccd1 vccd1 _12099_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_284_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18715_ _20958_/Q _18220_/Y _18719_/S vssd1 vssd1 vccd1 vccd1 _18716_/B sky130_fd_sc_hd__mux2_1
Xinput6 coreIndex[5] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_4
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15927_ _12036_/B _12466_/Y _12471_/X _12288_/A _15365_/A vssd1 vssd1 vccd1 vccd1
+ _15927_/X sky130_fd_sc_hd__o221a_1
XFILLER_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19695_ _19695_/CLK _19695_/D vssd1 vssd1 vccd1 vccd1 _19695_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_49_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18646_ _20935_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18646_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ _16017_/C1 _15857_/X _15853_/X vssd1 vssd1 vccd1 vccd1 _15858_/X sky130_fd_sc_hd__o21a_2
XFILLER_213_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14809_ _14809_/A _15246_/A vssd1 vssd1 vccd1 vccd1 _14809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_206_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18577_ _20917_/Q _18592_/B vssd1 vssd1 vccd1 vccd1 _18577_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15789_ _15789_/A _15789_/B _15981_/B vssd1 vssd1 vccd1 vccd1 _15789_/X sky130_fd_sc_hd__and3_1
XFILLER_178_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17528_ _20299_/Q _17528_/B _17528_/C vssd1 vssd1 vccd1 vccd1 _17528_/X sky130_fd_sc_hd__or3_1
XFILLER_221_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17459_ _17452_/A _17456_/Y _17457_/X _17458_/X vssd1 vssd1 vccd1 vccd1 _17459_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20470_ _20679_/CLK _20470_/D vssd1 vssd1 vccd1 vccd1 _20470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19129_ _19506_/CLK _19129_/D vssd1 vssd1 vccd1 vccd1 _19129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput310 _13617_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[14] sky130_fd_sc_hd__buf_4
Xoutput321 _13627_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[24] sky130_fd_sc_hd__buf_4
Xoutput332 _13597_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[9] sky130_fd_sc_hd__buf_4
XFILLER_273_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput343 _13716_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[18] sky130_fd_sc_hd__buf_4
Xoutput354 _13765_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[28] sky130_fd_sc_hd__buf_4
Xoutput365 _13674_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[9] sky130_fd_sc_hd__buf_4
Xoutput376 _13791_/X vssd1 vssd1 vccd1 vccd1 din0[0] sky130_fd_sc_hd__buf_6
XFILLER_0_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21022_ _21022_/CLK _21022_/D vssd1 vssd1 vccd1 vccd1 _21022_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput387 _13792_/X vssd1 vssd1 vccd1 vccd1 din0[1] sky130_fd_sc_hd__buf_6
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput398 _13793_/X vssd1 vssd1 vccd1 vccd1 din0[2] sky130_fd_sc_hd__buf_6
XFILLER_87_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09715_ _11988_/S _09714_/X _09713_/X _12144_/A1 vssd1 vssd1 vccd1 vccd1 _09715_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09646_ _19658_/Q _19695_/Q vssd1 vssd1 vccd1 vccd1 _09646_/Y sky130_fd_sc_hd__nand2_2
XFILLER_283_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09577_ _12967_/B _19096_/Q _09609_/A vssd1 vssd1 vccd1 vccd1 _10020_/B sky130_fd_sc_hd__o21ba_2
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20806_ _21029_/CLK _20806_/D vssd1 vssd1 vccd1 vccd1 _20806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20737_ _20860_/CLK _20737_/D vssd1 vssd1 vccd1 vccd1 _20737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ _19640_/Q _19946_/Q _12182_/S vssd1 vssd1 vccd1 vccd1 _11471_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20668_ _20668_/CLK _20668_/D vssd1 vssd1 vccd1 vccd1 _20668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10421_ _10419_/X _10420_/X _12071_/S vssd1 vssd1 vccd1 vccd1 _10421_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20599_ _20635_/CLK _20599_/D vssd1 vssd1 vccd1 vccd1 _20599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ _19214_/Q _13140_/B vssd1 vssd1 vccd1 vccd1 _13242_/B sky130_fd_sc_hd__or2_4
XFILLER_152_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10352_ _20411_/Q _20347_/Q _20639_/Q _20603_/Q _11203_/S _11026_/C vssd1 vssd1 vccd1
+ vccd1 _10352_/X sky130_fd_sc_hd__mux4_1
XFILLER_124_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13071_ _13039_/Y _13316_/A _13315_/B vssd1 vssd1 vccd1 vccd1 _13290_/C sky130_fd_sc_hd__o21ai_4
X_10283_ _19573_/Q _10282_/X _11243_/S vssd1 vssd1 vccd1 vccd1 _10283_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12022_ _20145_/Q _20113_/Q _12025_/S vssd1 vssd1 vccd1 vccd1 _12022_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1502 _12041_/B vssd1 vssd1 vccd1 vccd1 _12213_/B sky130_fd_sc_hd__buf_8
XFILLER_183_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1513 fanout1534/X vssd1 vssd1 vccd1 vccd1 _11599_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_266_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1524 _11665_/S vssd1 vssd1 vccd1 vccd1 _11978_/S sky130_fd_sc_hd__buf_6
XFILLER_278_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1535 _10303_/S vssd1 vssd1 vccd1 vccd1 _11255_/S sky130_fd_sc_hd__buf_6
X_16830_ _16932_/B1 _16827_/X _16829_/X _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16831_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1546 fanout1566/X vssd1 vssd1 vccd1 vccd1 _10316_/S sky130_fd_sc_hd__buf_4
Xfanout1557 _11358_/S vssd1 vssd1 vccd1 vccd1 _12296_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_66_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout570 _16490_/X vssd1 vssd1 vccd1 vccd1 _16522_/S sky130_fd_sc_hd__buf_12
Xfanout1568 _09625_/Y vssd1 vssd1 vccd1 vccd1 _12073_/A1 sky130_fd_sc_hd__buf_4
XFILLER_266_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1579 _09688_/A vssd1 vssd1 vccd1 vccd1 _11274_/B2 sky130_fd_sc_hd__buf_6
Xfanout581 _16199_/X vssd1 vssd1 vccd1 vccd1 _16227_/S sky130_fd_sc_hd__buf_4
XFILLER_47_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout592 _14704_/X vssd1 vssd1 vccd1 vccd1 _14733_/S sky130_fd_sc_hd__buf_8
X_13973_ _19190_/Q _14061_/C _14003_/S vssd1 vssd1 vccd1 vccd1 _13973_/X sky130_fd_sc_hd__mux2_1
X_16761_ _16726_/X _16760_/Y _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16761_/X sky130_fd_sc_hd__a21o_2
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18500_ _20893_/Q _18474_/S _18499_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18501_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12924_ _14237_/A2 _17461_/A vssd1 vssd1 vccd1 vccd1 _12962_/S sky130_fd_sc_hd__nand2b_4
X_15712_ _15710_/Y _15711_/X _15708_/Y vssd1 vssd1 vccd1 vccd1 _15712_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_206_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19480_ _20081_/CLK _19480_/D vssd1 vssd1 vccd1 vccd1 _19480_/Q sky130_fd_sc_hd__dfxtp_1
X_16692_ _19947_/Q _17695_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19947_/D sky130_fd_sc_hd__mux2_1
XFILLER_234_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18431_ _20870_/Q _18260_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18432_/B sky130_fd_sc_hd__mux2_1
X_15643_ _16049_/A1 _15631_/X _15642_/X vssd1 vssd1 vccd1 vccd1 _16878_/B sky130_fd_sc_hd__a21oi_4
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12855_ _19510_/Q _12855_/B vssd1 vssd1 vccd1 vccd1 _12855_/X sky130_fd_sc_hd__xor2_2
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11806_ _12039_/A1 _11236_/C split7/X vssd1 vssd1 vccd1 vccd1 _11806_/X sky130_fd_sc_hd__a21o_4
XFILLER_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15574_ _15606_/A1 _15563_/X _15573_/X vssd1 vssd1 vccd1 vccd1 _16860_/B sky130_fd_sc_hd__a21oi_4
XFILLER_61_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18362_ _20836_/Q _18363_/B _18361_/Y _18728_/A vssd1 vssd1 vccd1 vccd1 _20836_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12786_ _19503_/Q _12786_/B vssd1 vssd1 vccd1 vccd1 _12786_/X sky130_fd_sc_hd__and2_1
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _20210_/Q _17328_/A2 _17312_/X _17974_/B1 vssd1 vssd1 vccd1 vccd1 _20210_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _19299_/Q _14525_/B _14738_/B vssd1 vssd1 vccd1 vccd1 _14525_/X sky130_fd_sc_hd__and3_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11651_/A _11737_/B vssd1 vssd1 vccd1 vccd1 _11737_/Y sky130_fd_sc_hd__nand2b_1
X_18293_ _19554_/Q _18313_/B vssd1 vssd1 vccd1 vccd1 _18293_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_30_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17244_ _20187_/Q _17268_/A2 _17242_/X _17243_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1
+ _20187_/D sky130_fd_sc_hd__o221a_1
X_14456_ _18692_/A _14456_/B vssd1 vssd1 vccd1 vccd1 _19252_/D sky130_fd_sc_hd__and2_1
XFILLER_175_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11668_ _11660_/X _11661_/X _12056_/S vssd1 vssd1 vccd1 vccd1 _11668_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13407_ _13033_/X _13034_/Y _13073_/Y _13355_/B _13406_/Y vssd1 vssd1 vccd1 vccd1
+ _13407_/Y sky130_fd_sc_hd__a311oi_2
X_17175_ _20141_/Q _17666_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20141_/D sky130_fd_sc_hd__mux2_1
X_10619_ _20374_/Q _20438_/Q _10622_/S vssd1 vssd1 vccd1 vccd1 _10619_/X sky130_fd_sc_hd__mux2_1
X_14387_ _14383_/B _14386_/X _14417_/S vssd1 vssd1 vccd1 vccd1 _14387_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11599_ _19385_/Q _20676_/Q _11599_/S vssd1 vssd1 vccd1 vccd1 _11599_/X sky130_fd_sc_hd__mux2_1
X_16126_ _10039_/X _16126_/A2 _16125_/X vssd1 vssd1 vccd1 vccd1 _19587_/D sky130_fd_sc_hd__o21a_1
X_13338_ _20931_/Q _13350_/B _13323_/C _13337_/X _18628_/B vssd1 vssd1 vccd1 vccd1
+ _13338_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_143_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16057_ _14882_/A _16057_/A2 _12440_/A vssd1 vssd1 vccd1 vccd1 _16057_/X sky130_fd_sc_hd__a21bo_1
X_13269_ _13334_/A _13264_/X _13265_/Y _13268_/X vssd1 vssd1 vccd1 vccd1 _13269_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_143_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _19702_/Q _15454_/S _14949_/X _15007_/X _14941_/X vssd1 vssd1 vccd1 vccd1
+ _15008_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_142_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19816_ _20081_/CLK _19816_/D vssd1 vssd1 vccd1 vccd1 _19816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19747_ _20856_/CLK _19747_/D vssd1 vssd1 vccd1 vccd1 _19747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16959_ input60/X input95/X _17009_/S vssd1 vssd1 vccd1 vccd1 _16959_/X sky130_fd_sc_hd__mux2_8
XFILLER_271_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09500_ _19179_/Q vssd1 vssd1 vccd1 vccd1 _12517_/C sky130_fd_sc_hd__inv_6
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19678_ _20482_/CLK _19678_/D vssd1 vssd1 vccd1 vccd1 _19678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18629_ _18514_/X _18688_/A2 _18627_/Y _18628_/Y vssd1 vssd1 vccd1 vccd1 _18630_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_253_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_11 _15431_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_22 _15600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20522_ _20686_/CLK _20522_/D vssd1 vssd1 vccd1 vccd1 _20522_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_33 _15890_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_44 _16856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 _16977_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_66 _18315_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_77 _09625_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20453_ _21046_/A _20453_/D vssd1 vssd1 vccd1 vccd1 _20453_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_88 _11610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_99 _16009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_284_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20384_ _20480_/CLK _20384_/D vssd1 vssd1 vccd1 vccd1 _20384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21005_ _21009_/CLK _21005_/D vssd1 vssd1 vccd1 vccd1 _21005_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10970_ _10968_/Y _15226_/A vssd1 vssd1 vccd1 vccd1 _13523_/A sky130_fd_sc_hd__nand2b_4
XFILLER_216_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09629_ _16454_/A _11169_/B vssd1 vssd1 vccd1 vccd1 _09630_/D sky130_fd_sc_hd__xnor2_1
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _14803_/A1 _12657_/A2 _12682_/B _12639_/X vssd1 vssd1 vccd1 vccd1 _12640_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ _12513_/A _12513_/B _12588_/A _12570_/X _12464_/C vssd1 vssd1 vccd1 vccd1
+ _12574_/B sky130_fd_sc_hd__o311a_1
XFILLER_196_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14310_ _20285_/Q _14330_/A2 _14330_/B1 input225/X vssd1 vssd1 vccd1 vccd1 _14312_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_197_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11522_ _11902_/S _11521_/X _11520_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _11522_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15290_ _15068_/X _15289_/X _15577_/S vssd1 vssd1 vccd1 vccd1 _15290_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _14240_/A _14240_/B _14240_/C vssd1 vssd1 vccd1 vccd1 _14250_/B sky130_fd_sc_hd__a21o_1
XFILLER_172_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11453_ _19544_/Q _12155_/A2 _12155_/B1 _19608_/Q vssd1 vssd1 vccd1 vccd1 _11453_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10404_ _12084_/A _20504_/Q _12081_/S0 _20536_/Q vssd1 vssd1 vccd1 vccd1 _10404_/X
+ sky130_fd_sc_hd__o22a_1
X_14172_ _14262_/A _14170_/Y _14171_/X _18763_/A1 vssd1 vssd1 vccd1 vccd1 _14172_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11384_ _11383_/X _11375_/X _11384_/S vssd1 vssd1 vccd1 vccd1 _11384_/X sky130_fd_sc_hd__mux2_2
XFILLER_3_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123_ _20974_/Q _13272_/B _13122_/Y _18767_/A vssd1 vssd1 vccd1 vccd1 _13124_/B
+ sky130_fd_sc_hd__a211o_1
X_10335_ _10332_/X _10333_/X _10334_/X _12504_/B _10516_/S vssd1 vssd1 vccd1 vccd1
+ _10335_/X sky130_fd_sc_hd__a221o_1
XFILLER_98_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18980_ _18980_/A _18980_/B vssd1 vssd1 vccd1 vccd1 _21011_/D sky130_fd_sc_hd__nor2_1
XFILLER_180_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout2000 _17998_/A vssd1 vssd1 vccd1 vccd1 _17012_/C1 sky130_fd_sc_hd__buf_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _20951_/Q _20885_/Q vssd1 vssd1 vccd1 vccd1 _13064_/C sky130_fd_sc_hd__or2_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _20700_/Q _17931_/A1 _17946_/S vssd1 vssd1 vccd1 vccd1 _20700_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10266_ _11021_/A _20508_/Q _11035_/S _20540_/Q vssd1 vssd1 vccd1 vccd1 _10266_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_239_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1310 _14837_/S vssd1 vssd1 vccd1 vccd1 _14882_/B sky130_fd_sc_hd__clkbuf_8
X_12005_ _19650_/Q _19956_/Q _19294_/Q _20081_/Q _10622_/S _09834_/C vssd1 vssd1 vccd1
+ vccd1 _12005_/X sky130_fd_sc_hd__mux4_1
XFILLER_267_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1321 _15500_/A0 vssd1 vssd1 vccd1 vccd1 _16058_/A2 sky130_fd_sc_hd__clkbuf_4
X_17862_ _20635_/Q _10474_/X _17883_/S vssd1 vssd1 vccd1 vccd1 _20635_/D sky130_fd_sc_hd__mux2_1
Xfanout1332 _12085_/A2 vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__buf_6
XFILLER_278_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1343 _17378_/A2 vssd1 vssd1 vccd1 vccd1 _17390_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10197_ _10197_/A _11411_/B vssd1 vssd1 vccd1 vccd1 _15549_/S sky130_fd_sc_hd__nand2_4
XFILLER_238_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1354 _16593_/A vssd1 vssd1 vccd1 vccd1 _16591_/A sky130_fd_sc_hd__clkbuf_4
X_19601_ _19603_/CLK _19601_/D vssd1 vssd1 vccd1 vccd1 _19601_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1365 _17320_/S vssd1 vssd1 vccd1 vccd1 _17329_/S sky130_fd_sc_hd__buf_4
XFILLER_267_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16813_ _16849_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16813_/Y sky130_fd_sc_hd__nor2_1
Xfanout1376 _11213_/B vssd1 vssd1 vccd1 vccd1 _11379_/B sky130_fd_sc_hd__buf_8
XFILLER_19_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17793_ _20570_/Q _17933_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20570_/D sky130_fd_sc_hd__mux2_1
Xfanout1387 _09736_/Y vssd1 vssd1 vccd1 vccd1 _11860_/B2 sky130_fd_sc_hd__buf_4
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1398 _12081_/S0 vssd1 vssd1 vccd1 vccd1 _11698_/B2 sky130_fd_sc_hd__buf_4
XFILLER_266_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19532_ _19620_/CLK _19532_/D vssd1 vssd1 vccd1 vccd1 _19532_/Q sky130_fd_sc_hd__dfxtp_2
X_16744_ _20399_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16744_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13956_ _19152_/Q _13863_/B _14004_/B1 _13955_/X _16193_/A vssd1 vssd1 vccd1 vccd1
+ _19152_/D sky130_fd_sc_hd__o221a_1
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19463_ _20638_/CLK _19463_/D vssd1 vssd1 vccd1 vccd1 _19463_/Q sky130_fd_sc_hd__dfxtp_1
X_12907_ _13106_/B _12907_/B vssd1 vssd1 vccd1 vccd1 _12908_/A sky130_fd_sc_hd__and2_1
X_16675_ _19930_/Q _17051_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19930_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13887_ _19105_/Q _14738_/B _13889_/B1 _19171_/Q _13887_/C1 vssd1 vssd1 vccd1 vccd1
+ _19105_/D sky130_fd_sc_hd__o221a_1
XFILLER_235_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18414_ _18414_/A _18414_/B vssd1 vssd1 vccd1 vccd1 _20861_/D sky130_fd_sc_hd__and2_1
XFILLER_146_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12838_ _19512_/Q _12857_/B vssd1 vssd1 vccd1 vccd1 _12839_/D sky130_fd_sc_hd__nor2_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ _15983_/A _15626_/B vssd1 vssd1 vccd1 vccd1 _15626_/Y sky130_fd_sc_hd__nand2_1
X_19394_ _20685_/CLK _19394_/D vssd1 vssd1 vccd1 vccd1 _19394_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18345_ _18496_/B _18349_/B vssd1 vssd1 vccd1 vccd1 _18345_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15557_ _15977_/A1 _12741_/Y _15556_/X vssd1 vssd1 vccd1 vccd1 _15557_/X sky130_fd_sc_hd__o21a_1
X_12769_ _12517_/B split6/A _12767_/A _12767_/B vssd1 vssd1 vccd1 vccd1 _12771_/D
+ sky130_fd_sc_hd__a211o_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_168_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21041_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14508_ _19286_/Q _17696_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19286_/D sky130_fd_sc_hd__mux2_1
X_18276_ _20809_/Q _18275_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18277_/B sky130_fd_sc_hd__mux2_1
X_15488_ _12578_/B _12754_/X _15589_/S vssd1 vssd1 vccd1 vccd1 _15488_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17227_ _20265_/Q _20264_/Q vssd1 vssd1 vccd1 vccd1 _17441_/C sky130_fd_sc_hd__nor2_2
Xinput20 core_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_4
Xinput31 core_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
X_14439_ _17441_/A _17442_/A _17457_/B vssd1 vssd1 vccd1 vccd1 _14443_/B sky130_fd_sc_hd__or3b_2
XFILLER_128_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput42 core_wb_error_i vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_2
Xinput53 dout0[19] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_2
Xinput64 dout0[29] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_2
X_17158_ _20124_/Q _17926_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20124_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput75 dout0[39] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput86 dout0[49] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput97 dout0[59] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16109_ _19579_/Q _16127_/A2 _16127_/B1 vssd1 vssd1 vccd1 vccd1 _16109_/X sky130_fd_sc_hd__o21a_1
X_17089_ _20059_/Q _17751_/A1 _17114_/S vssd1 vssd1 vccd1 vccd1 _20059_/D sky130_fd_sc_hd__mux2_1
X_09980_ _12144_/C1 _09969_/X _09972_/X _09979_/X _12152_/A1 vssd1 vssd1 vccd1 vccd1
+ _09980_/X sky130_fd_sc_hd__a311o_1
XFILLER_66_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20505_ _20669_/CLK _20505_/D vssd1 vssd1 vccd1 vccd1 _20505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20436_ _20491_/CLK _20436_/D vssd1 vssd1 vccd1 vccd1 _20436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20367_ _20463_/CLK _20367_/D vssd1 vssd1 vccd1 vccd1 _20367_/Q sky130_fd_sc_hd__dfxtp_1
X_10120_ _10032_/Y _10119_/Y _09638_/Y vssd1 vssd1 vccd1 vccd1 _10120_/X sky130_fd_sc_hd__a21o_1
X_20298_ _20300_/CLK _20298_/D vssd1 vssd1 vccd1 vccd1 _20298_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10051_ _11259_/S _10049_/X _10050_/X vssd1 vssd1 vccd1 vccd1 _10051_/X sky130_fd_sc_hd__o21a_1
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _13810_/A1 _13721_/B split9/A input225/X vssd1 vssd1 vccd1 vccd1 _13810_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14790_ _19142_/Q _14802_/A2 _14789_/X _14794_/C1 vssd1 vssd1 vccd1 vccd1 _19519_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ _13777_/A _13741_/B vssd1 vssd1 vccd1 vccd1 _13741_/Y sky130_fd_sc_hd__nand2_8
X_10953_ _12429_/A1 _10951_/X _10952_/X vssd1 vssd1 vccd1 vccd1 _10953_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_272_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16460_ _19769_/Q _17189_/A1 _16471_/S vssd1 vssd1 vccd1 vccd1 _19769_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13672_ _13718_/A _13670_/Y _13671_/Y _13655_/A vssd1 vssd1 vccd1 vccd1 _13674_/B
+ sky130_fd_sc_hd__a211o_4
X_10884_ _10884_/A _11322_/B vssd1 vssd1 vccd1 vccd1 _10885_/B sky130_fd_sc_hd__nor2_4
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12623_ _19522_/Q _12901_/B _19523_/Q vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__a21oi_1
XFILLER_71_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15411_ _10642_/B _10638_/B _12468_/X _15410_/X vssd1 vssd1 vccd1 vccd1 _15411_/X
+ sky130_fd_sc_hd__a22o_1
X_16391_ _19742_/Q _16394_/C _18064_/A vssd1 vssd1 vccd1 vccd1 _16391_/Y sky130_fd_sc_hd__a21oi_1
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15342_ input261/X _15341_/X _15452_/S vssd1 vssd1 vccd1 vccd1 _15342_/X sky130_fd_sc_hd__mux2_1
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18130_ _14119_/B _19104_/Q _18134_/A vssd1 vssd1 vccd1 vccd1 _18320_/A sky130_fd_sc_hd__mux2_4
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12554_ _12554_/A _12554_/B _12554_/C vssd1 vssd1 vccd1 vccd1 _12555_/B sky130_fd_sc_hd__or3_4
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11505_ _20477_/Q _20317_/Q _11527_/S vssd1 vssd1 vccd1 vccd1 _11505_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18061_ _20760_/Q _20759_/Q _18061_/C vssd1 vssd1 vccd1 vccd1 _18063_/B sky130_fd_sc_hd__and3_1
X_15273_ _20919_/Q _15337_/A2 _15272_/X vssd1 vssd1 vccd1 vccd1 _15273_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12485_ _12716_/B _12731_/B vssd1 vssd1 vccd1 vccd1 _12485_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17012_ _19992_/Q _17012_/A2 _17011_/Y _17012_/C1 vssd1 vssd1 vccd1 vccd1 _19992_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14224_ _14255_/A _16068_/B _14224_/C vssd1 vssd1 vccd1 vccd1 _14224_/X sky130_fd_sc_hd__or3_1
X_11436_ _11981_/C1 _11435_/X _11432_/X _12137_/C1 vssd1 vssd1 vccd1 vccd1 _11436_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14155_ _19218_/Q _14256_/A2 _14154_/X _18698_/A vssd1 vssd1 vccd1 vccd1 _19218_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11367_ _11367_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__or2_1
XFILLER_4_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13106_ _13106_/A _13106_/B _13106_/C _13106_/D vssd1 vssd1 vccd1 vccd1 _13106_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ _10316_/X _10317_/X _11256_/S vssd1 vssd1 vccd1 vccd1 _10318_/X sky130_fd_sc_hd__mux2_1
X_14086_ _19202_/Q _14104_/A2 _14085_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1 _19202_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_258_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18963_ _18679_/Y _18970_/A2 _18962_/X _18901_/S vssd1 vssd1 vccd1 vccd1 _18963_/X
+ sky130_fd_sc_hd__a22o_1
X_11298_ _19398_/Q _20557_/Q _11303_/S vssd1 vssd1 vccd1 vccd1 _11298_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17914_ _20685_/Q _17914_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20685_/D sky130_fd_sc_hd__mux2_1
X_13037_ _20959_/Q _20893_/Q vssd1 vssd1 vccd1 vccd1 _13290_/A sky130_fd_sc_hd__or2_2
X_10249_ _19677_/Q _20165_/Q _11042_/B vssd1 vssd1 vccd1 vccd1 _10249_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18894_ _19136_/Q _18976_/A2 _18767_/B vssd1 vssd1 vccd1 vccd1 _18894_/Y sky130_fd_sc_hd__a21oi_1
Xfanout1140 _17941_/A1 vssd1 vssd1 vccd1 vccd1 _17801_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1151 _17909_/A1 vssd1 vssd1 vccd1 vccd1 _17107_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17845_ _20620_/Q _17917_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20620_/D sky130_fd_sc_hd__mux2_1
XFILLER_227_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1162 _09573_/Y vssd1 vssd1 vccd1 vccd1 _12403_/B1 sky130_fd_sc_hd__buf_6
XFILLER_67_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1173 _14895_/Y vssd1 vssd1 vccd1 vccd1 _16009_/B sky130_fd_sc_hd__buf_6
Xfanout1184 _15977_/A1 vssd1 vssd1 vccd1 vccd1 _12578_/B sky130_fd_sc_hd__buf_6
Xfanout1195 _17290_/C vssd1 vssd1 vccd1 vccd1 _17269_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_254_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17776_ _20555_/Q _17916_/A1 _17776_/S vssd1 vssd1 vccd1 vccd1 _20555_/D sky130_fd_sc_hd__mux2_1
XFILLER_226_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14988_ _15012_/B _14988_/B vssd1 vssd1 vccd1 vccd1 _14988_/Y sky130_fd_sc_hd__nor2_1
XFILLER_240_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19515_ _21004_/CLK _19515_/D vssd1 vssd1 vccd1 vccd1 _19515_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16727_ input68/X _16799_/S vssd1 vssd1 vccd1 vccd1 _16727_/Y sky130_fd_sc_hd__nand2_1
XFILLER_223_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13939_ _19143_/Q _13946_/B1 _13906_/X _13230_/X vssd1 vssd1 vccd1 vccd1 _19143_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19446_ _20710_/CLK _19446_/D vssd1 vssd1 vccd1 vccd1 _19446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16658_ _19915_/Q _17870_/A1 _16666_/S vssd1 vssd1 vccd1 vccd1 _19915_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _16052_/B2 _13426_/A _15608_/X vssd1 vssd1 vccd1 vccd1 _15609_/X sky130_fd_sc_hd__a21o_1
XFILLER_222_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19377_ _20668_/CLK _19377_/D vssd1 vssd1 vccd1 vccd1 _19377_/Q sky130_fd_sc_hd__dfxtp_1
X_16589_ _16591_/A _16589_/B vssd1 vssd1 vccd1 vccd1 _19860_/D sky130_fd_sc_hd__or2_1
XFILLER_176_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18328_ _20819_/Q _18343_/B _18327_/Y _18694_/A vssd1 vssd1 vccd1 vccd1 _20819_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18259_ _18299_/A1 _14322_/B _18258_/Y vssd1 vssd1 vccd1 vccd1 _18526_/B sky130_fd_sc_hd__o21ai_4
XFILLER_175_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20221_ _20816_/CLK _20221_/D vssd1 vssd1 vccd1 vccd1 _20221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20152_ _20563_/CLK _20152_/D vssd1 vssd1 vccd1 vccd1 _20152_/Q sky130_fd_sc_hd__dfxtp_1
X_09963_ _09955_/X _09956_/X _11902_/S vssd1 vssd1 vccd1 vccd1 _09963_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20630_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20083_ _20662_/CLK _20083_/D vssd1 vssd1 vccd1 vccd1 _20083_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _19387_/Q _20678_/Q _12146_/S vssd1 vssd1 vccd1 vccd1 _09894_/X sky130_fd_sc_hd__mux2_1
XFILLER_246_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_507 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_518 _16278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20985_ _21017_/CLK _20985_/D vssd1 vssd1 vccd1 vccd1 _20985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_529 _19499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12270_ _20490_/Q _12272_/B2 _12270_/B1 vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__o21a_1
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ _15155_/S _11223_/B vssd1 vssd1 vccd1 vccd1 _15071_/S sky130_fd_sc_hd__and2b_2
X_20419_ _20683_/CLK _20419_/D vssd1 vssd1 vccd1 vccd1 _20419_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_150_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11152_ _09595_/Y _11151_/X _11146_/Y _15103_/A1 vssd1 vssd1 vccd1 vccd1 _11152_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10103_ _12084_/A _19314_/Q _12084_/C vssd1 vssd1 vccd1 vccd1 _10103_/X sky130_fd_sc_hd__or3_1
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11083_ _20627_/Q _20591_/Q _12316_/S vssd1 vssd1 vccd1 vccd1 _11083_/X sky130_fd_sc_hd__mux2_1
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15960_ _15960_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15960_/X sky130_fd_sc_hd__and2_1
XFILLER_89_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput210 localMemory_wb_adr_i[6] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput221 localMemory_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_hd__buf_12
XFILLER_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput232 localMemory_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_hd__buf_12
X_14911_ _12945_/A _13897_/A _14917_/A vssd1 vssd1 vccd1 vccd1 _14951_/A sky130_fd_sc_hd__mux2_2
X_10034_ _10032_/Y _10033_/Y _09638_/Y vssd1 vssd1 vccd1 vccd1 _10034_/X sky130_fd_sc_hd__a21o_1
XFILLER_191_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput243 localMemory_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_hd__buf_12
Xinput254 manufacturerID[10] vssd1 vssd1 vccd1 vccd1 _17269_/A sky130_fd_sc_hd__buf_2
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _13439_/C _15925_/B _16056_/B1 vssd1 vssd1 vccd1 vccd1 _15891_/X sky130_fd_sc_hd__a21o_1
Xinput265 partID[10] vssd1 vssd1 vccd1 vccd1 _17302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_264_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput276 partID[6] vssd1 vssd1 vccd1 vccd1 _17290_/A sky130_fd_sc_hd__buf_2
X_17630_ _20386_/Q _17941_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20386_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ _10016_/B _10641_/B _14882_/B vssd1 vssd1 vccd1 vccd1 _14842_/X sky130_fd_sc_hd__mux2_1
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17561_ _20321_/Q _17800_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20321_/D sky130_fd_sc_hd__mux2_1
X_11985_ _11917_/S _11984_/X _11983_/X _12151_/A1 vssd1 vssd1 vccd1 vccd1 _11985_/X
+ sky130_fd_sc_hd__a211o_1
X_14773_ _19511_/Q _14773_/B vssd1 vssd1 vccd1 vccd1 _14773_/X sky130_fd_sc_hd__or2_1
XFILLER_263_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19300_ _19697_/CLK _19300_/D vssd1 vssd1 vccd1 vccd1 _19300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16512_ _19819_/Q _17835_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19819_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10936_ _10937_/A _19901_/Q _11211_/S _20026_/Q vssd1 vssd1 vccd1 vccd1 _10936_/X
+ sky130_fd_sc_hd__o22a_1
X_13724_ _13776_/B1 _13762_/B _13723_/X vssd1 vssd1 vccd1 vccd1 _13725_/B sky130_fd_sc_hd__a21oi_4
X_17492_ _20281_/Q _17494_/B vssd1 vssd1 vccd1 vccd1 _17492_/Y sky130_fd_sc_hd__nand2_1
XFILLER_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19231_ _19232_/CLK _19231_/D vssd1 vssd1 vccd1 vccd1 _19231_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_177_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16443_ _18835_/A _16443_/B _16444_/B vssd1 vssd1 vccd1 vccd1 _19761_/D sky130_fd_sc_hd__nor3_1
X_10867_ _19870_/Q _19771_/Q _12352_/S vssd1 vssd1 vccd1 vccd1 _10867_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13655_ _13655_/A _13655_/B vssd1 vssd1 vccd1 vccd1 _13656_/B sky130_fd_sc_hd__nor2_8
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19162_ _20670_/CLK _19162_/D vssd1 vssd1 vccd1 vccd1 _19162_/Q sky130_fd_sc_hd__dfxtp_1
X_12606_ _19511_/Q _19510_/Q _12855_/B vssd1 vssd1 vccd1 vccd1 _12845_/A sky130_fd_sc_hd__and3_1
X_16374_ _16378_/C _16374_/B vssd1 vssd1 vccd1 vccd1 _19735_/D sky130_fd_sc_hd__nor2_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _13586_/A _13586_/B _13586_/C vssd1 vssd1 vccd1 vccd1 _13586_/X sky130_fd_sc_hd__or3_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10798_ _10799_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10798_/X sky130_fd_sc_hd__and2_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18113_ _20779_/Q _18111_/B _18112_/Y vssd1 vssd1 vccd1 vccd1 _20779_/D sky130_fd_sc_hd__o21a_1
XFILLER_185_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15325_ _15283_/A _15304_/Y _15457_/B1 vssd1 vssd1 vccd1 vccd1 _15325_/Y sky130_fd_sc_hd__a21oi_1
X_12537_ _20874_/Q _12549_/B _12537_/C vssd1 vssd1 vccd1 vccd1 _12552_/A sky130_fd_sc_hd__and3_2
X_19093_ _19620_/CLK _19093_/D vssd1 vssd1 vccd1 vccd1 _19093_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ _20753_/Q _18045_/C _20754_/Q vssd1 vssd1 vccd1 vccd1 _18046_/B sky130_fd_sc_hd__a21oi_1
XFILLER_157_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15256_ _15407_/S _15251_/X _15253_/X _15578_/S vssd1 vssd1 vccd1 vccd1 _15256_/X
+ sky130_fd_sc_hd__o211a_1
X_12468_ _14894_/A _12468_/B _12468_/C vssd1 vssd1 vccd1 vccd1 _12468_/X sky130_fd_sc_hd__or3_4
X_11419_ _20382_/Q _20446_/Q _12121_/S vssd1 vssd1 vccd1 vccd1 _11419_/X sky130_fd_sc_hd__mux2_1
X_14207_ _19503_/Q _14208_/B vssd1 vssd1 vccd1 vccd1 _14209_/A sky130_fd_sc_hd__or2_1
X_15187_ _15326_/A _15187_/B _15187_/C vssd1 vssd1 vccd1 vccd1 _15208_/A sky130_fd_sc_hd__or3_1
X_12399_ _12399_/A1 _12395_/X _12398_/X _12399_/C1 vssd1 vssd1 vccd1 vccd1 _12399_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14138_ _19496_/Q _14139_/B vssd1 vssd1 vccd1 vccd1 _14138_/Y sky130_fd_sc_hd__nor2_1
X_19995_ _20621_/CLK _19995_/D vssd1 vssd1 vccd1 vccd1 _19995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14069_ _14081_/A _14069_/B _14069_/C vssd1 vssd1 vccd1 vccd1 _14069_/X sky130_fd_sc_hd__or3_1
X_18946_ _18966_/A _18946_/B vssd1 vssd1 vccd1 vccd1 _21006_/D sky130_fd_sc_hd__nor2_1
XFILLER_101_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18877_ _18877_/A _18877_/B vssd1 vssd1 vccd1 vccd1 _20996_/D sky130_fd_sc_hd__nor2_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17828_ _20603_/Q _17866_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20603_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_255_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17759_ _20538_/Q _17899_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20538_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_183_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20261_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20770_ _20860_/CLK _20770_/D vssd1 vssd1 vccd1 vccd1 _20770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_112_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20017_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_222_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19429_ _20694_/CLK _19429_/D vssd1 vssd1 vccd1 vccd1 _19429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20204_ _20760_/CLK _20204_/D vssd1 vssd1 vccd1 vccd1 _20204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout900 _15388_/S vssd1 vssd1 vccd1 vccd1 _15996_/B1 sky130_fd_sc_hd__buf_6
Xfanout911 _16046_/A1 vssd1 vssd1 vccd1 vccd1 _16017_/C1 sky130_fd_sc_hd__buf_6
Xfanout1909 _18726_/A vssd1 vssd1 vccd1 vccd1 _14776_/C1 sky130_fd_sc_hd__buf_4
Xfanout922 _14938_/Y vssd1 vssd1 vccd1 vccd1 _14983_/A sky130_fd_sc_hd__buf_6
X_20135_ _20641_/CLK _20135_/D vssd1 vssd1 vccd1 vccd1 _20135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09946_ _12366_/A1 _10033_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _09946_/X sky130_fd_sc_hd__a21o_4
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout933 _15039_/A vssd1 vssd1 vccd1 vccd1 _15061_/S sky130_fd_sc_hd__buf_6
Xfanout944 _15577_/S vssd1 vssd1 vccd1 vccd1 _15611_/S sky130_fd_sc_hd__buf_4
Xfanout955 _14262_/A vssd1 vssd1 vccd1 vccd1 _14325_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_246_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout966 _17687_/A1 vssd1 vssd1 vccd1 vccd1 _17930_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout977 _17866_/A1 vssd1 vssd1 vccd1 vccd1 _17691_/A1 sky130_fd_sc_hd__buf_2
X_20066_ _20472_/CLK _20066_/D vssd1 vssd1 vccd1 vccd1 _20066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _11977_/A1 _20710_/Q _11916_/S _09876_/X vssd1 vssd1 vccd1 vccd1 _09877_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout988 _17096_/A1 vssd1 vssd1 vccd1 vccd1 _17932_/A1 sky130_fd_sc_hd__buf_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout999 _16000_/A1 vssd1 vssd1 vccd1 vccd1 _15941_/B2 sky130_fd_sc_hd__buf_6
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_304 input231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 _17269_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_326 _13645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 _19495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_348 _17782_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11770_ _10801_/Y _11775_/B _10803_/Y vssd1 vssd1 vccd1 vccd1 _11771_/B sky130_fd_sc_hd__a21bo_1
XFILLER_246_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_359 _12295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20968_ _21040_/CLK _20968_/D vssd1 vssd1 vccd1 vccd1 _20968_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _19533_/Q _09613_/A _11225_/B _19597_/Q vssd1 vssd1 vccd1 vccd1 _10721_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20899_ _20998_/CLK _20899_/D vssd1 vssd1 vccd1 vccd1 _20899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13440_ _13440_/A _15954_/A _15981_/A vssd1 vssd1 vccd1 vccd1 _13440_/X sky130_fd_sc_hd__or3b_1
X_10652_ _19669_/Q _20157_/Q _12368_/S vssd1 vssd1 vccd1 vccd1 _10652_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13371_ _13368_/Y _13369_/X _13370_/Y _18671_/B vssd1 vssd1 vccd1 vccd1 _13371_/X
+ sky130_fd_sc_hd__o211a_1
X_10583_ _20634_/Q _20598_/Q _11676_/S vssd1 vssd1 vccd1 vccd1 _10583_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12322_ _20053_/Q _19928_/Q _12323_/S vssd1 vssd1 vccd1 vccd1 _12322_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15110_ _14844_/X _14854_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15110_/X sky130_fd_sc_hd__mux2_1
X_16090_ _10459_/X _16106_/A2 _16089_/X vssd1 vssd1 vccd1 vccd1 _19569_/D sky130_fd_sc_hd__o21a_1
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15041_ _15155_/S _15038_/X _15040_/X vssd1 vssd1 vccd1 vccd1 _15041_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_108_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12253_ _12337_/A _20522_/Q _12339_/S0 _20554_/Q vssd1 vssd1 vccd1 vccd1 _12253_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ _11202_/X _11203_/X _11204_/S vssd1 vssd1 vccd1 vccd1 _11204_/X sky130_fd_sc_hd__mux2_1
X_12184_ _19426_/Q _20585_/Q _12185_/S vssd1 vssd1 vccd1 vccd1 _12184_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18800_ _18480_/X _18819_/B _18798_/X _18799_/Y vssd1 vssd1 vccd1 vccd1 _18801_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11135_ _11138_/B vssd1 vssd1 vccd1 vccd1 _11136_/B sky130_fd_sc_hd__inv_2
X_19780_ _20557_/CLK _19780_/D vssd1 vssd1 vccd1 vccd1 _19780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16992_ _16950_/Y _16991_/X _16875_/B2 vssd1 vssd1 vccd1 vccd1 _16992_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18731_ _20966_/Q _18260_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18732_/B sky130_fd_sc_hd__mux2_1
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11066_ _19867_/Q _19768_/Q _11342_/S vssd1 vssd1 vccd1 vccd1 _11066_/X sky130_fd_sc_hd__mux2_1
X_15943_ _16000_/A1 _15932_/X _15933_/X _15942_/X vssd1 vssd1 vccd1 vccd1 _15943_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_283_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10017_ _13415_/A _11758_/B _10016_/Y vssd1 vssd1 vccd1 vccd1 _11761_/B sky130_fd_sc_hd__o21ai_2
XFILLER_276_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18662_ _20939_/Q _18686_/B vssd1 vssd1 vccd1 vccd1 _18662_/Y sky130_fd_sc_hd__nand2_1
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _20875_/Q _16018_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15874_/X sky130_fd_sc_hd__o21ba_1
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17613_ _20369_/Q _17647_/A1 _17623_/S vssd1 vssd1 vccd1 vccd1 _20369_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _14824_/X _14817_/X _15215_/S vssd1 vssd1 vccd1 vccd1 _14825_/X sky130_fd_sc_hd__mux2_1
XFILLER_252_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _12634_/A _18593_/A2 _18487_/X _18564_/A vssd1 vssd1 vccd1 vccd1 _18593_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17544_ _20304_/Q _17923_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20304_/D sky130_fd_sc_hd__mux2_1
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _19125_/Q _14764_/A2 _14755_/X _18476_/A vssd1 vssd1 vccd1 vccd1 _19502_/D
+ sky130_fd_sc_hd__o211a_1
X_11968_ _12051_/A1 _19361_/Q _20716_/Q _11978_/S _12051_/C1 vssd1 vssd1 vccd1 vccd1
+ _11968_/X sky130_fd_sc_hd__a221o_1
XFILLER_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13707_ _13707_/A _13742_/B vssd1 vssd1 vccd1 vccd1 _13747_/B sky130_fd_sc_hd__or2_2
XFILLER_220_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17475_ _17487_/A1 _17474_/Y _18048_/A vssd1 vssd1 vccd1 vccd1 _20272_/D sky130_fd_sc_hd__a21oi_1
X_10919_ _10914_/X _10918_/X _12310_/C1 vssd1 vssd1 vccd1 vccd1 _10919_/X sky130_fd_sc_hd__a21o_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11899_ _20143_/Q _20111_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _11899_/X sky130_fd_sc_hd__mux2_1
X_14687_ _19446_/Q _17936_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19446_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19214_ _19214_/CLK _19214_/D vssd1 vssd1 vccd1 vccd1 _19214_/Q sky130_fd_sc_hd__dfxtp_1
X_16426_ _19754_/Q _19755_/Q _16426_/C vssd1 vssd1 vccd1 vccd1 _16428_/B sky130_fd_sc_hd__and3_1
X_13638_ _15954_/A _13189_/B _16237_/B _13478_/B vssd1 vssd1 vccd1 vccd1 _13638_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_32_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19145_ _20291_/CLK _19145_/D vssd1 vssd1 vccd1 vccd1 _19145_/Q sky130_fd_sc_hd__dfxtp_1
X_16357_ _19729_/Q _16356_/B _18718_/A vssd1 vssd1 vccd1 vccd1 _16358_/B sky130_fd_sc_hd__o21ai_1
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13569_ _13142_/X _13566_/Y _13568_/Y _13624_/B2 vssd1 vssd1 vccd1 vccd1 _13569_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_145_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ _20888_/Q _15308_/B _15308_/C vssd1 vssd1 vccd1 vccd1 _15308_/X sky130_fd_sc_hd__and3_1
X_19076_ _20421_/Q vssd1 vssd1 vccd1 vccd1 _20421_/D sky130_fd_sc_hd__clkbuf_2
X_16288_ _19702_/Q _19703_/Q _19704_/Q vssd1 vssd1 vccd1 vccd1 _16290_/B sky130_fd_sc_hd__a21oi_1
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18027_ _20748_/Q _18030_/C vssd1 vssd1 vccd1 vccd1 _18028_/B sky130_fd_sc_hd__and2_1
X_15239_ _17284_/A _15482_/A2 _15232_/X _15238_/X vssd1 vssd1 vccd1 vccd1 _15239_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_246_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09800_ _20547_/Q _11665_/S vssd1 vssd1 vccd1 vccd1 _09800_/X sky130_fd_sc_hd__or2_1
XFILLER_87_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19978_ _19978_/CLK _19978_/D vssd1 vssd1 vccd1 vccd1 _19978_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09731_ _09731_/A _10979_/C vssd1 vssd1 vccd1 vccd1 _09731_/Y sky130_fd_sc_hd__nand2_2
X_18929_ _18659_/Y _18970_/A2 _18927_/Y _18928_/Y vssd1 vssd1 vccd1 vccd1 _18929_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09662_ _19695_/Q _19656_/Q vssd1 vssd1 vccd1 vccd1 _09662_/Y sky130_fd_sc_hd__nand2_2
XFILLER_227_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09593_ _09610_/A _09585_/A _19088_/Q _09592_/X vssd1 vssd1 vccd1 vccd1 _09593_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_282_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20822_ _20949_/CLK _20822_/D vssd1 vssd1 vccd1 vccd1 _20822_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20753_ _21020_/CLK _20753_/D vssd1 vssd1 vccd1 vccd1 _20753_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20684_ _20706_/CLK _20684_/D vssd1 vssd1 vccd1 vccd1 _20684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_80_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19603_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1706 _11537_/A1 vssd1 vssd1 vccd1 vccd1 _12100_/B1 sky130_fd_sc_hd__buf_6
Xfanout1717 _11309_/A1 vssd1 vssd1 vccd1 vccd1 _11375_/S sky130_fd_sc_hd__buf_8
XFILLER_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1728 _11258_/A1 vssd1 vssd1 vccd1 vccd1 _11008_/A1 sky130_fd_sc_hd__buf_6
Xfanout730 _18985_/X vssd1 vssd1 vccd1 vccd1 _19016_/B1 sky130_fd_sc_hd__buf_8
XFILLER_278_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout741 _14114_/X vssd1 vssd1 vccd1 vccd1 _14204_/A sky130_fd_sc_hd__buf_4
XFILLER_131_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1739 _12304_/C1 vssd1 vssd1 vccd1 vccd1 _11338_/A1 sky130_fd_sc_hd__buf_6
X_20118_ _20557_/CLK _20118_/D vssd1 vssd1 vccd1 vccd1 _20118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09929_ _09927_/X _09928_/X _11945_/S vssd1 vssd1 vccd1 vccd1 _09929_/X sky130_fd_sc_hd__mux2_1
Xfanout752 _18458_/X vssd1 vssd1 vccd1 vccd1 _18474_/S sky130_fd_sc_hd__buf_6
XFILLER_120_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout763 _18565_/Y vssd1 vssd1 vccd1 vccd1 _18619_/B sky130_fd_sc_hd__buf_6
XFILLER_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout774 _18902_/A vssd1 vssd1 vccd1 vccd1 _18671_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_258_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout785 _12911_/A vssd1 vssd1 vccd1 vccd1 _12906_/A sky130_fd_sc_hd__buf_8
XFILLER_246_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout796 _12488_/X vssd1 vssd1 vccd1 vccd1 _12652_/B sky130_fd_sc_hd__buf_8
X_12940_ _19256_/Q _12964_/A2 _16945_/B _20004_/Q vssd1 vssd1 vccd1 vccd1 _14921_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20049_ _20438_/CLK _20049_/D vssd1 vssd1 vccd1 vccd1 _20049_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12871_/A _12871_/B vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _12465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_112 _15303_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ _19374_/Q _17058_/A1 _14632_/S vssd1 vssd1 vccd1 vccd1 _19374_/D sky130_fd_sc_hd__mux2_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 _13676_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11812_/X _11814_/X _11821_/X _11904_/S _12137_/A1 vssd1 vssd1 vccd1 vccd1
+ _11822_/X sky130_fd_sc_hd__o221a_1
XANTENNA_134 _13683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _14895_/A _16063_/A2 _15589_/X vssd1 vssd1 vccd1 vccd1 _15591_/B sky130_fd_sc_hd__a21oi_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _13729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _13780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _19099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_178 _19115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14541_ _19311_/Q _17686_/A1 _14558_/S vssd1 vssd1 vccd1 vccd1 _19311_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _11772_/A _11405_/X _13425_/A _10645_/X vssd1 vssd1 vccd1 vccd1 _11754_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 _19172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _11118_/A _10703_/Y _10700_/Y _12431_/A1 vssd1 vssd1 vccd1 vccd1 _10704_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ input261/X _17275_/B vssd1 vssd1 vccd1 vccd1 _17260_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_202_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14472_ _18702_/A _14472_/B vssd1 vssd1 vccd1 vccd1 _19260_/D sky130_fd_sc_hd__and2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11684_/A1 _11683_/X _11680_/X _12072_/C1 vssd1 vssd1 vccd1 vccd1 _11684_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16211_ _19634_/Q _17095_/A1 _16227_/S vssd1 vssd1 vccd1 vccd1 _19634_/D sky130_fd_sc_hd__mux2_1
X_13423_ _13423_/A _13423_/B vssd1 vssd1 vccd1 vccd1 _13426_/B sky130_fd_sc_hd__xnor2_4
X_10635_ _12581_/A _15413_/A _10600_/Y vssd1 vssd1 vccd1 vccd1 _10638_/B sky130_fd_sc_hd__o21bai_4
X_17191_ _20155_/Q _17925_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20155_/D sky130_fd_sc_hd__mux2_1
XFILLER_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16142_ _19595_/Q _15243_/X _16196_/S vssd1 vssd1 vccd1 vccd1 _16143_/B sky130_fd_sc_hd__mux2_1
X_13354_ _13354_/A _13354_/B vssd1 vssd1 vccd1 vccd1 _13354_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_155_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10566_ _20159_/Q _12044_/B vssd1 vssd1 vccd1 vccd1 _10566_/X sky130_fd_sc_hd__or2_1
XFILLER_155_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12305_ _12306_/A1 _12396_/A1 _19493_/Q _12302_/S vssd1 vssd1 vccd1 vccd1 _12305_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16073_ _16073_/A _16081_/B vssd1 vssd1 vccd1 vccd1 _16073_/Y sky130_fd_sc_hd__nand2_1
X_13285_ _19227_/Q _13450_/A _19228_/Q vssd1 vssd1 vccd1 vccd1 _13287_/A sky130_fd_sc_hd__a21oi_1
X_10497_ _19277_/Q _09688_/B _11274_/B2 vssd1 vssd1 vccd1 vccd1 _10497_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _19652_/Q _12316_/S _12213_/X _12241_/S vssd1 vssd1 vccd1 vccd1 _12236_/X
+ sky130_fd_sc_hd__o211a_1
X_19901_ _20690_/CLK _19901_/D vssd1 vssd1 vccd1 vccd1 _19901_/Q sky130_fd_sc_hd__dfxtp_1
X_15024_ _12468_/B _12468_/C _14897_/A vssd1 vssd1 vccd1 vccd1 _15096_/B sky130_fd_sc_hd__o21ai_4
XFILLER_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19832_ _20621_/CLK _19832_/D vssd1 vssd1 vccd1 vccd1 _19832_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_268_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12167_ _11849_/S _12164_/X _12166_/X _12183_/C1 vssd1 vssd1 vccd1 vccd1 _12167_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11118_ _11118_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11118_/Y sky130_fd_sc_hd__nor2_1
X_19763_ _20268_/CLK _19763_/D vssd1 vssd1 vccd1 vccd1 _19763_/Q sky130_fd_sc_hd__dfxtp_2
X_16975_ input62/X input97/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16975_/X sky130_fd_sc_hd__mux2_8
X_12098_ _12102_/A1 _19488_/Q _19456_/Q _12097_/S _12100_/B1 vssd1 vssd1 vccd1 vccd1
+ _12098_/X sky130_fd_sc_hd__a221o_1
XFILLER_283_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18714_ _18714_/A _18714_/B vssd1 vssd1 vccd1 vccd1 _20957_/D sky130_fd_sc_hd__and2_1
XFILLER_77_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ _09750_/Y _11048_/X _11049_/B1 _12277_/A1 vssd1 vssd1 vccd1 vccd1 _12658_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_15926_ _12290_/C _12290_/D _16028_/C vssd1 vssd1 vccd1 vccd1 _15926_/Y sky130_fd_sc_hd__o21ai_1
X_19694_ _20704_/CLK _19694_/D vssd1 vssd1 vccd1 vccd1 _19694_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 coreIndex[6] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18645_ _18643_/Y _18644_/X _18966_/A vssd1 vssd1 vccd1 vccd1 _20934_/D sky130_fd_sc_hd__a21oi_1
XFILLER_92_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _20970_/Q _16045_/A2 _16016_/S _20842_/Q _15856_/X vssd1 vssd1 vccd1 vccd1
+ _15857_/X sky130_fd_sc_hd__a221o_1
XFILLER_37_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14808_ _14808_/A _15096_/A vssd1 vssd1 vccd1 vccd1 _14808_/Y sky130_fd_sc_hd__nand2_2
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18576_ _18783_/A _18576_/B vssd1 vssd1 vccd1 vccd1 _20916_/D sky130_fd_sc_hd__nor2_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _19548_/Q _15980_/A2 _15787_/X _16191_/A vssd1 vssd1 vccd1 vccd1 _19548_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17527_ _20249_/Q _20248_/Q vssd1 vssd1 vccd1 vccd1 _17528_/C sky130_fd_sc_hd__nor2_1
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14739_ _19494_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14739_/X sky130_fd_sc_hd__or2_1
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17458_ _17446_/A _17443_/D _17454_/D _17438_/B vssd1 vssd1 vccd1 vccd1 _17458_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16409_ _19748_/Q _16410_/C _19749_/Q vssd1 vssd1 vccd1 vccd1 _16411_/B sky130_fd_sc_hd__a21oi_1
XFILLER_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ _20243_/Q _17401_/A2 _17388_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _20243_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19128_ _19505_/CLK _19128_/D vssd1 vssd1 vccd1 vccd1 _19128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19059_ _20404_/Q vssd1 vssd1 vccd1 vccd1 _20404_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_146_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput300 _13787_/X vssd1 vssd1 vccd1 vccd1 addr1[6] sky130_fd_sc_hd__buf_4
XFILLER_133_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput311 _13618_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[15] sky130_fd_sc_hd__buf_4
Xoutput322 _13628_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[25] sky130_fd_sc_hd__buf_4
Xoutput333 _13191_/X vssd1 vssd1 vccd1 vccd1 core_wb_cyc_o sky130_fd_sc_hd__buf_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput344 _13721_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[19] sky130_fd_sc_hd__buf_4
Xoutput355 _13770_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[29] sky130_fd_sc_hd__buf_4
XFILLER_273_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21021_ _21021_/CLK _21021_/D vssd1 vssd1 vccd1 vccd1 _21021_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput366 _13632_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[0] sky130_fd_sc_hd__buf_4
Xoutput377 _13801_/X vssd1 vssd1 vccd1 vccd1 din0[10] sky130_fd_sc_hd__buf_4
Xoutput388 _13811_/X vssd1 vssd1 vccd1 vccd1 din0[20] sky130_fd_sc_hd__buf_4
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput399 _13821_/X vssd1 vssd1 vccd1 vccd1 din0[30] sky130_fd_sc_hd__buf_4
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09714_ _19389_/Q _20680_/Q _12124_/S vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_262_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09645_ _10373_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _10553_/B sky130_fd_sc_hd__nand2_8
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09576_ _09609_/A _12967_/B _19096_/Q _19098_/Q vssd1 vssd1 vccd1 vccd1 _09576_/X
+ sky130_fd_sc_hd__or4bb_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20805_ _21029_/CLK _20805_/D vssd1 vssd1 vccd1 vccd1 _20805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20736_ _20860_/CLK _20736_/D vssd1 vssd1 vccd1 vccd1 _20736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20667_ _20667_/CLK _20667_/D vssd1 vssd1 vccd1 vccd1 _20667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10420_ _19673_/Q _20161_/Q _10428_/S vssd1 vssd1 vccd1 vccd1 _10420_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20598_ _20698_/CLK _20598_/D vssd1 vssd1 vccd1 vccd1 _20598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10351_ _19380_/Q _12085_/A2 _10349_/X _11291_/B2 _10350_/X vssd1 vssd1 vccd1 vccd1
+ _10351_/X sky130_fd_sc_hd__o221a_1
XFILLER_125_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ _13453_/A _13453_/C _13453_/B vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__a21boi_4
XFILLER_279_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10282_ _09672_/A _09664_/B _10281_/X _11228_/B1 _19845_/Q vssd1 vssd1 vccd1 vccd1
+ _10282_/X sky130_fd_sc_hd__o32a_1
XFILLER_183_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12021_ _19689_/Q _20177_/Q _12025_/S vssd1 vssd1 vccd1 vccd1 _12021_/X sky130_fd_sc_hd__mux2_1
XFILLER_279_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1503 _09628_/Y vssd1 vssd1 vccd1 vccd1 _12041_/B sky130_fd_sc_hd__buf_8
XFILLER_238_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1514 _12149_/S vssd1 vssd1 vccd1 vccd1 _12133_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_215_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20482_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1525 _11682_/S vssd1 vssd1 vccd1 vccd1 _11994_/S sky130_fd_sc_hd__buf_6
Xfanout1536 _10303_/S vssd1 vssd1 vccd1 vccd1 _10485_/S sky130_fd_sc_hd__clkbuf_8
Xfanout1547 fanout1556/X vssd1 vssd1 vccd1 vccd1 _12375_/S sky130_fd_sc_hd__buf_6
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout560 _16666_/S vssd1 vssd1 vccd1 vccd1 _16668_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1558 _11358_/S vssd1 vssd1 vccd1 vccd1 _12300_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_219_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout571 _16490_/X vssd1 vssd1 vccd1 vccd1 _16521_/S sky130_fd_sc_hd__buf_8
Xfanout1569 _09625_/Y vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_120_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout582 _16199_/X vssd1 vssd1 vccd1 vccd1 _16231_/S sky130_fd_sc_hd__buf_12
X_16760_ _16760_/A vssd1 vssd1 vccd1 vccd1 _16760_/Y sky130_fd_sc_hd__clkinv_4
Xfanout593 _14719_/S vssd1 vssd1 vccd1 vccd1 _14736_/S sky130_fd_sc_hd__buf_12
X_13972_ _14002_/A1 _13978_/A2 _11231_/X _14002_/B1 _19839_/Q vssd1 vssd1 vccd1 vccd1
+ _14061_/C sky130_fd_sc_hd__o32a_1
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15711_ _14843_/S _15498_/Y _15499_/X _15258_/A vssd1 vssd1 vccd1 vccd1 _15711_/X
+ sky130_fd_sc_hd__o22a_2
X_12923_ _17526_/C _17522_/B vssd1 vssd1 vccd1 vccd1 _17461_/A sky130_fd_sc_hd__or2_4
X_16691_ _19946_/Q _17869_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19946_/D sky130_fd_sc_hd__mux2_1
XFILLER_280_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18430_ _18730_/A _18430_/B vssd1 vssd1 vccd1 vccd1 _20869_/D sky130_fd_sc_hd__and2_1
XFILLER_234_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15642_ _19718_/Q _15933_/B _15641_/X vssd1 vssd1 vccd1 vccd1 _15642_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _15649_/A1 _12832_/B _13350_/A _12710_/B vssd1 vssd1 vccd1 vccd1 _12860_/A
+ sky130_fd_sc_hd__o211a_2
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _19551_/Q _12155_/A2 _12155_/B1 _19615_/Q vssd1 vssd1 vccd1 vccd1 _11805_/X
+ sky130_fd_sc_hd__a22o_1
X_18361_ _18520_/B _18363_/B vssd1 vssd1 vccd1 vccd1 _18361_/Y sky130_fd_sc_hd__nand2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _19716_/Q _15395_/S _15572_/X vssd1 vssd1 vccd1 vccd1 _15573_/X sky130_fd_sc_hd__o21a_1
XFILLER_215_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _12783_/X _12784_/Y _12716_/B vssd1 vssd1 vccd1 vccd1 _12785_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_15_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17312_ _20209_/Q _17321_/A2 _17305_/C _17311_/X _17330_/C1 vssd1 vssd1 vccd1 vccd1
+ _17312_/X sky130_fd_sc_hd__a221o_1
XFILLER_199_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14524_ _14524_/A1 _14523_/X _14524_/B1 vssd1 vssd1 vccd1 vccd1 _14524_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18292_ _18746_/A _18292_/B vssd1 vssd1 vccd1 vccd1 _20812_/D sky130_fd_sc_hd__and2_1
X_11736_ _13420_/A _11794_/B _11734_/Y vssd1 vssd1 vccd1 vccd1 _11736_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17243_ _20186_/Q _17235_/Y _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17243_/X sky130_fd_sc_hd__a21o_1
X_14455_ _20223_/Q _19252_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14456_/B sky130_fd_sc_hd__mux2_1
XFILLER_159_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11667_ _11657_/X _11659_/X _11666_/X _11670_/S _12136_/B1 vssd1 vssd1 vccd1 vccd1
+ _11667_/X sky130_fd_sc_hd__o221a_1
X_13406_ _13033_/X _13034_/Y _13073_/Y vssd1 vssd1 vccd1 vccd1 _13406_/Y sky130_fd_sc_hd__a21oi_1
X_10618_ _20470_/Q _20310_/Q _10622_/S vssd1 vssd1 vccd1 vccd1 _10618_/X sky130_fd_sc_hd__mux2_1
X_17174_ _20140_/Q _17942_/A1 _17178_/S vssd1 vssd1 vccd1 vccd1 _20140_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14386_ _14386_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _14386_/X sky130_fd_sc_hd__xor2_1
X_11598_ _20416_/Q _11965_/B _11584_/X _11917_/S vssd1 vssd1 vccd1 vccd1 _11598_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16125_ _19587_/Q _16131_/A2 _16129_/B1 vssd1 vssd1 vccd1 vccd1 _16125_/X sky130_fd_sc_hd__o21a_1
X_10549_ _10549_/A vssd1 vssd1 vccd1 vccd1 _10549_/Y sky130_fd_sc_hd__inv_2
X_13337_ _19232_/Q _13350_/C vssd1 vssd1 vccd1 vccd1 _13337_/X sky130_fd_sc_hd__xor2_1
XFILLER_182_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16056_ _13181_/B _15982_/C _16056_/B1 _16055_/X vssd1 vssd1 vccd1 vccd1 _16056_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13268_ _14110_/B _13390_/B _13266_/Y _13267_/Y vssd1 vssd1 vccd1 vccd1 _13268_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_131_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15007_ _17239_/A _14983_/A _14987_/B _15006_/X _14980_/X vssd1 vssd1 vccd1 vccd1
+ _15007_/X sky130_fd_sc_hd__o311a_1
XFILLER_29_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12219_ _20394_/Q _20458_/Q _12219_/S vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13199_ _13199_/A _13199_/B vssd1 vssd1 vccd1 vccd1 _13199_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_116_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19815_ _20646_/CLK _19815_/D vssd1 vssd1 vccd1 vccd1 _19815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19746_ _20861_/CLK _19746_/D vssd1 vssd1 vccd1 vccd1 _19746_/Q sky130_fd_sc_hd__dfxtp_1
X_16958_ _16974_/A1 _16957_/X _16982_/B1 vssd1 vssd1 vccd1 vccd1 _16958_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_244_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15909_ _21038_/Q _21006_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _15909_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19677_ _20702_/CLK _19677_/D vssd1 vssd1 vccd1 vccd1 _19677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16889_ _20414_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16889_/X sky130_fd_sc_hd__a21o_2
XFILLER_38_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18628_ _19510_/Q _18628_/B vssd1 vssd1 vccd1 vccd1 _18628_/Y sky130_fd_sc_hd__nand2_1
XFILLER_266_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18559_ _20913_/Q _18559_/B vssd1 vssd1 vccd1 vccd1 _18559_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20679_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_12 _15449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20521_ _20685_/CLK _20521_/D vssd1 vssd1 vccd1 vccd1 _20521_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_23 _16869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 _16021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_45 _16856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_56 _16993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 _18324_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 _09647_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20452_ _20712_/CLK _20452_/D vssd1 vssd1 vccd1 vccd1 _20452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_89 _11687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20383_ _20715_/CLK _20383_/D vssd1 vssd1 vccd1 vccd1 _20383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21004_ _21004_/CLK _21004_/D vssd1 vssd1 vccd1 vccd1 _21004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09628_ _11268_/A _10979_/C vssd1 vssd1 vccd1 vccd1 _09628_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ _12513_/A _12513_/B _12517_/B vssd1 vssd1 vccd1 vccd1 _09561_/D sky130_fd_sc_hd__or3b_1
XFILLER_270_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _15220_/A _12463_/B _09560_/X vssd1 vssd1 vccd1 vccd1 _12570_/X sky130_fd_sc_hd__a21o_1
XFILLER_197_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20719_ _20719_/CLK _20719_/D vssd1 vssd1 vccd1 vccd1 _20719_/Q sky130_fd_sc_hd__dfxtp_1
X_11521_ _19382_/Q _20673_/Q _12133_/S vssd1 vssd1 vccd1 vccd1 _11521_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ _12039_/A1 _10553_/D split7/A vssd1 vssd1 vccd1 vccd1 _11452_/X sky130_fd_sc_hd__a21o_4
XFILLER_183_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14240_ _14240_/A _14240_/B _14240_/C vssd1 vssd1 vccd1 vccd1 _14242_/B sky130_fd_sc_hd__and3_1
XFILLER_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10403_ _10260_/S _10402_/X _09839_/A vssd1 vssd1 vccd1 vccd1 _10403_/X sky130_fd_sc_hd__o21a_1
XFILLER_125_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14171_ _14233_/S _14171_/B vssd1 vssd1 vccd1 vccd1 _14171_/X sky130_fd_sc_hd__or2_1
XFILLER_109_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11383_ _11375_/S _11378_/X _11382_/X vssd1 vssd1 vccd1 vccd1 _11383_/X sky130_fd_sc_hd__o21a_1
XFILLER_178_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10334_ _10356_/A _19476_/Q _19444_/Q _10345_/S vssd1 vssd1 vccd1 vccd1 _10334_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13122_ _13272_/B _13122_/B vssd1 vssd1 vccd1 vccd1 _13122_/Y sky130_fd_sc_hd__nor2_1
Xfanout2001 fanout2002/X vssd1 vssd1 vccd1 vccd1 _17998_/A sky130_fd_sc_hd__buf_6
XFILLER_180_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13053_ _20952_/Q _20886_/Q vssd1 vssd1 vccd1 vccd1 _13064_/B sky130_fd_sc_hd__or2_1
X_17930_ _20699_/Q _17930_/A1 _17934_/S vssd1 vssd1 vccd1 vccd1 _20699_/D sky130_fd_sc_hd__mux2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _10263_/X _10264_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _10265_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1300 _14267_/B1 vssd1 vssd1 vccd1 vccd1 _14216_/B1 sky130_fd_sc_hd__clkbuf_16
X_12004_ _19825_/Q _12009_/A2 _12002_/X _11641_/S _12003_/X vssd1 vssd1 vccd1 vccd1
+ _12004_/X sky130_fd_sc_hd__o221a_1
XFILLER_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1311 _14836_/S vssd1 vssd1 vccd1 vccd1 _14837_/S sky130_fd_sc_hd__buf_6
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17861_ _20634_/Q _17861_/A1 _17878_/S vssd1 vssd1 vccd1 vccd1 _20634_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10196_ _10197_/A _11411_/B vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__or2_4
Xfanout1322 _12465_/X vssd1 vssd1 vccd1 vccd1 _15500_/A0 sky130_fd_sc_hd__buf_6
Xfanout1333 _09738_/Y vssd1 vssd1 vccd1 vccd1 _12085_/A2 sky130_fd_sc_hd__buf_8
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1344 _17230_/Y vssd1 vssd1 vccd1 vccd1 _17378_/A2 sky130_fd_sc_hd__buf_8
Xfanout1355 _16557_/A vssd1 vssd1 vccd1 vccd1 _16593_/A sky130_fd_sc_hd__clkbuf_4
X_19600_ _19603_/CLK _19600_/D vssd1 vssd1 vccd1 vccd1 _19600_/Q sky130_fd_sc_hd__dfxtp_1
X_16812_ _17008_/B1 _16808_/X _16811_/X _16875_/B2 vssd1 vssd1 vccd1 vccd1 _16813_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_93_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1366 _13839_/X vssd1 vssd1 vccd1 vccd1 _17320_/S sky130_fd_sc_hd__buf_4
XFILLER_254_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17792_ _20569_/Q _17932_/A1 _17794_/S vssd1 vssd1 vccd1 vccd1 _20569_/D sky130_fd_sc_hd__mux2_1
XFILLER_226_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1377 _11213_/B vssd1 vssd1 vccd1 vccd1 _11305_/B sky130_fd_sc_hd__buf_8
XFILLER_219_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1388 _12188_/S vssd1 vssd1 vccd1 vccd1 _12174_/S sky130_fd_sc_hd__buf_6
X_19531_ _19606_/CLK _19531_/D vssd1 vssd1 vccd1 vccd1 _19531_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1399 _10400_/S vssd1 vssd1 vccd1 vccd1 _10397_/S sky130_fd_sc_hd__buf_6
XFILLER_282_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16743_ _16869_/A _16743_/B vssd1 vssd1 vccd1 vccd1 _16743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13955_ _19184_/Q _14049_/C _14003_/S vssd1 vssd1 vccd1 vccd1 _13955_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19462_ _20704_/CLK _19462_/D vssd1 vssd1 vccd1 vccd1 _19462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12906_ _12906_/A _12906_/B vssd1 vssd1 vccd1 vccd1 _12907_/B sky130_fd_sc_hd__or2_1
X_16674_ _19929_/Q _17886_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19929_/D sky130_fd_sc_hd__mux2_1
XFILLER_59_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _19104_/Q _14738_/B _13889_/B1 _11281_/A _16189_/A vssd1 vssd1 vccd1 vccd1
+ _19104_/D sky130_fd_sc_hd__o221a_1
XFILLER_250_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18413_ _20861_/Q _18215_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18414_/B sky130_fd_sc_hd__mux2_1
XFILLER_222_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _11792_/X _16028_/C _15624_/X vssd1 vssd1 vccd1 vccd1 _15625_/Y sky130_fd_sc_hd__a21oi_1
X_19393_ _20698_/CLK _19393_/D vssd1 vssd1 vccd1 vccd1 _19393_/Q sky130_fd_sc_hd__dfxtp_1
X_12837_ _12833_/Y _12836_/X _15703_/B2 vssd1 vssd1 vccd1 vccd1 _12839_/C sky130_fd_sc_hd__a21oi_4
XFILLER_222_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18344_ _20827_/Q _18343_/B _18343_/Y _18710_/A vssd1 vssd1 vccd1 vccd1 _20827_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _15544_/X _15555_/X _12716_/B vssd1 vssd1 vccd1 vccd1 _15556_/X sky130_fd_sc_hd__a21o_1
XFILLER_203_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12767_/A _12767_/B _12517_/B split6/A vssd1 vssd1 vccd1 vccd1 _12771_/C
+ sky130_fd_sc_hd__o211ai_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _19285_/Q _17695_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19285_/D sky130_fd_sc_hd__mux2_1
X_18275_ _18535_/B vssd1 vssd1 vccd1 vccd1 _18275_/Y sky130_fd_sc_hd__inv_2
X_11719_ _19641_/Q _19947_/Q _19285_/Q _20072_/Q _10621_/S _09834_/C vssd1 vssd1 vccd1
+ vccd1 _11719_/X sky130_fd_sc_hd__mux4_1
X_15487_ _15644_/A1 _16833_/B _15473_/Y vssd1 vssd1 vccd1 vccd1 _15487_/Y sky130_fd_sc_hd__o21ai_1
X_12699_ _13501_/B _12699_/B _12699_/C _12678_/B vssd1 vssd1 vccd1 vccd1 _12701_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_238_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17226_ _17443_/A _17226_/B vssd1 vssd1 vccd1 vccd1 _17235_/A sky130_fd_sc_hd__nor2_8
X_14438_ _19246_/Q _14438_/A2 _14437_/X _14802_/C1 vssd1 vssd1 vccd1 vccd1 _19246_/D
+ sky130_fd_sc_hd__o211a_1
Xinput10 core_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_6
Xinput21 core_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_4
Xinput32 core_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_8
Xinput43 dout0[0] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
Xinput54 dout0[1] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17157_ _20123_/Q _17925_/A1 _17166_/S vssd1 vssd1 vccd1 vccd1 _20123_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14369_ _13205_/Y _14368_/X _14437_/B _14437_/A vssd1 vssd1 vccd1 vccd1 _14369_/X
+ sky130_fd_sc_hd__a211o_1
Xinput65 dout0[2] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_2
Xinput76 dout0[3] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_2
Xinput87 dout0[4] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_2
X_16108_ _10375_/X _16126_/A2 _16107_/X vssd1 vssd1 vccd1 vccd1 _19578_/D sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_137_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _19223_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput98 dout0[5] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_2
X_17088_ _20058_/Q _17890_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20058_/D sky130_fd_sc_hd__mux2_1
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16039_ _19733_/Q _16039_/B vssd1 vssd1 vccd1 vccd1 _16039_/X sky130_fd_sc_hd__or2_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19729_ _20990_/CLK _19729_/D vssd1 vssd1 vccd1 vccd1 _19729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20504_ _20668_/CLK _20504_/D vssd1 vssd1 vccd1 vccd1 _20504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20435_ _20467_/CLK _20435_/D vssd1 vssd1 vccd1 vccd1 _20435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20366_ _20694_/CLK _20366_/D vssd1 vssd1 vccd1 vccd1 _20366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20297_ _20300_/CLK _20297_/D vssd1 vssd1 vccd1 vccd1 _20297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10050_ _11273_/A1 _19346_/Q _20701_/Q _10485_/S _12519_/C vssd1 vssd1 vccd1 vccd1
+ _10050_/X sky130_fd_sc_hd__a221o_1
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13740_ _13740_/A _13740_/B vssd1 vssd1 vccd1 vccd1 _13741_/B sky130_fd_sc_hd__nand2_8
XFILLER_244_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10952_ _11021_/A _19466_/Q _19434_/Q _11211_/S _11212_/S vssd1 vssd1 vccd1 vccd1
+ _10952_/X sky130_fd_sc_hd__a221o_1
XFILLER_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ _13718_/A _13708_/B vssd1 vssd1 vccd1 vccd1 _13671_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10883_ _10884_/A _11322_/B vssd1 vssd1 vccd1 vccd1 _10885_/A sky130_fd_sc_hd__and2_4
XFILLER_231_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15410_ _12471_/X _12466_/Y _15410_/S vssd1 vssd1 vccd1 vccd1 _15410_/X sky130_fd_sc_hd__mux2_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ _12911_/A _12911_/B vssd1 vssd1 vccd1 vccd1 _12912_/A sky130_fd_sc_hd__nand2_1
X_16390_ _19741_/Q _16388_/B _16389_/Y vssd1 vssd1 vccd1 vccd1 _19741_/D sky130_fd_sc_hd__o21a_1
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15341_ _17293_/A _15482_/A2 _15334_/X _15340_/X vssd1 vssd1 vccd1 vccd1 _15341_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12553_ _12553_/A _12553_/B _12553_/C _12553_/D vssd1 vssd1 vccd1 vccd1 _12554_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18060_ _20759_/Q _18061_/C _20760_/Q vssd1 vssd1 vccd1 vccd1 _18062_/B sky130_fd_sc_hd__a21oi_1
X_11504_ _11514_/A1 _20705_/Q _11818_/B2 _11503_/X vssd1 vssd1 vccd1 vccd1 _11504_/X
+ sky130_fd_sc_hd__a31o_1
X_15272_ _20887_/Q _14971_/A _15323_/B _15271_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15272_/X sky130_fd_sc_hd__a221o_1
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ split8/X _12847_/A2 _15526_/A vssd1 vssd1 vccd1 vccd1 _12484_/X sky130_fd_sc_hd__a21o_2
X_17011_ _17008_/Y _17010_/Y _17011_/B1 vssd1 vssd1 vccd1 vccd1 _17011_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14223_ _13609_/A _14222_/X _13609_/Y vssd1 vssd1 vccd1 vccd1 _14224_/C sky130_fd_sc_hd__o21a_1
X_11435_ _11433_/X _11434_/X _12058_/S vssd1 vssd1 vccd1 vccd1 _11435_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11366_ _12245_/A1 _11397_/A2 _11365_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _13664_/A
+ sky130_fd_sc_hd__o211a_4
X_14154_ _14255_/A _14204_/B _14154_/C vssd1 vssd1 vccd1 vccd1 _14154_/X sky130_fd_sc_hd__or3_1
XFILLER_152_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ _19380_/Q _20671_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__mux2_1
X_13105_ _13001_/B _13104_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _13105_/X sky130_fd_sc_hd__a21o_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14085_ _14099_/A _14107_/B _14085_/C vssd1 vssd1 vccd1 vccd1 _14085_/X sky130_fd_sc_hd__or3_1
X_11297_ _11295_/X _11296_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11297_/X sky130_fd_sc_hd__mux2_1
X_18962_ _09490_/Y _18961_/X _18975_/A vssd1 vssd1 vccd1 vccd1 _18962_/X sky130_fd_sc_hd__mux2_2
XFILLER_152_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10248_ _20133_/Q _20101_/Q _11303_/S vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__mux2_1
X_17913_ _20684_/Q _17913_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20684_/D sky130_fd_sc_hd__mux2_1
X_13036_ _20960_/Q _20894_/Q vssd1 vssd1 vccd1 vccd1 _13382_/B sky130_fd_sc_hd__nand2_2
X_18893_ _18955_/A _18893_/B vssd1 vssd1 vccd1 vccd1 _18893_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1130 _17937_/A1 vssd1 vssd1 vccd1 vccd1 _17592_/A1 sky130_fd_sc_hd__buf_2
Xfanout1141 _09936_/A2 vssd1 vssd1 vccd1 vccd1 _17941_/A1 sky130_fd_sc_hd__buf_2
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17844_ _20619_/Q _17916_/A1 _17844_/S vssd1 vssd1 vccd1 vccd1 _20619_/D sky130_fd_sc_hd__mux2_1
XFILLER_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10179_ _10176_/X _10177_/X _10178_/X _12504_/B _12514_/C vssd1 vssd1 vccd1 vccd1
+ _10179_/X sky130_fd_sc_hd__a221o_1
Xfanout1152 _09687_/X vssd1 vssd1 vccd1 vccd1 _17909_/A1 sky130_fd_sc_hd__buf_6
Xfanout1163 _18811_/S vssd1 vssd1 vccd1 vccd1 _18901_/S sky130_fd_sc_hd__buf_8
Xfanout1174 _14808_/Y vssd1 vssd1 vccd1 vccd1 _15246_/A sky130_fd_sc_hd__buf_6
Xfanout1185 _15977_/A1 vssd1 vssd1 vccd1 vccd1 _15348_/B2 sky130_fd_sc_hd__buf_2
X_17775_ _20554_/Q _17881_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20554_/D sky130_fd_sc_hd__mux2_1
Xfanout1196 _17302_/C vssd1 vssd1 vccd1 vccd1 _17290_/C sky130_fd_sc_hd__buf_2
XFILLER_282_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14987_ _14987_/A _14987_/B vssd1 vssd1 vccd1 vccd1 _14987_/Y sky130_fd_sc_hd__nor2_1
XFILLER_208_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16726_ _19701_/Q _19696_/Q vssd1 vssd1 vccd1 vccd1 _16726_/X sky130_fd_sc_hd__and2_4
X_19514_ _20913_/CLK _19514_/D vssd1 vssd1 vccd1 vccd1 _19514_/Q sky130_fd_sc_hd__dfxtp_4
X_13938_ _19142_/Q _13946_/B1 _13906_/X _13240_/X vssd1 vssd1 vccd1 vccd1 _19142_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19445_ _20702_/CLK _19445_/D vssd1 vssd1 vccd1 vccd1 _19445_/Q sky130_fd_sc_hd__dfxtp_1
X_16657_ _19914_/Q _17903_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19914_/D sky130_fd_sc_hd__mux2_1
X_13869_ _13869_/A _13902_/B vssd1 vssd1 vccd1 vccd1 _13869_/Y sky130_fd_sc_hd__nand2_1
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15608_ _16052_/A1 _15594_/X _15607_/Y _15544_/A vssd1 vssd1 vccd1 vccd1 _15608_/X
+ sky130_fd_sc_hd__a31o_1
X_19376_ _20667_/CLK _19376_/D vssd1 vssd1 vccd1 vccd1 _19376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16588_ _19860_/Q _16592_/A2 _16592_/B1 input31/X vssd1 vssd1 vccd1 vccd1 _16589_/B
+ sky130_fd_sc_hd__o22a_1
X_18327_ _18463_/B _18341_/B vssd1 vssd1 vccd1 vccd1 _18327_/Y sky130_fd_sc_hd__nand2_1
XFILLER_148_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _19747_/Q _15604_/A2 _15538_/X _16048_/C1 vssd1 vssd1 vccd1 vccd1 _15539_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_231_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18258_ _19547_/Q _18308_/B vssd1 vssd1 vccd1 vccd1 _18258_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_191_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17209_ _20173_/Q _17943_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20173_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18189_ _18134_/A _14177_/B _18188_/Y vssd1 vssd1 vccd1 vccd1 _18483_/B sky130_fd_sc_hd__o21ai_4
XFILLER_200_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20220_ _20268_/CLK _20220_/D vssd1 vssd1 vccd1 vccd1 _20220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20151_ _20561_/CLK _20151_/D vssd1 vssd1 vccd1 vccd1 _20151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09962_ _09952_/X _09954_/X _09961_/X _11904_/S _12137_/A1 vssd1 vssd1 vccd1 vccd1
+ _09962_/X sky130_fd_sc_hd__o221a_1
XFILLER_89_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20082_ _20446_/CLK _20082_/D vssd1 vssd1 vccd1 vccd1 _20082_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _20418_/Q _12146_/S _09871_/X _12150_/S vssd1 vssd1 vccd1 vccd1 _09893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_281_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_273_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20657_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_508 input215/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ _21016_/CLK _20984_/D vssd1 vssd1 vccd1 vccd1 _20984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_519 _16278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11220_ _11189_/B _11219_/X _11189_/Y vssd1 vssd1 vccd1 vccd1 _11223_/B sky130_fd_sc_hd__a21oi_4
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20418_ _20421_/CLK _20418_/D vssd1 vssd1 vccd1 vccd1 _20418_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ _11246_/A1 _11147_/Y _11150_/X _11149_/X vssd1 vssd1 vccd1 vccd1 _11151_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20349_ _20641_/CLK _20349_/D vssd1 vssd1 vccd1 vccd1 _20349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10102_ _12084_/A _19909_/Q _10092_/S _20034_/Q vssd1 vssd1 vccd1 vccd1 _10102_/X
+ sky130_fd_sc_hd__o22a_1
X_11082_ _20527_/Q _12316_/S _11081_/X _12317_/S vssd1 vssd1 vccd1 vccd1 _11082_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput200 localMemory_wb_adr_i[19] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput211 localMemory_wb_adr_i[7] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__clkbuf_2
XFILLER_276_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910_ _14950_/A _14950_/B _14973_/A vssd1 vssd1 vccd1 vccd1 _14920_/A sky130_fd_sc_hd__or3_1
Xinput222 localMemory_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_hd__buf_12
X_10033_ _10033_/A _10465_/A vssd1 vssd1 vccd1 vccd1 _10033_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput233 localMemory_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_hd__buf_12
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _15890_/A _15890_/B _15890_/C vssd1 vssd1 vccd1 vccd1 _15893_/B sky130_fd_sc_hd__or3_1
XFILLER_248_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput244 localMemory_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_hd__buf_12
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput255 manufacturerID[1] vssd1 vssd1 vccd1 vccd1 _17242_/A sky130_fd_sc_hd__clkbuf_4
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput266 partID[11] vssd1 vssd1 vccd1 vccd1 _17305_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_264_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput277 partID[7] vssd1 vssd1 vccd1 vccd1 _17293_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14841_ _14825_/X _14840_/X _14841_/S vssd1 vssd1 vccd1 vccd1 _14841_/X sky130_fd_sc_hd__mux2_1
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _20320_/Q _17696_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20320_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ _19133_/Q _14774_/A2 _14771_/X _14772_/C1 vssd1 vssd1 vccd1 vccd1 _19510_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_217_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ _20652_/Q _20616_/Q _12124_/S vssd1 vssd1 vccd1 vccd1 _11984_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16511_ _19818_/Q _17872_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19818_/D sky130_fd_sc_hd__mux2_1
X_13723_ _13655_/A _13684_/Y _13651_/Y _13714_/S vssd1 vssd1 vccd1 vccd1 _13723_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10935_ _19498_/Q _10935_/B vssd1 vssd1 vccd1 vccd1 _10935_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17491_ _17495_/A1 _17490_/Y _18835_/A vssd1 vssd1 vccd1 vccd1 _20280_/D sky130_fd_sc_hd__a21oi_1
XFILLER_232_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19230_ _19695_/CLK _19230_/D vssd1 vssd1 vccd1 vccd1 _19230_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_231_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16442_ _19760_/Q _19761_/Q _16442_/C vssd1 vssd1 vccd1 vccd1 _16444_/B sky130_fd_sc_hd__and3_1
X_13654_ _13658_/A _13689_/C vssd1 vssd1 vccd1 vccd1 _13655_/B sky130_fd_sc_hd__or2_4
X_10866_ _10866_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10866_/Y sky130_fd_sc_hd__nor2_1
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19161_ _19577_/CLK _19161_/D vssd1 vssd1 vccd1 vccd1 _19161_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _19509_/Q _12718_/A vssd1 vssd1 vccd1 vccd1 _12855_/B sky130_fd_sc_hd__and2_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _19735_/Q _16372_/B _17963_/B1 vssd1 vssd1 vccd1 vccd1 _16374_/B sky130_fd_sc_hd__o21ai_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13586_/A _13586_/C _13586_/B vssd1 vssd1 vccd1 vccd1 _13585_/Y sky130_fd_sc_hd__o21ai_1
X_10797_ _15150_/C1 _15304_/A _10766_/Y vssd1 vssd1 vccd1 vccd1 _10803_/B sky130_fd_sc_hd__o21ba_2
XFILLER_157_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _18112_/A _18117_/C vssd1 vssd1 vccd1 vccd1 _18112_/Y sky130_fd_sc_hd__nor2_1
X_15324_ _15282_/A _16784_/B _15304_/Y vssd1 vssd1 vccd1 vccd1 _15324_/X sky130_fd_sc_hd__o21a_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19092_ _19620_/CLK _19092_/D vssd1 vssd1 vccd1 vccd1 _19092_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12536_ _20871_/Q _12549_/B _12536_/C vssd1 vssd1 vccd1 vccd1 _12551_/A sky130_fd_sc_hd__and3_1
XFILLER_8_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18043_ _20753_/Q _18045_/C _18042_/Y vssd1 vssd1 vccd1 vccd1 _20753_/D sky130_fd_sc_hd__o21a_1
XFILLER_185_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15255_ _15121_/Y _15254_/X _15545_/A vssd1 vssd1 vccd1 vccd1 _15255_/X sky130_fd_sc_hd__mux2_4
X_12467_ _14894_/A _12468_/B _12468_/C vssd1 vssd1 vccd1 vccd1 _12467_/Y sky130_fd_sc_hd__nor3_4
XFILLER_144_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14206_ _20275_/Q _14237_/A2 _14216_/B1 input246/X vssd1 vssd1 vccd1 vccd1 _14208_/B
+ sky130_fd_sc_hd__a22o_4
X_11418_ _20478_/Q _20318_/Q _12149_/S vssd1 vssd1 vccd1 vccd1 _11418_/X sky130_fd_sc_hd__mux2_1
X_15186_ _11786_/B _15127_/B _15185_/X _12579_/D vssd1 vssd1 vccd1 vccd1 _15187_/C
+ sky130_fd_sc_hd__o211a_1
X_12398_ _11094_/S _12397_/X _12396_/X _12398_/C1 vssd1 vssd1 vccd1 vccd1 _12398_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_99_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14137_ _19494_/Q _14123_/B _14131_/B _14129_/X vssd1 vssd1 vccd1 vccd1 _14141_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_4_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11349_ _20341_/Q _12295_/B vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__or2_1
X_19994_ _20621_/CLK _19994_/D vssd1 vssd1 vccd1 vccd1 _19994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14068_ _19193_/Q _14108_/A2 _14067_/X _16107_/B1 vssd1 vssd1 vccd1 vccd1 _19193_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18945_ _18544_/X _18964_/B _18943_/X _18944_/Y vssd1 vssd1 vccd1 vccd1 _18946_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13019_ _20969_/Q _20903_/Q vssd1 vssd1 vccd1 vccd1 _13258_/A sky130_fd_sc_hd__or2_2
X_18876_ _18514_/X _18937_/B _18874_/X _18875_/Y vssd1 vssd1 vccd1 vccd1 _18877_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_239_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17827_ _20602_/Q _17899_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20602_/D sky130_fd_sc_hd__mux2_1
XFILLER_255_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17758_ _20537_/Q _17898_/A1 _17772_/S vssd1 vssd1 vccd1 vccd1 _20537_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16709_ _16719_/A _16710_/A _16720_/D vssd1 vssd1 vccd1 vccd1 _16709_/X sky130_fd_sc_hd__or3_4
X_17689_ _20473_/Q _17689_/A1 _17706_/S vssd1 vssd1 vccd1 vccd1 _20473_/D sky130_fd_sc_hd__mux2_1
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19428_ _20719_/CLK _19428_/D vssd1 vssd1 vccd1 vccd1 _19428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19359_ _20714_/CLK _19359_/D vssd1 vssd1 vccd1 vccd1 _19359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_152_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21024_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20203_ _20760_/CLK _20203_/D vssd1 vssd1 vccd1 vccd1 _20203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout901 _15388_/S vssd1 vssd1 vccd1 vccd1 _15568_/B1 sky130_fd_sc_hd__clkbuf_16
X_20134_ _20573_/CLK _20134_/D vssd1 vssd1 vccd1 vccd1 _20134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09945_ _19579_/Q _09944_/X _11229_/S vssd1 vssd1 vccd1 vccd1 _10033_/A sky130_fd_sc_hd__mux2_2
Xfanout912 _15322_/B vssd1 vssd1 vccd1 vccd1 _16046_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout923 _15989_/B1 vssd1 vssd1 vccd1 vccd1 _15961_/B1 sky130_fd_sc_hd__buf_4
Xfanout934 _11282_/Y vssd1 vssd1 vccd1 vccd1 _15039_/A sky130_fd_sc_hd__buf_4
Xfanout945 _15545_/A vssd1 vssd1 vccd1 vccd1 _15577_/S sky130_fd_sc_hd__buf_6
XFILLER_131_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout956 _14120_/Y vssd1 vssd1 vccd1 vccd1 _14262_/A sky130_fd_sc_hd__buf_8
XFILLER_57_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20065_ _20669_/CLK _20065_/D vssd1 vssd1 vccd1 vccd1 _20065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout967 _17060_/A1 vssd1 vssd1 vccd1 vccd1 _17687_/A1 sky130_fd_sc_hd__buf_2
X_09876_ _11977_/A1 _12120_/A1 _19355_/Q _12129_/S vssd1 vssd1 vccd1 vccd1 _09876_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout978 _10294_/X vssd1 vssd1 vccd1 vccd1 _17866_/A1 sky130_fd_sc_hd__buf_6
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout989 _17898_/A1 vssd1 vssd1 vccd1 vccd1 _17096_/A1 sky130_fd_sc_hd__buf_4
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_305 input232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_316 _13783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_327 _13649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 _19495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_349 _17892_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20967_ _21040_/CLK _20967_/D vssd1 vssd1 vccd1 vccd1 _20967_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_54_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10720_ _10720_/A _10720_/B vssd1 vssd1 vccd1 vccd1 _13567_/A sky130_fd_sc_hd__nor2_8
XFILLER_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _21027_/CLK _20898_/D vssd1 vssd1 vccd1 vccd1 _20898_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_201_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10651_ _09503_/A _10650_/X _10649_/X vssd1 vssd1 vccd1 vccd1 _10651_/X sky130_fd_sc_hd__o21a_1
XFILLER_213_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _20966_/Q _13370_/B vssd1 vssd1 vccd1 vccd1 _13370_/Y sky130_fd_sc_hd__nand2_1
X_10582_ _12063_/C1 _10580_/X _10581_/X _11680_/C1 vssd1 vssd1 vccd1 vccd1 _10582_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_221_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12321_ _12309_/S _12320_/X _12319_/X _12399_/A1 vssd1 vssd1 vccd1 vccd1 _12321_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15040_ _15039_/A _14869_/X _15039_/Y _15167_/S vssd1 vssd1 vccd1 vccd1 _15040_/X
+ sky130_fd_sc_hd__a211o_1
X_12252_ _12250_/X _12251_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _12252_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11203_ _19663_/Q _20151_/Q _11203_/S vssd1 vssd1 vccd1 vccd1 _11203_/X sky130_fd_sc_hd__mux2_1
X_12183_ _11849_/S _12182_/X _12181_/X _12183_/C1 vssd1 vssd1 vccd1 vccd1 _12183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ _11189_/B _12668_/A _11103_/Y vssd1 vssd1 vccd1 vccd1 _11138_/B sky130_fd_sc_hd__a21o_2
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16991_ input64/X input100/X _17009_/S vssd1 vssd1 vccd1 vccd1 _16991_/X sky130_fd_sc_hd__mux2_8
XFILLER_122_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11065_ _20367_/Q _20431_/Q _12397_/S vssd1 vssd1 vccd1 vccd1 _11065_/X sky130_fd_sc_hd__mux2_1
X_18730_ _18730_/A _18730_/B vssd1 vssd1 vccd1 vccd1 _20965_/D sky130_fd_sc_hd__and2_1
XFILLER_122_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15942_ _19761_/Q _15942_/A2 _15941_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15942_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ _09939_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _10016_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_264_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ _18932_/A _18661_/B vssd1 vssd1 vccd1 vccd1 _20938_/D sky130_fd_sc_hd__nor2_1
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _20747_/Q _15934_/A2 _15934_/B1 _20779_/Q vssd1 vssd1 vccd1 vccd1 _15873_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ _20368_/Q _17923_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20368_/D sky130_fd_sc_hd__mux2_1
X_14824_ _14820_/X _14823_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _14824_/X sky130_fd_sc_hd__mux2_1
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18592_ _20921_/Q _18592_/B vssd1 vssd1 vccd1 vccd1 _18592_/Y sky130_fd_sc_hd__nand2_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17543_ _20303_/Q _17679_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20303_/D sky130_fd_sc_hd__mux2_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _19502_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14755_/X sky130_fd_sc_hd__or2_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _19425_/Q _20584_/Q _11978_/S vssd1 vssd1 vccd1 vccd1 _11967_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13706_ _13780_/A _13706_/B vssd1 vssd1 vccd1 vccd1 _13706_/X sky130_fd_sc_hd__and2_1
X_17474_ _20272_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17474_/Y sky130_fd_sc_hd__nand2_1
X_10918_ _09618_/A _20090_/Q _10983_/S _10916_/X _10917_/X vssd1 vssd1 vccd1 vccd1
+ _10918_/X sky130_fd_sc_hd__a311o_1
XFILLER_204_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14686_ _19445_/Q _17935_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19445_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11898_ _19687_/Q _20175_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19213_ _19704_/CLK _19213_/D vssd1 vssd1 vccd1 vccd1 _19213_/Q sky130_fd_sc_hd__dfxtp_1
X_16425_ _19754_/Q _16426_/C _19755_/Q vssd1 vssd1 vccd1 vccd1 _16427_/B sky130_fd_sc_hd__a21oi_1
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13637_ _13637_/A _14525_/B _13637_/C vssd1 vssd1 vccd1 vccd1 _16237_/B sky130_fd_sc_hd__and3_4
X_10849_ _19175_/Q _11367_/B vssd1 vssd1 vccd1 vccd1 _10849_/X sky130_fd_sc_hd__or2_1
XFILLER_60_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19144_ _19523_/CLK _19144_/D vssd1 vssd1 vccd1 vccd1 _19144_/Q sky130_fd_sc_hd__dfxtp_1
X_16356_ _19729_/Q _16356_/B vssd1 vssd1 vccd1 vccd1 _16362_/C sky130_fd_sc_hd__and2_2
XFILLER_157_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ _13568_/A vssd1 vssd1 vccd1 vccd1 _13568_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15307_ _19740_/Q _15453_/A2 _15306_/X _15396_/A1 _16048_/C1 vssd1 vssd1 vccd1 vccd1
+ _15307_/X sky130_fd_sc_hd__a221o_1
X_12519_ _12519_/A _12584_/B _12519_/C _12588_/B vssd1 vssd1 vccd1 vccd1 _12520_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_157_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19075_ _20420_/Q vssd1 vssd1 vccd1 vccd1 _20420_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16287_ _19702_/Q _19703_/Q _16286_/Y vssd1 vssd1 vccd1 vccd1 _19703_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13499_ _13499_/A _13499_/B vssd1 vssd1 vccd1 vccd1 _13499_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18026_ _20747_/Q _18022_/B _18025_/Y vssd1 vssd1 vccd1 vccd1 _20747_/D sky130_fd_sc_hd__o21a_1
X_15238_ _20790_/Q _15016_/A _15021_/X _15237_/X vssd1 vssd1 vccd1 vccd1 _15238_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_173_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_114_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15169_ _15168_/A _15166_/A _15357_/S vssd1 vssd1 vccd1 vccd1 _15175_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19977_ _20004_/CLK _19977_/D vssd1 vssd1 vccd1 vccd1 _19977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09730_ _09730_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09730_/Y sky130_fd_sc_hd__nor2_2
X_18928_ _19141_/Q _18976_/A2 _18767_/B vssd1 vssd1 vccd1 vccd1 _18928_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09661_ _09666_/B _09657_/X _11326_/A _09660_/X vssd1 vssd1 vccd1 vccd1 _09678_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_269_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18859_ _19131_/Q _12533_/B _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18859_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_283_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09592_ _09592_/A _09592_/B _09592_/C vssd1 vssd1 vccd1 vccd1 _09592_/X sky130_fd_sc_hd__and3_1
XFILLER_209_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20821_ _20982_/CLK _20821_/D vssd1 vssd1 vccd1 vccd1 _20821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20752_ _21020_/CLK _20752_/D vssd1 vssd1 vccd1 vccd1 _20752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20683_ _20683_/CLK _20683_/D vssd1 vssd1 vccd1 vccd1 _20683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1707 _09730_/A vssd1 vssd1 vccd1 vccd1 _11304_/S sky130_fd_sc_hd__buf_6
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1718 _09505_/Y vssd1 vssd1 vccd1 vccd1 _11309_/A1 sky130_fd_sc_hd__buf_8
XFILLER_172_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout720 _13775_/A vssd1 vssd1 vccd1 vccd1 _13624_/B2 sky130_fd_sc_hd__buf_6
X_20117_ _20720_/CLK _20117_/D vssd1 vssd1 vccd1 vccd1 _20117_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1729 _18765_/A vssd1 vssd1 vccd1 vccd1 _11258_/A1 sky130_fd_sc_hd__buf_6
Xfanout731 _18985_/X vssd1 vssd1 vccd1 vccd1 _19002_/B1 sky130_fd_sc_hd__buf_4
XFILLER_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09928_ _20139_/Q _20107_/Q _09928_/S vssd1 vssd1 vccd1 vccd1 _09928_/X sky130_fd_sc_hd__mux2_1
Xfanout742 _19017_/X vssd1 vssd1 vccd1 vccd1 _19048_/B1 sky130_fd_sc_hd__buf_6
Xfanout753 _18458_/X vssd1 vssd1 vccd1 vccd1 fanout753/X sky130_fd_sc_hd__clkbuf_4
XFILLER_213_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout764 _18565_/Y vssd1 vssd1 vccd1 vccd1 _18592_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_172_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout775 _18902_/A vssd1 vssd1 vccd1 vccd1 _18628_/B sky130_fd_sc_hd__buf_6
Xfanout786 _12628_/A vssd1 vssd1 vccd1 vccd1 _12911_/A sky130_fd_sc_hd__buf_4
X_20048_ _20669_/CLK _20048_/D vssd1 vssd1 vccd1 vccd1 _20048_/Q sky130_fd_sc_hd__dfxtp_1
X_09859_ _09861_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09859_/X sky130_fd_sc_hd__and2b_1
Xfanout797 _12487_/Y vssd1 vssd1 vccd1 vccd1 _13334_/A sky130_fd_sc_hd__buf_8
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12870_ _12822_/Y _13362_/B _12869_/Y vssd1 vssd1 vccd1 vccd1 _12871_/B sky130_fd_sc_hd__o21a_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 _12493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11819_/X _11820_/X _11902_/S vssd1 vssd1 vccd1 vccd1 _11821_/X sky130_fd_sc_hd__mux2_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 _15303_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_124 _13718_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _13683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _13729_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _13780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ _19310_/Q _17058_/A1 _14562_/S vssd1 vssd1 vccd1 vccd1 _19310_/D sky130_fd_sc_hd__mux2_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _19108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _13419_/A _11752_/B vssd1 vssd1 vccd1 vccd1 _11752_/X sky130_fd_sc_hd__xor2_2
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _19115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _12420_/B1 _10701_/X _10702_/X vssd1 vssd1 vccd1 vccd1 _10703_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_241_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _20231_/Q _19260_/Q _14477_/S vssd1 vssd1 vccd1 vccd1 _14472_/B sky130_fd_sc_hd__mux2_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11681_/X _11682_/X _11995_/S vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _19633_/Q _17896_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19633_/D sky130_fd_sc_hd__mux2_1
X_13422_ _13422_/A _13422_/B vssd1 vssd1 vccd1 vccd1 _13426_/A sky130_fd_sc_hd__xnor2_4
X_17190_ _20154_/Q _17647_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20154_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10634_ _12107_/A1 _17895_/A1 _10633_/X _11397_/B2 vssd1 vssd1 vccd1 vccd1 _15413_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_195_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16141_ _19594_/Q _16194_/S _16140_/Y _16195_/A vssd1 vssd1 vccd1 vccd1 _19594_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13353_ _13031_/Y _13353_/B vssd1 vssd1 vccd1 vccd1 _13354_/B sky130_fd_sc_hd__nand2b_1
X_10565_ _12056_/S _10563_/X _10564_/X vssd1 vssd1 vccd1 vccd1 _10565_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12304_ _19797_/Q _12295_/B _12303_/X _12304_/C1 vssd1 vssd1 vccd1 vccd1 _12304_/X
+ sky130_fd_sc_hd__o211a_1
X_16072_ _19560_/Q _16081_/B _16071_/Y _16087_/B1 vssd1 vssd1 vccd1 vccd1 _19560_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13284_ _19226_/Q _13449_/B vssd1 vssd1 vccd1 vccd1 _13450_/A sky130_fd_sc_hd__and2_2
X_10496_ _11281_/A _20064_/Q _11268_/C vssd1 vssd1 vccd1 vccd1 _10496_/X sky130_fd_sc_hd__and3_1
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19900_ _20660_/CLK _19900_/D vssd1 vssd1 vccd1 vccd1 _19900_/Q sky130_fd_sc_hd__dfxtp_1
X_15023_ _15644_/A1 _16708_/B _14896_/X vssd1 vssd1 vccd1 vccd1 _15023_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12235_ _12309_/S _12234_/X _12233_/X _12318_/A1 vssd1 vssd1 vccd1 vccd1 _12235_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_136_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19831_ _19978_/CLK _19831_/D vssd1 vssd1 vccd1 vccd1 _19831_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12166_ _12186_/S _12166_/B vssd1 vssd1 vccd1 vccd1 _12166_/X sky130_fd_sc_hd__or2_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11117_ _11115_/X _11116_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _11118_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19762_ _19970_/CLK _19762_/D vssd1 vssd1 vccd1 vccd1 _19762_/Q sky130_fd_sc_hd__dfxtp_1
X_16974_ _16974_/A1 _16973_/X _16982_/B1 vssd1 vssd1 vccd1 vccd1 _16974_/Y sky130_fd_sc_hd__o21ai_2
X_12097_ _19891_/Q _19792_/Q _12097_/S vssd1 vssd1 vccd1 vccd1 _12097_/X sky130_fd_sc_hd__mux2_1
X_18713_ _20957_/Q _18215_/Y _18719_/S vssd1 vssd1 vccd1 vccd1 _18714_/B sky130_fd_sc_hd__mux2_1
XFILLER_283_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11048_ _11201_/A _11030_/X _11038_/X _11047_/Y vssd1 vssd1 vccd1 vccd1 _11048_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15925_ _15949_/B _15925_/B vssd1 vssd1 vccd1 vccd1 _15925_/Y sky130_fd_sc_hd__nand2_1
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19693_ _20155_/CLK _19693_/D vssd1 vssd1 vccd1 vccd1 _19693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 coreIndex[7] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15856_ _20938_/Q _16044_/A2 _15855_/X vssd1 vssd1 vccd1 vccd1 _15856_/X sky130_fd_sc_hd__o21a_1
X_18644_ _19514_/Q _18902_/A _18526_/X _18684_/A2 vssd1 vssd1 vccd1 vccd1 _18644_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_225_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14807_ _15220_/A _15095_/B _14808_/A vssd1 vssd1 vccd1 vccd1 _14807_/X sky130_fd_sc_hd__and3_1
XFILLER_52_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18575_ _18467_/B _18621_/A2 _18573_/Y _18574_/Y vssd1 vssd1 vccd1 vccd1 _18576_/B
+ sky130_fd_sc_hd__o211a_1
X_15787_ _15787_/A _15787_/B _15980_/A2 vssd1 vssd1 vccd1 vccd1 _15787_/X sky130_fd_sc_hd__or3b_1
XFILLER_224_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _19244_/Q _19243_/Q _13114_/B vssd1 vssd1 vccd1 vccd1 _13104_/B sky130_fd_sc_hd__and3_1
XFILLER_229_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17526_ _20300_/Q _17526_/B _17526_/C _20299_/Q vssd1 vssd1 vccd1 vccd1 _17537_/A
+ sky130_fd_sc_hd__or4b_2
X_14738_ _19149_/Q _14738_/B vssd1 vssd1 vccd1 vccd1 _14738_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_233_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17457_ _17457_/A _17457_/B _17457_/C vssd1 vssd1 vccd1 vccd1 _17457_/X sky130_fd_sc_hd__and3_1
X_14669_ _17918_/A _16604_/B vssd1 vssd1 vccd1 vccd1 _14670_/C sky130_fd_sc_hd__nor2_1
XFILLER_221_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16408_ _19748_/Q _16410_/C _16407_/Y vssd1 vssd1 vccd1 vccd1 _19748_/D sky130_fd_sc_hd__o21a_1
XFILLER_177_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17388_ _20242_/Q _17337_/B _17530_/A2 _20291_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17388_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16339_ _18863_/A _16339_/B _16340_/B vssd1 vssd1 vccd1 vccd1 _19722_/D sky130_fd_sc_hd__nor3_1
X_19127_ _19506_/CLK _19127_/D vssd1 vssd1 vccd1 vccd1 _19127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19058_ _20403_/Q vssd1 vssd1 vccd1 vccd1 _20403_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_195_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput301 _13788_/X vssd1 vssd1 vccd1 vccd1 addr1[7] sky130_fd_sc_hd__buf_4
XFILLER_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput312 _13619_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[16] sky130_fd_sc_hd__buf_4
X_18009_ _20741_/Q _18011_/C _18008_/Y vssd1 vssd1 vccd1 vccd1 _20741_/D sky130_fd_sc_hd__o21a_1
XFILLER_127_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput323 _13629_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[26] sky130_fd_sc_hd__buf_4
XFILLER_145_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput334 _13643_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[0] sky130_fd_sc_hd__buf_4
Xoutput345 _13645_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[1] sky130_fd_sc_hd__buf_4
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21020_ _21020_/CLK _21020_/D vssd1 vssd1 vccd1 vccd1 _21020_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput356 _13647_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[2] sky130_fd_sc_hd__buf_4
Xoutput367 _13634_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[1] sky130_fd_sc_hd__buf_4
XFILLER_113_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput378 _13802_/X vssd1 vssd1 vccd1 vccd1 din0[11] sky130_fd_sc_hd__buf_4
XFILLER_102_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput389 _13812_/X vssd1 vssd1 vccd1 vccd1 din0[21] sky130_fd_sc_hd__buf_4
XFILLER_248_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09713_ _20420_/Q _11987_/S _09690_/X _11833_/C1 vssd1 vssd1 vccd1 vccd1 _09713_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09644_ _11234_/A _11235_/A vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__and2_4
XFILLER_228_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ _12967_/B _09592_/A vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__nor2_4
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20804_ _20962_/CLK _20804_/D vssd1 vssd1 vccd1 vccd1 _20804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20735_ _20796_/CLK _20735_/D vssd1 vssd1 vccd1 vccd1 _20735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20666_ _20666_/CLK _20666_/D vssd1 vssd1 vccd1 vccd1 _20666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20597_ _20633_/CLK _20597_/D vssd1 vssd1 vccd1 vccd1 _20597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10350_ _11290_/A _20671_/Q _11026_/C vssd1 vssd1 vccd1 vccd1 _10350_/X sky130_fd_sc_hd__or3_1
XFILLER_192_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10281_ input112/X input147/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10281_/X sky130_fd_sc_hd__mux2_8
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12020_ _09776_/S _12015_/Y _12019_/Y _12020_/C1 vssd1 vssd1 vccd1 vccd1 _12020_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1504 _11891_/B vssd1 vssd1 vccd1 vccd1 _11899_/S sky130_fd_sc_hd__buf_6
XFILLER_250_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1515 fanout1522/X vssd1 vssd1 vccd1 vccd1 _12149_/S sky130_fd_sc_hd__buf_6
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1526 _11665_/S vssd1 vssd1 vccd1 vccd1 _11682_/S sky130_fd_sc_hd__buf_6
XFILLER_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1537 _10303_/S vssd1 vssd1 vccd1 vccd1 _10324_/S sky130_fd_sc_hd__buf_6
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1548 fanout1556/X vssd1 vssd1 vccd1 vccd1 _12368_/S sky130_fd_sc_hd__buf_4
Xfanout550 _17083_/X vssd1 vssd1 vccd1 vccd1 _17115_/S sky130_fd_sc_hd__buf_12
XFILLER_265_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1559 fanout1566/X vssd1 vssd1 vccd1 vccd1 _11358_/S sky130_fd_sc_hd__buf_6
Xfanout561 _16639_/X vssd1 vssd1 vccd1 vccd1 _16666_/S sky130_fd_sc_hd__buf_6
XFILLER_265_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout572 _16456_/X vssd1 vssd1 vccd1 vccd1 _16485_/S sky130_fd_sc_hd__buf_12
XFILLER_247_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout583 _16199_/X vssd1 vssd1 vccd1 vccd1 _16230_/S sky130_fd_sc_hd__buf_6
XFILLER_219_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13971_ _19157_/Q _14004_/A2 _14004_/B1 _13970_/X _16165_/C1 vssd1 vssd1 vccd1 vccd1
+ _19157_/D sky130_fd_sc_hd__o221a_1
XFILLER_19_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout594 _14704_/X vssd1 vssd1 vccd1 vccd1 _14719_/S sky130_fd_sc_hd__buf_12
XFILLER_247_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15710_ _13418_/A _12565_/B _15709_/X vssd1 vssd1 vccd1 vccd1 _15710_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_246_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12922_ _20300_/Q _20299_/Q vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__or2_4
XFILLER_246_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16690_ _19945_/Q _17202_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19945_/D sky130_fd_sc_hd__mux2_1
XFILLER_207_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15641_ _19750_/Q _15942_/A2 _15640_/X _15999_/C1 vssd1 vssd1 vccd1 vccd1 _15641_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12853_ _12851_/Y _12853_/B vssd1 vssd1 vccd1 vccd1 _13332_/A sky130_fd_sc_hd__nand2b_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11804_ _11804_/A _11804_/B vssd1 vssd1 vccd1 vccd1 _11880_/A sky130_fd_sc_hd__nand2_2
X_18360_ _20835_/Q _18363_/B _18359_/Y _18728_/A vssd1 vssd1 vccd1 vccd1 _20835_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _19748_/Q _15604_/A2 _15571_/X _16048_/C1 vssd1 vssd1 vccd1 vccd1 _15572_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _15413_/A _12784_/B vssd1 vssd1 vccd1 vccd1 _12784_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ input2/X input268/X _17329_/S vssd1 vssd1 vccd1 vccd1 _17311_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14523_ _13631_/B _16068_/A _16133_/A vssd1 vssd1 vccd1 vccd1 _14523_/X sky130_fd_sc_hd__o21ba_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _20812_/Q _18290_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18292_/B sky130_fd_sc_hd__mux2_1
X_11735_ _11574_/A _11735_/B vssd1 vssd1 vccd1 vccd1 _11794_/B sky130_fd_sc_hd__nand2b_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17242_/A _17290_/B _17269_/C vssd1 vssd1 vccd1 vccd1 _17242_/X sky130_fd_sc_hd__and3_1
XFILLER_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14454_ _18694_/A _14454_/B vssd1 vssd1 vccd1 vccd1 _19251_/D sky130_fd_sc_hd__and2_1
XFILLER_175_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11666_ _11664_/X _11665_/X _12056_/S vssd1 vssd1 vccd1 vccd1 _11666_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13405_ _13401_/Y _13402_/X _13404_/X vssd1 vssd1 vccd1 vccd1 _13405_/X sky130_fd_sc_hd__a21o_1
X_17173_ _20139_/Q _17801_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20139_/D sky130_fd_sc_hd__mux2_1
X_10617_ _10608_/X _10616_/X _09839_/A vssd1 vssd1 vccd1 vccd1 _10617_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14385_ _14372_/Y _14376_/B _14374_/B vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__o21a_1
X_11597_ _11917_/S _11596_/X _11595_/X _11597_/C1 vssd1 vssd1 vccd1 vccd1 _11597_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_259_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16124_ _10380_/X _16132_/A2 _16123_/X vssd1 vssd1 vccd1 vccd1 _19586_/D sky130_fd_sc_hd__o21a_1
X_13336_ _19231_/Q _19230_/Q _13403_/B vssd1 vssd1 vccd1 vccd1 _13350_/C sky130_fd_sc_hd__and3_1
XFILLER_128_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10548_ _09643_/A _09636_/B _10020_/Y _10547_/Y _15103_/A1 vssd1 vssd1 vccd1 vccd1
+ _10549_/A sky130_fd_sc_hd__a2111o_2
XFILLER_155_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16055_ _12449_/X _12451_/Y _16028_/C vssd1 vssd1 vccd1 vccd1 _16055_/X sky130_fd_sc_hd__o21a_1
XFILLER_127_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13267_ _20935_/Q _13363_/B _18667_/B vssd1 vssd1 vccd1 vccd1 _13267_/Y sky130_fd_sc_hd__a21oi_1
X_10479_ _19408_/Q _20567_/Q _10485_/S vssd1 vssd1 vccd1 vccd1 _10479_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15006_ _15004_/X _15005_/X _14983_/Y _14986_/X vssd1 vssd1 vccd1 vccd1 _15006_/X
+ sky130_fd_sc_hd__a211o_1
X_12218_ _20490_/Q _20330_/Q _12381_/S vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13198_ _12871_/A _12871_/B _13199_/B vssd1 vssd1 vccd1 vccd1 _13233_/C sky130_fd_sc_hd__a21boi_1
XFILLER_124_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19814_ _20673_/CLK _19814_/D vssd1 vssd1 vccd1 vccd1 _19814_/Q sky130_fd_sc_hd__dfxtp_1
X_12149_ _19295_/Q _20082_/Q _12149_/S vssd1 vssd1 vccd1 vccd1 _12149_/X sky130_fd_sc_hd__mux2_1
XFILLER_284_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19745_ _20795_/CLK _19745_/D vssd1 vssd1 vccd1 vccd1 _19745_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16957_ _16981_/A1 _15882_/X _16945_/X _16956_/X vssd1 vssd1 vccd1 vccd1 _16957_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_77_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15908_ _20876_/Q _16018_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15908_/X sky130_fd_sc_hd__o21ba_1
X_19676_ _20315_/CLK _19676_/D vssd1 vssd1 vccd1 vccd1 _19676_/Q sky130_fd_sc_hd__dfxtp_1
X_16888_ _19977_/Q _16887_/A _16887_/Y _16896_/C1 vssd1 vssd1 vccd1 vccd1 _19977_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_264_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18627_ _20930_/Q _18686_/B vssd1 vssd1 vccd1 vccd1 _18627_/Y sky130_fd_sc_hd__nand2_1
XFILLER_280_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15839_ _15948_/A1 _12817_/X _15838_/X _15921_/B2 vssd1 vssd1 vccd1 vccd1 _15841_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_253_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_252_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18558_ _18973_/A _18558_/B vssd1 vssd1 vccd1 vccd1 _20912_/D sky130_fd_sc_hd__nor2_1
XFILLER_240_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17509_ _17525_/A1 _17508_/Y _18932_/A vssd1 vssd1 vccd1 vccd1 _20289_/D sky130_fd_sc_hd__a21oi_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18489_ _18598_/A _18489_/B vssd1 vssd1 vccd1 vccd1 _20889_/D sky130_fd_sc_hd__nor2_1
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 _15449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20520_ _20706_/CLK _20520_/D vssd1 vssd1 vccd1 vccd1 _20520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_24 _15632_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_35 _16021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_46 _16858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20720_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_57 _17003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20451_ _20451_/CLK _20451_/D vssd1 vssd1 vccd1 vccd1 _20451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_68 _18913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _09685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20382_ _20677_/CLK _20382_/D vssd1 vssd1 vccd1 vccd1 _20382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_273_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21003_ _21010_/CLK _21003_/D vssd1 vssd1 vccd1 vccd1 _21003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ _18765_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09627_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09558_ _12708_/A _12517_/B _09561_/C vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__or3_4
XFILLER_43_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09489_ _19525_/Q vssd1 vssd1 vccd1 vccd1 _14433_/A sky130_fd_sc_hd__inv_2
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11520_ _20413_/Q _12133_/S _11498_/X _09901_/S vssd1 vssd1 vccd1 vccd1 _11520_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20718_ _20718_/CLK _20718_/D vssd1 vssd1 vccd1 vccd1 _20718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ _11436_/X _11450_/X _12153_/A1 vssd1 vssd1 vccd1 vccd1 _11451_/X sky130_fd_sc_hd__a21o_1
XFILLER_183_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20649_ _20649_/CLK _20649_/D vssd1 vssd1 vccd1 vccd1 _20649_/Q sky130_fd_sc_hd__dfxtp_1
X_10402_ _10398_/X _10401_/X _10516_/S vssd1 vssd1 vccd1 vccd1 _10402_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14170_ _14170_/A _14170_/B vssd1 vssd1 vccd1 vccd1 _14170_/Y sky130_fd_sc_hd__xnor2_1
X_11382_ _11379_/X _11380_/X _11381_/X _12420_/B1 _12265_/A vssd1 vssd1 vccd1 vccd1
+ _11382_/X sky130_fd_sc_hd__a221o_1
XFILLER_178_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13121_ _13121_/A _13121_/B vssd1 vssd1 vccd1 vccd1 _13122_/B sky130_fd_sc_hd__xnor2_1
X_10333_ _19780_/Q _11305_/B _09730_/A vssd1 vssd1 vccd1 vccd1 _10333_/X sky130_fd_sc_hd__o21a_1
XFILLER_191_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13052_ _20952_/Q _20886_/Q vssd1 vssd1 vccd1 vccd1 _13064_/A sky130_fd_sc_hd__nand2_1
Xfanout2002 _16278_/A vssd1 vssd1 vccd1 vccd1 fanout2002/X sky130_fd_sc_hd__buf_8
XFILLER_140_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10264_ _19638_/Q _19944_/Q _19282_/Q _20069_/Q _11035_/S _11021_/C vssd1 vssd1 vccd1
+ vccd1 _10264_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12003_ _12003_/A _19329_/Q _12003_/C vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__or3_1
XFILLER_121_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1301 _14117_/Y vssd1 vssd1 vccd1 vccd1 _14267_/B1 sky130_fd_sc_hd__buf_8
X_17860_ _20633_/Q _17894_/A1 _17882_/S vssd1 vssd1 vccd1 vccd1 _20633_/D sky130_fd_sc_hd__mux2_1
Xfanout1312 _12474_/Y vssd1 vssd1 vccd1 vccd1 _14836_/S sky130_fd_sc_hd__buf_4
X_10195_ _19507_/Q _15528_/A _11398_/S vssd1 vssd1 vccd1 vccd1 _11411_/B sky130_fd_sc_hd__mux2_4
XFILLER_266_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1323 _12463_/B vssd1 vssd1 vccd1 vccd1 _16053_/A sky130_fd_sc_hd__buf_4
XFILLER_238_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1334 _11192_/A2 vssd1 vssd1 vccd1 vccd1 _11291_/A2 sky130_fd_sc_hd__buf_8
XFILLER_239_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1345 _17321_/A2 vssd1 vssd1 vccd1 vccd1 _17330_/A2 sky130_fd_sc_hd__buf_4
X_16811_ _16846_/A _09521_/Y _16809_/X _16810_/Y vssd1 vssd1 vccd1 vccd1 _16811_/X
+ sky130_fd_sc_hd__o211a_4
Xfanout1356 _16551_/A vssd1 vssd1 vccd1 vccd1 _16557_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_282_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1367 _14330_/A2 vssd1 vssd1 vccd1 vccd1 _14431_/A2 sky130_fd_sc_hd__buf_6
XFILLER_94_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17791_ _20568_/Q _17931_/A1 _17806_/S vssd1 vssd1 vccd1 vccd1 _20568_/D sky130_fd_sc_hd__mux2_1
Xfanout1378 _09737_/Y vssd1 vssd1 vccd1 vccd1 _11213_/B sky130_fd_sc_hd__buf_12
XFILLER_94_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1389 _11848_/S0 vssd1 vssd1 vccd1 vccd1 _12188_/S sky130_fd_sc_hd__buf_6
XFILLER_253_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19530_ _19620_/CLK _19530_/D vssd1 vssd1 vccd1 vccd1 _19530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13954_ _14002_/A1 _13960_/A2 _11059_/X _14002_/B1 _19833_/Q vssd1 vssd1 vccd1 vccd1
+ _14049_/C sky130_fd_sc_hd__o32a_1
X_16742_ _19962_/Q _16822_/A _16741_/Y _18801_/A vssd1 vssd1 vccd1 vccd1 _19962_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_143_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12905_ _12906_/A _12906_/B vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__nand2_2
X_19461_ _20155_/CLK _19461_/D vssd1 vssd1 vccd1 vccd1 _19461_/Q sky130_fd_sc_hd__dfxtp_1
X_16673_ _17919_/A _17574_/B _16673_/C vssd1 vssd1 vccd1 vccd1 _16673_/X sky130_fd_sc_hd__and3_4
XFILLER_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13885_ _19103_/Q _14738_/B _13889_/B1 _18765_/B _16189_/A vssd1 vssd1 vccd1 vccd1
+ _19103_/D sky130_fd_sc_hd__o221a_1
XFILLER_185_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18412_ _18416_/A _18412_/B vssd1 vssd1 vccd1 vccd1 _20860_/D sky130_fd_sc_hd__and2_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12836_ split8/X _12847_/A2 _15526_/A _12835_/Y vssd1 vssd1 vccd1 vccd1 _12836_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _13427_/C _15982_/C _16056_/B1 vssd1 vssd1 vccd1 vccd1 _15624_/X sky130_fd_sc_hd__a21o_1
XFILLER_222_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _20683_/CLK _19392_/D vssd1 vssd1 vccd1 vccd1 _19392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18343_ _18493_/B _18343_/B vssd1 vssd1 vccd1 vccd1 _18343_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _15552_/X _15554_/Y _15527_/B vssd1 vssd1 vccd1 vccd1 _15555_/X sky130_fd_sc_hd__a21o_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12767_/A _12767_/B vssd1 vssd1 vccd1 vccd1 _12767_/X sky130_fd_sc_hd__or2_1
XFILLER_187_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _19284_/Q _17903_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19284_/D sky130_fd_sc_hd__mux2_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18274_ _18299_/A1 _14352_/B _18273_/Y vssd1 vssd1 vccd1 vccd1 _18535_/B sky130_fd_sc_hd__o21ai_4
X_11718_ _11716_/X _11717_/X _11718_/S vssd1 vssd1 vccd1 vccd1 _11718_/X sky130_fd_sc_hd__mux2_1
X_15486_ _15021_/A _15475_/X _15485_/X vssd1 vssd1 vccd1 vccd1 _16833_/B sky130_fd_sc_hd__a21oi_4
XFILLER_203_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _12698_/A _12698_/B _12698_/C _12698_/D vssd1 vssd1 vccd1 vccd1 _12699_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_202_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17225_ _14123_/B _17219_/Y _17224_/X _18698_/A vssd1 vssd1 vccd1 vccd1 _20184_/D
+ sky130_fd_sc_hd__o211a_1
X_14437_ _14437_/A _14437_/B _14437_/C vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__or3_1
X_11649_ _19513_/Q _11648_/Y _11649_/S vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__mux2_4
Xinput11 core_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_4
Xinput22 core_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_4
XFILLER_156_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput33 core_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
X_17156_ _20122_/Q _17647_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20122_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput44 dout0[10] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_2
X_14368_ _14427_/A _14364_/B _14367_/Y _13205_/A vssd1 vssd1 vccd1 vccd1 _14368_/X
+ sky130_fd_sc_hd__a211o_1
Xinput55 dout0[20] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput66 dout0[30] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_2
Xinput77 dout0[40] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ _19578_/Q _16079_/B _16107_/B1 vssd1 vssd1 vccd1 vccd1 _16107_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput88 dout0[50] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_2
X_13319_ _13314_/Y _13318_/Y _14275_/A1 vssd1 vssd1 vccd1 vccd1 _13319_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17087_ _20057_/Q _17855_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20057_/D sky130_fd_sc_hd__mux2_1
Xinput99 dout0[60] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ _19512_/Q _14300_/B vssd1 vssd1 vccd1 vccd1 _14301_/A sky130_fd_sc_hd__nand2_1
XFILLER_115_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16038_ _19733_/Q _14933_/Y _14935_/Y _19765_/Q vssd1 vssd1 vccd1 vccd1 _16038_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_177_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19520_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_106_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20795_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_257_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17989_ _18080_/A _17989_/B vssd1 vssd1 vccd1 vccd1 _17989_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19728_ _19970_/CLK _19728_/D vssd1 vssd1 vccd1 vccd1 _19728_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1890 _13887_/C1 vssd1 vssd1 vccd1 vccd1 _17432_/A sky130_fd_sc_hd__buf_4
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19659_ _19695_/CLK _19659_/D vssd1 vssd1 vccd1 vccd1 _19659_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20503_ _20635_/CLK _20503_/D vssd1 vssd1 vccd1 vccd1 _20503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20434_ _20630_/CLK _20434_/D vssd1 vssd1 vccd1 vccd1 _20434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20365_ _21047_/A _20365_/D vssd1 vssd1 vccd1 vccd1 _20365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20296_ _20296_/CLK _20296_/D vssd1 vssd1 vccd1 vccd1 _20296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10951_ _19869_/Q _19770_/Q _11211_/S vssd1 vssd1 vccd1 vccd1 _10951_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13670_ _13670_/A1 _17895_/A1 _10595_/X _13684_/B vssd1 vssd1 vccd1 vccd1 _13670_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_251_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10882_ _15150_/C1 _15267_/A _10851_/Y vssd1 vssd1 vccd1 vccd1 _11322_/B sky130_fd_sc_hd__o21ba_4
XFILLER_216_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _12916_/B2 _12618_/X _12916_/A2 _19524_/Q vssd1 vssd1 vccd1 vccd1 _12911_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ _20793_/Q _15016_/A _15021_/X _15339_/X vssd1 vssd1 vccd1 vccd1 _15340_/X
+ sky130_fd_sc_hd__a211o_4
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _12552_/A _12552_/B _12552_/C _12552_/D vssd1 vssd1 vccd1 vccd1 _12554_/B
+ sky130_fd_sc_hd__or4_1
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11503_ _11514_/A1 _12120_/A1 _19350_/Q _12046_/B1 vssd1 vssd1 vccd1 vccd1 _11503_/X
+ sky130_fd_sc_hd__a31o_1
X_15271_ _21017_/Q _20985_/Q _15508_/S vssd1 vssd1 vccd1 vccd1 _15271_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12483_ split8/X _12847_/A2 _15526_/A vssd1 vssd1 vccd1 vccd1 _12483_/Y sky130_fd_sc_hd__a21oi_4
X_17010_ _16950_/Y _17009_/X _16875_/B2 vssd1 vssd1 vccd1 vccd1 _17010_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_200_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14222_ _14218_/B _14221_/Y _14233_/S vssd1 vssd1 vccd1 vccd1 _14222_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11434_ _12125_/A1 _11420_/X _11421_/X vssd1 vssd1 vccd1 vccd1 _11434_/X sky130_fd_sc_hd__o21a_1
XFILLER_184_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14153_ _18763_/A1 _14152_/X _13507_/X vssd1 vssd1 vccd1 vccd1 _14154_/C sky130_fd_sc_hd__a21o_1
X_11365_ _11347_/X _11364_/X _12401_/A1 vssd1 vssd1 vccd1 vccd1 _11365_/X sky130_fd_sc_hd__a21o_2
XFILLER_138_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20077_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_256_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13104_ _19245_/Q _13104_/B vssd1 vssd1 vccd1 vccd1 _13104_/X sky130_fd_sc_hd__or2_1
X_10316_ _20411_/Q _20347_/Q _10316_/S vssd1 vssd1 vccd1 vccd1 _10316_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14084_ _19201_/Q _14104_/A2 _14083_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1 _19201_/D
+ sky130_fd_sc_hd__o211a_1
X_18961_ _19113_/Q _18974_/A2 _12591_/X _15981_/A vssd1 vssd1 vccd1 vccd1 _18961_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11296_ _19662_/Q _20150_/Q _11303_/S vssd1 vssd1 vccd1 vccd1 _11296_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17912_ _20683_/Q _12040_/X _17912_/S vssd1 vssd1 vccd1 vccd1 _20683_/D sky130_fd_sc_hd__mux2_1
X_13035_ _20960_/Q _20894_/Q vssd1 vssd1 vccd1 vccd1 _13035_/Y sky130_fd_sc_hd__nor2_2
X_10247_ _12429_/A1 _10245_/X _10246_/X vssd1 vssd1 vccd1 vccd1 _10247_/X sky130_fd_sc_hd__o21a_1
X_18892_ _19103_/Q _18954_/A2 _18967_/B1 _13428_/C vssd1 vssd1 vccd1 vccd1 _18893_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1120 _17939_/A1 vssd1 vssd1 vccd1 vccd1 _17696_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_239_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1131 _11454_/X vssd1 vssd1 vccd1 vccd1 _17937_/A1 sky130_fd_sc_hd__buf_4
X_17843_ _20618_/Q _17881_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20618_/D sky130_fd_sc_hd__mux2_1
Xfanout1142 _09936_/A2 vssd1 vssd1 vccd1 vccd1 _17835_/A1 sky130_fd_sc_hd__buf_4
XFILLER_79_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10178_ _10262_/A _20378_/Q _20442_/Q _11303_/S vssd1 vssd1 vccd1 vccd1 _10178_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1153 _13670_/A1 vssd1 vssd1 vccd1 vccd1 _12157_/A1 sky130_fd_sc_hd__buf_12
XFILLER_94_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1164 _15673_/B1 vssd1 vssd1 vccd1 vccd1 _16051_/B1 sky130_fd_sc_hd__buf_4
Xfanout1175 _13730_/B vssd1 vssd1 vccd1 vccd1 _13742_/B sky130_fd_sc_hd__buf_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1186 _12485_/Y vssd1 vssd1 vccd1 vccd1 _15977_/A1 sky130_fd_sc_hd__buf_6
Xfanout1197 _17302_/C vssd1 vssd1 vccd1 vccd1 _17305_/C sky130_fd_sc_hd__buf_4
X_17774_ _20553_/Q _17914_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20553_/D sky130_fd_sc_hd__mux2_1
X_14986_ _17272_/A _15308_/B _14986_/C vssd1 vssd1 vccd1 vccd1 _14986_/X sky130_fd_sc_hd__and3_1
XFILLER_208_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19513_ _20913_/CLK _19513_/D vssd1 vssd1 vccd1 vccd1 _19513_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_263_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16725_ _16723_/X _16724_/X _12930_/B vssd1 vssd1 vccd1 vccd1 _16725_/X sky130_fd_sc_hd__a21bo_1
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13937_ _19141_/Q _13941_/B _13946_/B1 _13242_/C vssd1 vssd1 vccd1 vccd1 _19141_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_263_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19444_ _20703_/CLK _19444_/D vssd1 vssd1 vccd1 vccd1 _19444_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13868_ _19087_/Q _13902_/B _13867_/Y _15288_/C1 vssd1 vssd1 vccd1 vccd1 _19087_/D
+ sky130_fd_sc_hd__o211a_1
X_16656_ _19913_/Q _17693_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19913_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12819_ _19517_/Q _12916_/A2 _12818_/X _12916_/B2 vssd1 vssd1 vccd1 vccd1 _12820_/B
+ sky130_fd_sc_hd__o22a_2
X_15607_ _15644_/A1 _16869_/B _15593_/Y vssd1 vssd1 vccd1 vccd1 _15607_/Y sky130_fd_sc_hd__o21ai_1
X_19375_ _20666_/CLK _19375_/D vssd1 vssd1 vccd1 vccd1 _19375_/Q sky130_fd_sc_hd__dfxtp_1
X_16587_ _16591_/A _16587_/B vssd1 vssd1 vccd1 vccd1 _19859_/D sky130_fd_sc_hd__or2_1
X_13799_ _13816_/A1 _13668_/Y split9/A input245/X vssd1 vssd1 vccd1 vccd1 _13799_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18326_ _20818_/Q _18341_/B _18325_/Y _18692_/A vssd1 vssd1 vccd1 vccd1 _20818_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15538_ _20799_/Q _15016_/A _15536_/X _15537_/X vssd1 vssd1 vccd1 vccd1 _15538_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_148_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18257_ _18728_/A _18257_/B vssd1 vssd1 vccd1 vccd1 _20805_/D sky130_fd_sc_hd__and2_1
X_15469_ _15610_/A1 _15212_/X _15610_/B1 vssd1 vssd1 vccd1 vccd1 _15736_/B sky130_fd_sc_hd__o21ai_4
XFILLER_191_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17208_ _20172_/Q _17942_/A1 _17212_/S vssd1 vssd1 vccd1 vccd1 _20172_/D sky130_fd_sc_hd__mux2_1
XFILLER_200_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ _19533_/Q _18198_/B vssd1 vssd1 vccd1 vccd1 _18188_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_156_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _20107_/Q _17801_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20107_/D sky130_fd_sc_hd__mux2_1
XFILLER_265_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20150_ _20557_/CLK _20150_/D vssd1 vssd1 vccd1 vccd1 _20150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09961_ _09959_/X _09960_/X _11902_/S vssd1 vssd1 vccd1 vccd1 _09961_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20081_ _20081_/CLK _20081_/D vssd1 vssd1 vccd1 vccd1 _20081_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _12150_/S _09891_/X _09890_/X _12140_/C1 vssd1 vssd1 vccd1 vccd1 _09892_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20983_ _21015_/CLK _20983_/D vssd1 vssd1 vccd1 vccd1 _20983_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_509 input215/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_74_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20694_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_214_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20417_ _20425_/CLK _20417_/D vssd1 vssd1 vccd1 vccd1 _20417_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_135_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11150_ _11234_/A _11150_/B vssd1 vssd1 vccd1 vccd1 _11150_/X sky130_fd_sc_hd__and2_1
XFILLER_175_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20348_ _20465_/CLK _20348_/D vssd1 vssd1 vccd1 vccd1 _20348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10101_ _10409_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10101_/X sky130_fd_sc_hd__or2_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11081_ _20495_/Q _12213_/B vssd1 vssd1 vccd1 vccd1 _11081_/X sky130_fd_sc_hd__or2_1
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20279_ _20990_/CLK _20279_/D vssd1 vssd1 vccd1 vccd1 _20279_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput201 localMemory_wb_adr_i[1] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_hd__clkbuf_2
XFILLER_103_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10032_ _10465_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _10032_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput212 localMemory_wb_adr_i[8] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput223 localMemory_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_hd__buf_12
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput234 localMemory_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_hd__buf_12
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 localMemory_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_hd__buf_12
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput256 manufacturerID[2] vssd1 vssd1 vccd1 vccd1 _17245_/A sky130_fd_sc_hd__buf_2
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput267 partID[12] vssd1 vssd1 vccd1 vccd1 input267/X sky130_fd_sc_hd__clkbuf_2
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _14839_/X _14832_/X _15215_/S vssd1 vssd1 vccd1 vccd1 _14840_/X sky130_fd_sc_hd__mux2_1
Xinput278 partID[8] vssd1 vssd1 vccd1 vccd1 _17296_/A sky130_fd_sc_hd__clkbuf_2
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14771_ _19510_/Q _14773_/B vssd1 vssd1 vccd1 vccd1 _14771_/X sky130_fd_sc_hd__or2_1
X_11983_ _11983_/A1 _20520_/Q _11980_/S _11965_/X vssd1 vssd1 vccd1 vccd1 _11983_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13722_ _13722_/A _13742_/B vssd1 vssd1 vccd1 vccd1 _13762_/B sky130_fd_sc_hd__or2_2
X_16510_ _19817_/Q _17905_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19817_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ _10931_/X _10932_/Y _11313_/B vssd1 vssd1 vccd1 vccd1 _15118_/S sky130_fd_sc_hd__a21o_4
XFILLER_232_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17490_ _20280_/Q _17494_/B vssd1 vssd1 vccd1 vccd1 _17490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_216_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13653_ _13653_/A _13653_/B vssd1 vssd1 vccd1 vccd1 _13689_/C sky130_fd_sc_hd__nand2_2
X_16441_ _19760_/Q _16442_/C _19761_/Q vssd1 vssd1 vccd1 vccd1 _16443_/B sky130_fd_sc_hd__a21oi_1
X_10865_ _10863_/X _10864_/X _12414_/S vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12604_ _19508_/Q _19507_/Q _12740_/B vssd1 vssd1 vccd1 vccd1 _12718_/A sky130_fd_sc_hd__and3_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _19735_/Q _16372_/B vssd1 vssd1 vccd1 vccd1 _16378_/C sky130_fd_sc_hd__and2_2
X_19160_ _19560_/CLK _19160_/D vssd1 vssd1 vccd1 vccd1 _19160_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _13624_/B2 _15369_/A _13583_/Y _13478_/B vssd1 vssd1 vccd1 vccd1 _13584_/X
+ sky130_fd_sc_hd__a22o_4
X_10796_ _12277_/A1 _17926_/A1 _10795_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _15304_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_158_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15323_ _15323_/A _15323_/B _15388_/S vssd1 vssd1 vccd1 vccd1 _15323_/X sky130_fd_sc_hd__or3_2
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _20779_/Q _18111_/B vssd1 vssd1 vccd1 vccd1 _18117_/C sky130_fd_sc_hd__and2_2
XFILLER_200_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ _20873_/Q _12549_/B _12535_/C vssd1 vssd1 vccd1 vccd1 _12553_/A sky130_fd_sc_hd__and3_1
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19091_ _19620_/CLK _19091_/D vssd1 vssd1 vccd1 vccd1 _19091_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_173_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18042_ _20753_/Q _18045_/C _18704_/A vssd1 vssd1 vccd1 vccd1 _18042_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_172_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15254_ _15056_/X _15063_/X _15254_/S vssd1 vssd1 vccd1 vccd1 _15254_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12466_ _14895_/A _15026_/A vssd1 vssd1 vccd1 vccd1 _12466_/Y sky130_fd_sc_hd__nand2_8
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14205_ _19223_/Q _14205_/A2 _14204_/X _18710_/A vssd1 vssd1 vccd1 vccd1 _19223_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ _11415_/A _10367_/Y _11413_/Y _11415_/X _11416_/Y vssd1 vssd1 vccd1 vccd1
+ _11791_/B sky130_fd_sc_hd__o311a_2
X_15185_ _15185_/A _15185_/B vssd1 vssd1 vccd1 vccd1 _15185_/X sky130_fd_sc_hd__or2_1
X_12397_ _19297_/Q _20084_/Q _12397_/S vssd1 vssd1 vccd1 vccd1 _12397_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14136_ _20268_/Q _14117_/A _14216_/B1 input237/X vssd1 vssd1 vccd1 vccd1 _14139_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ _20030_/Q _12300_/S vssd1 vssd1 vccd1 vccd1 _11348_/X sky130_fd_sc_hd__or2_1
XFILLER_113_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19993_ _20621_/CLK _19993_/D vssd1 vssd1 vccd1 vccd1 _19993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14067_ _14107_/A _14069_/B _14067_/C vssd1 vssd1 vccd1 vccd1 _14067_/X sky130_fd_sc_hd__or3_1
X_18944_ _21006_/Q _18964_/B vssd1 vssd1 vccd1 vccd1 _18944_/Y sky130_fd_sc_hd__nand2_1
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11279_ _19157_/Q _12569_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11279_/X sky130_fd_sc_hd__o21ba_1
XFILLER_267_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13018_ _20970_/Q _20904_/Q vssd1 vssd1 vccd1 vccd1 _13194_/B sky130_fd_sc_hd__nand2_2
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18875_ _20996_/Q _18937_/B vssd1 vssd1 vccd1 vccd1 _18875_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17826_ _20601_/Q _17898_/A1 _17840_/S vssd1 vssd1 vccd1 vccd1 _20601_/D sky130_fd_sc_hd__mux2_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17757_ _20536_/Q split4/A _17772_/S vssd1 vssd1 vccd1 vccd1 _20536_/D sky130_fd_sc_hd__mux2_1
XFILLER_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14969_ _15314_/D _15019_/A _15021_/B vssd1 vssd1 vccd1 vccd1 _14971_/B sky130_fd_sc_hd__and3b_1
XFILLER_208_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16708_ _16878_/A _16708_/B vssd1 vssd1 vccd1 vccd1 _16708_/Y sky130_fd_sc_hd__nand2_1
X_17688_ _20472_/Q _17931_/A1 _17703_/S vssd1 vssd1 vccd1 vccd1 _20472_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19427_ _20586_/CLK _19427_/D vssd1 vssd1 vccd1 vccd1 _19427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16639_ _17851_/A _17676_/B _16639_/C vssd1 vssd1 vccd1 vccd1 _16639_/X sky130_fd_sc_hd__and3_4
XFILLER_251_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19358_ _20713_/CLK _19358_/D vssd1 vssd1 vccd1 vccd1 _19358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18309_ _18308_/B _14423_/B _18308_/Y vssd1 vssd1 vccd1 vccd1 _18556_/B sky130_fd_sc_hd__o21ai_4
XFILLER_148_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19289_ _20479_/CLK _19289_/D vssd1 vssd1 vccd1 vccd1 _19289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_192_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19607_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_128_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20202_ _20760_/CLK _20202_/D vssd1 vssd1 vccd1 vccd1 _20202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_121_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20751_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _11242_/A1 _14011_/A2 _09943_/X _11242_/B1 _19851_/Q vssd1 vssd1 vccd1 vccd1
+ _09944_/X sky130_fd_sc_hd__o32a_1
Xfanout902 _15020_/Y vssd1 vssd1 vccd1 vccd1 _15388_/S sky130_fd_sc_hd__buf_6
X_20133_ _20557_/CLK _20133_/D vssd1 vssd1 vccd1 vccd1 _20133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout913 _14995_/Y vssd1 vssd1 vccd1 vccd1 _15322_/B sky130_fd_sc_hd__buf_6
XFILLER_131_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout924 _14935_/Y vssd1 vssd1 vccd1 vccd1 _15989_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout935 _11223_/A vssd1 vssd1 vccd1 vccd1 _15165_/S sky130_fd_sc_hd__buf_6
XFILLER_225_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout946 _11017_/X vssd1 vssd1 vccd1 vccd1 _15545_/A sky130_fd_sc_hd__buf_6
X_20064_ _20671_/CLK _20064_/D vssd1 vssd1 vccd1 vccd1 _20064_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout957 _17788_/A1 vssd1 vssd1 vccd1 vccd1 _17928_/A1 sky130_fd_sc_hd__clkbuf_4
X_09875_ _19419_/Q _11818_/B2 _09874_/X _11892_/C1 vssd1 vssd1 vccd1 vccd1 _09875_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout968 _10474_/X vssd1 vssd1 vccd1 vccd1 _17060_/A1 sky130_fd_sc_hd__buf_2
XFILLER_219_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout979 _17692_/A1 vssd1 vssd1 vccd1 vccd1 _17935_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 input233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_317 _13478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_328 _20258_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20966_ _21040_/CLK _20966_/D vssd1 vssd1 vccd1 vccd1 _20966_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_339 _19519_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20897_ _21027_/CLK _20897_/D vssd1 vssd1 vccd1 vccd1 _20897_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_201_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10650_ _19405_/Q _20564_/Q _12368_/S vssd1 vssd1 vccd1 vccd1 _10650_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10581_ _10581_/A1 _20666_/Q _12064_/S _19375_/Q _10585_/S vssd1 vssd1 vccd1 vccd1
+ _10581_/X sky130_fd_sc_hd__o221a_1
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12320_ _19829_/Q _19333_/Q _12323_/S vssd1 vssd1 vccd1 vccd1 _12320_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_209_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20717_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_214_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _19652_/Q _19958_/Q _19296_/Q _20083_/Q _12339_/S0 _12337_/C vssd1 vssd1
+ vccd1 vccd1 _12251_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11202_ _20119_/Q _20087_/Q _11203_/S vssd1 vssd1 vccd1 vccd1 _11202_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _19826_/Q _19330_/Q _12182_/S vssd1 vssd1 vccd1 vccd1 _12182_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11133_ _12277_/A1 _17782_/A1 _11132_/X _09750_/Y vssd1 vssd1 vccd1 vccd1 _12668_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16990_ _17008_/A1 _16989_/X _17008_/B1 vssd1 vssd1 vccd1 vccd1 _16990_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_150_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11064_ _20463_/Q _20303_/Q _12397_/S vssd1 vssd1 vccd1 vccd1 _11064_/X sky130_fd_sc_hd__mux2_1
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15941_ _20813_/Q _15941_/A2 _15934_/X _15941_/B2 _15940_/X vssd1 vssd1 vccd1 vccd1
+ _15941_/X sky130_fd_sc_hd__a221o_4
XFILLER_95_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10015_ _11742_/A _11742_/B vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__nand2b_2
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18660_ _18538_/X _18684_/A2 _18658_/Y _18659_/Y vssd1 vssd1 vccd1 vccd1 _18661_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15872_ _19727_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15872_/X sky130_fd_sc_hd__or2_1
XFILLER_264_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17611_ _20367_/Q _17922_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20367_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ _14821_/X _14822_/X _15039_/A vssd1 vssd1 vccd1 vccd1 _14823_/X sky130_fd_sc_hd__mux2_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _18783_/A _18591_/B vssd1 vssd1 vccd1 vccd1 _20920_/D sky130_fd_sc_hd__nor2_1
XFILLER_224_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17542_ _20302_/Q _17678_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20302_/D sky130_fd_sc_hd__mux2_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14754_ _19124_/Q _14764_/A2 _14753_/X _18710_/A vssd1 vssd1 vccd1 vccd1 _19501_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11966_ _19956_/Q _12044_/B vssd1 vssd1 vccd1 vccd1 _11966_/X sky130_fd_sc_hd__or2_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10917_ _09618_/A _11008_/A1 _20122_/Q _11345_/S vssd1 vssd1 vccd1 vccd1 _10917_/X
+ sky130_fd_sc_hd__a31o_1
X_13705_ _13703_/Y _13704_/X _13714_/S vssd1 vssd1 vccd1 vccd1 _13706_/B sky130_fd_sc_hd__mux2_8
X_17473_ _17487_/A1 _17472_/Y _18704_/A vssd1 vssd1 vccd1 vccd1 _20271_/D sky130_fd_sc_hd__a21oi_1
XFILLER_189_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14685_ _19444_/Q _17657_/A1 _14685_/S vssd1 vssd1 vccd1 vccd1 _19444_/D sky130_fd_sc_hd__mux2_1
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11897_ _19954_/Q _11897_/B vssd1 vssd1 vccd1 vccd1 _11897_/X sky130_fd_sc_hd__or2_1
XFILLER_260_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19212_ _20759_/CLK _19212_/D vssd1 vssd1 vccd1 vccd1 _19212_/Q sky130_fd_sc_hd__dfxtp_1
X_13636_ _13636_/A _13658_/A vssd1 vssd1 vccd1 vccd1 _13777_/A sky130_fd_sc_hd__nand2_8
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16424_ _19754_/Q _16426_/C _16423_/Y vssd1 vssd1 vccd1 vccd1 _19754_/D sky130_fd_sc_hd__o21a_1
X_10848_ _12245_/A1 _17925_/A1 _10847_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _13653_/B
+ sky130_fd_sc_hd__o211a_4
X_19143_ _19520_/CLK _19143_/D vssd1 vssd1 vccd1 vccd1 _19143_/Q sky130_fd_sc_hd__dfxtp_1
X_13567_ _13567_/A _13567_/B vssd1 vssd1 vccd1 vccd1 _13568_/A sky130_fd_sc_hd__xor2_4
XFILLER_13_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16355_ _18835_/A _16355_/B _16356_/B vssd1 vssd1 vccd1 vccd1 _19728_/D sky130_fd_sc_hd__nor3_1
X_10779_ _20467_/Q _20307_/Q _12268_/S vssd1 vssd1 vccd1 vccd1 _10779_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15306_ _20728_/Q _15445_/A2 _15445_/B1 _20760_/Q vssd1 vssd1 vccd1 vccd1 _15306_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12518_ _13192_/A _18765_/B _12518_/C _11367_/A vssd1 vssd1 vccd1 vccd1 _12520_/C
+ sky130_fd_sc_hd__or4b_1
X_16286_ _19702_/Q _19703_/Q _18054_/A vssd1 vssd1 vccd1 vccd1 _16286_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_146_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19074_ _20419_/Q vssd1 vssd1 vccd1 vccd1 _20419_/D sky130_fd_sc_hd__clkbuf_2
X_13498_ _19218_/Q _13498_/B vssd1 vssd1 vccd1 vccd1 _13499_/B sky130_fd_sc_hd__nor2_1
XFILLER_145_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18025_ _18112_/A _18030_/C vssd1 vssd1 vccd1 vccd1 _18025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_246_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15237_ _20854_/Q _15236_/X _15601_/S vssd1 vssd1 vccd1 vccd1 _15237_/X sky130_fd_sc_hd__mux2_1
X_12449_ _12449_/A _12450_/A _12449_/C vssd1 vssd1 vccd1 vccd1 _12449_/X sky130_fd_sc_hd__and3_1
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15168_ _15168_/A vssd1 vssd1 vccd1 vccd1 _15168_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14119_ _14119_/A _14119_/B vssd1 vssd1 vccd1 vccd1 _16710_/B sky130_fd_sc_hd__or2_2
X_19976_ _20014_/CLK _19976_/D vssd1 vssd1 vccd1 vccd1 _19976_/Q sky130_fd_sc_hd__dfxtp_1
X_15099_ _15365_/A _15076_/Y _15077_/X _15074_/X vssd1 vssd1 vccd1 vccd1 _15099_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_262_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18927_ _18975_/A _18927_/B vssd1 vssd1 vccd1 vccd1 _18927_/Y sky130_fd_sc_hd__nand2_2
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09660_ _19566_/Q _11243_/S vssd1 vssd1 vccd1 vccd1 _09660_/X sky130_fd_sc_hd__or2_1
XFILLER_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18858_ _18968_/A _18858_/B vssd1 vssd1 vccd1 vccd1 _18858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_267_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17809_ _20586_/Q _17949_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20586_/D sky130_fd_sc_hd__mux2_1
XFILLER_209_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09591_ _09592_/A _09592_/C vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__nand2_1
X_18789_ _18787_/X _18788_/X _18476_/A vssd1 vssd1 vccd1 vccd1 _20983_/D sky130_fd_sc_hd__o21a_1
XFILLER_283_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20820_ _21016_/CLK _20820_/D vssd1 vssd1 vccd1 vccd1 _20820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20751_ _20751_/CLK _20751_/D vssd1 vssd1 vccd1 vccd1 _20751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20682_ _20682_/CLK _20682_/D vssd1 vssd1 vccd1 vccd1 _20682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1708 _11537_/A1 vssd1 vssd1 vccd1 vccd1 _09730_/A sky130_fd_sc_hd__buf_6
Xfanout710 _13822_/A1 vssd1 vssd1 vccd1 vccd1 _13810_/A1 sky130_fd_sc_hd__buf_2
Xfanout1719 _11983_/A1 vssd1 vssd1 vccd1 vccd1 _12120_/A1 sky130_fd_sc_hd__buf_6
Xfanout721 _13775_/A vssd1 vssd1 vccd1 vccd1 _13780_/A sky130_fd_sc_hd__buf_2
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20116_ _20180_/CLK _20116_/D vssd1 vssd1 vccd1 vccd1 _20116_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout732 _19015_/B vssd1 vssd1 vccd1 vccd1 _19049_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_259_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _19683_/Q _20171_/Q _09928_/S vssd1 vssd1 vccd1 vccd1 _09927_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout743 _18818_/A2 vssd1 vssd1 vccd1 vccd1 _18970_/A2 sky130_fd_sc_hd__buf_6
Xfanout754 _18964_/B vssd1 vssd1 vccd1 vccd1 _18971_/B sky130_fd_sc_hd__buf_4
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout765 _13183_/Y vssd1 vssd1 vccd1 vccd1 _15954_/A sky130_fd_sc_hd__buf_8
XFILLER_246_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout776 _12592_/X vssd1 vssd1 vccd1 vccd1 _18902_/A sky130_fd_sc_hd__buf_6
X_09858_ _19516_/Q _15795_/A _15895_/S vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__mux2_8
X_20047_ _20047_/CLK _20047_/D vssd1 vssd1 vccd1 vccd1 _20047_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout787 _12525_/Y vssd1 vssd1 vccd1 vccd1 _13575_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_246_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout798 _12487_/Y vssd1 vssd1 vccd1 vccd1 _12982_/B sky130_fd_sc_hd__buf_4
XFILLER_207_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _12366_/A1 _10285_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__a21o_2
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _12486_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _20142_/Q _20110_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _11820_/X sky130_fd_sc_hd__mux2_1
XANTENNA_114 _13603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_125 _13656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_136 _13683_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _13738_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _13420_/A _11794_/C _11736_/Y vssd1 vssd1 vccd1 vccd1 _11752_/B sky130_fd_sc_hd__o21ba_2
XFILLER_82_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_158 _13780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_169 _19108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20949_ _20949_/CLK _20949_/D vssd1 vssd1 vccd1 vccd1 _20949_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _10692_/A _19469_/Q _19437_/Q _12268_/S _12419_/C1 vssd1 vssd1 vccd1 vccd1
+ _10702_/X sky130_fd_sc_hd__a221o_1
XFILLER_241_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14470_ _18700_/A _14470_/B vssd1 vssd1 vccd1 vccd1 _19259_/D sky130_fd_sc_hd__and2_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11682_ _19285_/Q _20072_/Q _11682_/S vssd1 vssd1 vccd1 vccd1 _11682_/X sky130_fd_sc_hd__mux2_1
XFILLER_241_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13421_ _13421_/A _13421_/B vssd1 vssd1 vccd1 vccd1 _13427_/C sky130_fd_sc_hd__xnor2_4
X_10633_ _12105_/A _10632_/X _10617_/X vssd1 vssd1 vccd1 vccd1 _10633_/X sky130_fd_sc_hd__o21a_2
XFILLER_167_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16140_ _16754_/B _16194_/S vssd1 vssd1 vccd1 vccd1 _16140_/Y sky130_fd_sc_hd__nand2_1
XFILLER_220_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _13352_/A _13352_/B _13352_/C vssd1 vssd1 vccd1 vccd1 _13352_/X sky130_fd_sc_hd__and3_1
X_10564_ _12051_/A1 _20374_/Q _20438_/Q _11994_/S _11995_/S vssd1 vssd1 vccd1 vccd1
+ _10564_/X sky130_fd_sc_hd__a221o_1
X_12303_ _19896_/Q _12389_/S vssd1 vssd1 vccd1 vccd1 _12303_/X sky130_fd_sc_hd__or2_1
XFILLER_6_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16071_ _16071_/A _16081_/B vssd1 vssd1 vccd1 vccd1 _16071_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13283_ _12748_/X _13281_/Y _13282_/Y vssd1 vssd1 vccd1 vccd1 _13283_/X sky130_fd_sc_hd__o21a_1
X_10495_ _19376_/Q _09689_/D _10493_/X _11274_/B2 _10494_/X vssd1 vssd1 vccd1 vccd1
+ _10495_/X sky130_fd_sc_hd__o221a_1
XFILLER_142_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15022_ _15022_/A _15022_/B _15022_/C _15022_/D vssd1 vssd1 vccd1 vccd1 _15334_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_182_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12234_ _19395_/Q _20686_/Q _12313_/S vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19830_ _21040_/CLK _19830_/D vssd1 vssd1 vccd1 vccd1 _19830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12165_ _20425_/Q _20361_/Q _12165_/S vssd1 vssd1 vccd1 vccd1 _12166_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ _20463_/Q _20303_/Q _11116_/S vssd1 vssd1 vccd1 vccd1 _11116_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19761_ _19970_/CLK _19761_/D vssd1 vssd1 vccd1 vccd1 _19761_/Q sky130_fd_sc_hd__dfxtp_1
X_12096_ _12828_/A _12091_/X _12095_/Y _12850_/A1 vssd1 vssd1 vccd1 vccd1 _12105_/B
+ sky130_fd_sc_hd__o211a_1
X_16973_ _16981_/A1 _15943_/X _16945_/X _16972_/X vssd1 vssd1 vccd1 vccd1 _16973_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_284_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18712_ _18985_/A _18712_/B vssd1 vssd1 vccd1 vccd1 _20956_/D sky130_fd_sc_hd__and2_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ _12275_/A _11047_/B vssd1 vssd1 vccd1 vccd1 _11047_/Y sky130_fd_sc_hd__nor2_1
X_15924_ _19553_/Q _15814_/A _15923_/X _16185_/A vssd1 vssd1 vccd1 vccd1 _19553_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19692_ _20586_/CLK _19692_/D vssd1 vssd1 vccd1 vccd1 _19692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_249_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput9 core_wb_ack_i vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18643_ _20934_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18643_/Y sky130_fd_sc_hd__nand2_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _20906_/Q _16043_/A2 _16043_/B1 _15854_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _15855_/X sky130_fd_sc_hd__a221o_1
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _15365_/A _15095_/B vssd1 vssd1 vccd1 vccd1 _14897_/B sky130_fd_sc_hd__nand2_2
X_18574_ _19496_/Q _18760_/B vssd1 vssd1 vccd1 vccd1 _18574_/Y sky130_fd_sc_hd__nand2_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15786_ _19171_/Q _15978_/A2 _15762_/A _16063_/B2 vssd1 vssd1 vccd1 vccd1 _15787_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _19243_/Q _13114_/B vssd1 vssd1 vccd1 vccd1 _12998_/Y sky130_fd_sc_hd__nand2_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ _17525_/A1 _17524_/Y _17430_/A vssd1 vssd1 vccd1 vccd1 _20297_/D sky130_fd_sc_hd__a21oi_1
XFILLER_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14737_ _19149_/Q _16133_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _14737_/X sky130_fd_sc_hd__and3b_4
X_11949_ _11945_/X _11948_/X _11949_/S vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17456_ _17443_/C _17456_/B vssd1 vssd1 vccd1 vccd1 _17456_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_60_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14668_ _19093_/Q _14668_/B _17538_/C vssd1 vssd1 vccd1 vccd1 _16604_/B sky130_fd_sc_hd__or3_2
XFILLER_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16407_ _19748_/Q _16410_/C _18094_/A vssd1 vssd1 vccd1 vccd1 _16407_/Y sky130_fd_sc_hd__a21oi_1
X_13619_ _13626_/A1 _13359_/Y _13427_/C _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13619_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_220_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17387_ _20242_/Q _17401_/A2 _17386_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _20242_/D
+ sky130_fd_sc_hd__o211a_1
X_14599_ _19365_/Q _17951_/A1 _14599_/S vssd1 vssd1 vccd1 vccd1 _19365_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19126_ _19505_/CLK _19126_/D vssd1 vssd1 vccd1 vccd1 _19126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16338_ _19721_/Q _19722_/Q _16338_/C vssd1 vssd1 vccd1 vccd1 _16340_/B sky130_fd_sc_hd__and3_1
XFILLER_9_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19057_ _20402_/Q vssd1 vssd1 vccd1 vccd1 _20402_/D sky130_fd_sc_hd__clkbuf_2
X_16269_ _19685_/Q _17943_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19685_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput302 _13789_/X vssd1 vssd1 vccd1 vccd1 addr1[8] sky130_fd_sc_hd__buf_4
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18008_ _20741_/Q _18011_/C _18096_/A vssd1 vssd1 vccd1 vccd1 _18008_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_161_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput313 _13620_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[17] sky130_fd_sc_hd__buf_4
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput324 _13630_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[27] sky130_fd_sc_hd__buf_4
Xoutput335 _13679_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[10] sky130_fd_sc_hd__buf_4
XFILLER_99_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput346 _13725_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[20] sky130_fd_sc_hd__buf_4
XFILLER_142_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput357 _13775_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[30] sky130_fd_sc_hd__buf_4
XFILLER_259_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput368 _13638_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[2] sky130_fd_sc_hd__buf_4
XFILLER_273_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput379 _13803_/X vssd1 vssd1 vccd1 vccd1 din0[12] sky130_fd_sc_hd__buf_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19959_ _20463_/CLK _19959_/D vssd1 vssd1 vccd1 vccd1 _19959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ _11917_/S _09711_/X _09710_/X _12151_/A1 vssd1 vssd1 vccd1 vccd1 _09712_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_101_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09643_ _09643_/A _09686_/D vssd1 vssd1 vccd1 vccd1 _09643_/Y sky130_fd_sc_hd__nor2_1
XFILLER_110_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _14112_/A _19096_/Q vssd1 vssd1 vccd1 vccd1 _09592_/A sky130_fd_sc_hd__nand2b_4
XFILLER_55_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20803_ _20990_/CLK _20803_/D vssd1 vssd1 vccd1 vccd1 _20803_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20734_ _20796_/CLK _20734_/D vssd1 vssd1 vccd1 vccd1 _20734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20665_ _20665_/CLK _20665_/D vssd1 vssd1 vccd1 vccd1 _20665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20596_ _20655_/CLK _20596_/D vssd1 vssd1 vccd1 vccd1 _20596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10280_ _19541_/Q _09596_/A _09613_/B _19605_/Q _11246_/A1 vssd1 vssd1 vccd1 vccd1
+ _10280_/X sky130_fd_sc_hd__a221o_1
XFILLER_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1505 _11818_/B2 vssd1 vssd1 vccd1 vccd1 _11891_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_132_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1516 fanout1522/X vssd1 vssd1 vccd1 vccd1 _12121_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_278_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1527 fanout1534/X vssd1 vssd1 vccd1 vccd1 _11665_/S sky130_fd_sc_hd__buf_4
Xfanout1538 _10316_/S vssd1 vssd1 vccd1 vccd1 _10303_/S sky130_fd_sc_hd__buf_6
Xfanout540 _17178_/S vssd1 vssd1 vccd1 vccd1 _17180_/S sky130_fd_sc_hd__buf_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout551 _17083_/X vssd1 vssd1 vccd1 vccd1 _17114_/S sky130_fd_sc_hd__buf_6
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1549 fanout1556/X vssd1 vssd1 vccd1 vccd1 _11342_/S sky130_fd_sc_hd__buf_6
Xfanout562 _16639_/X vssd1 vssd1 vccd1 vccd1 _16671_/S sky130_fd_sc_hd__buf_12
X_13970_ _19189_/Q _14059_/C _14042_/S vssd1 vssd1 vccd1 vccd1 _13970_/X sky130_fd_sc_hd__mux2_2
Xfanout573 _16456_/X vssd1 vssd1 vccd1 vccd1 _16483_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_281_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout584 _16126_/A2 vssd1 vssd1 vccd1 vccd1 _16132_/A2 sky130_fd_sc_hd__buf_4
XFILLER_219_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout595 _14699_/S vssd1 vssd1 vccd1 vccd1 _14698_/S sky130_fd_sc_hd__buf_12
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _20299_/Q _17526_/C _20300_/Q vssd1 vssd1 vccd1 vccd1 _12921_/X sky130_fd_sc_hd__and3b_4
XFILLER_47_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15640_ _20802_/Q _16047_/A2 _15632_/X _16000_/A1 _15639_/X vssd1 vssd1 vccd1 vccd1
+ _15640_/X sky130_fd_sc_hd__a221o_1
XFILLER_74_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12852_/A _12852_/B _12852_/C vssd1 vssd1 vccd1 vccd1 _12853_/B sky130_fd_sc_hd__nand3_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11803_ _13413_/A _11802_/Y _11799_/Y vssd1 vssd1 vccd1 vccd1 _11804_/B sky130_fd_sc_hd__o21a_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _20800_/Q _15016_/A _15569_/X _15570_/X vssd1 vssd1 vccd1 vccd1 _15571_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _14803_/A1 _12582_/C _12784_/B _12782_/X vssd1 vssd1 vccd1 vccd1 _12783_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _20209_/Q _17328_/A2 _17309_/X _18416_/A vssd1 vssd1 vccd1 vccd1 _20209_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _11495_/A _11734_/B vssd1 vssd1 vccd1 vccd1 _11734_/Y sky130_fd_sc_hd__nand2b_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _14522_/A _14522_/B vssd1 vssd1 vccd1 vccd1 _19299_/D sky130_fd_sc_hd__nor2_1
X_18290_ _18544_/B vssd1 vssd1 vccd1 vccd1 _18290_/Y sky130_fd_sc_hd__clkinv_2
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _20186_/Q _17268_/A2 _17239_/X _17240_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1
+ _20186_/D sky130_fd_sc_hd__o221a_1
X_14453_ _20222_/Q _19251_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14454_/B sky130_fd_sc_hd__mux2_1
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11665_ _20136_/Q _20104_/Q _11665_/S vssd1 vssd1 vccd1 vccd1 _11665_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10616_ _10610_/X _10612_/X _10615_/X _10409_/A vssd1 vssd1 vccd1 vccd1 _10616_/X
+ sky130_fd_sc_hd__a211o_1
X_13404_ _20929_/Q _13350_/B _13323_/C _13403_/X _18628_/B vssd1 vssd1 vccd1 vccd1
+ _13404_/X sky130_fd_sc_hd__a221o_1
X_17172_ _20138_/Q _17800_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20138_/D sky130_fd_sc_hd__mux2_1
X_14384_ _14382_/Y _14384_/B vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__nand2b_1
X_11596_ _20644_/Q _20608_/Q _11599_/S vssd1 vssd1 vccd1 vccd1 _11596_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16123_ _19586_/Q _16127_/A2 _16127_/B1 vssd1 vssd1 vccd1 vccd1 _16123_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13335_ _19229_/Q _19228_/Q _19227_/Q _13450_/A vssd1 vssd1 vccd1 vccd1 _13403_/B
+ sky130_fd_sc_hd__and4_2
X_10547_ _14524_/B1 _10546_/X _10544_/X vssd1 vssd1 vccd1 vccd1 _10547_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13266_ _19235_/Q _13365_/B _19236_/Q vssd1 vssd1 vccd1 vccd1 _13266_/Y sky130_fd_sc_hd__a21oi_2
X_16054_ _16054_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16054_/Y sky130_fd_sc_hd__nor2_1
X_10478_ _10476_/X _10477_/X _11250_/S vssd1 vssd1 vccd1 vccd1 _10478_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15005_ input280/X _15133_/B _15012_/B _14988_/B vssd1 vssd1 vccd1 vccd1 _15005_/X
+ sky130_fd_sc_hd__a211o_1
X_12217_ _09503_/A _20718_/Q _12375_/S _12216_/X vssd1 vssd1 vccd1 vccd1 _12217_/X
+ sky130_fd_sc_hd__a31o_1
X_13197_ _20970_/Q _13397_/B vssd1 vssd1 vccd1 vccd1 _13197_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19813_ _20692_/CLK _19813_/D vssd1 vssd1 vccd1 vccd1 _19813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12148_ _20050_/Q _19925_/Q _12148_/S vssd1 vssd1 vccd1 vccd1 _12148_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19744_ _20795_/CLK _19744_/D vssd1 vssd1 vccd1 vccd1 _19744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16956_ _19240_/Q _16980_/A2 _16980_/B1 _19109_/Q _16955_/X vssd1 vssd1 vccd1 vccd1
+ _16956_/X sky130_fd_sc_hd__o221a_2
X_12079_ _12084_/A _19328_/Q _12084_/C vssd1 vssd1 vccd1 vccd1 _12079_/X sky130_fd_sc_hd__or3_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15907_ _20748_/Q _15934_/A2 _15934_/B1 _20780_/Q vssd1 vssd1 vccd1 vccd1 _15907_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19675_ _20180_/CLK _19675_/D vssd1 vssd1 vccd1 vccd1 _19675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16887_ _16887_/A _16887_/B vssd1 vssd1 vccd1 vccd1 _16887_/Y sky130_fd_sc_hd__nor2_1
XFILLER_253_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18626_ _18877_/A _18626_/B vssd1 vssd1 vccd1 vccd1 _20929_/D sky130_fd_sc_hd__nor2_1
XFILLER_280_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_266_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _15890_/B _15821_/Y _15837_/X _15976_/B2 vssd1 vssd1 vccd1 vccd1 _15838_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18557_ _20912_/Q fanout750/X _18556_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18558_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_280_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15769_ _19723_/Q _15961_/A2 _15961_/B1 _19755_/Q vssd1 vssd1 vccd1 vccd1 _15769_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17508_ _20289_/Q _17524_/B vssd1 vssd1 vccd1 vccd1 _17508_/Y sky130_fd_sc_hd__nand2_1
X_18488_ _20889_/Q fanout753/X _18487_/X _18491_/B2 vssd1 vssd1 vccd1 vccd1 _18489_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_14 _15480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ _20265_/Q _20264_/Q _17457_/C _17421_/Y vssd1 vssd1 vccd1 vccd1 _17439_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_25 _15671_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_36 _16049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _16876_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 _17011_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20450_ _20714_/CLK _20450_/D vssd1 vssd1 vccd1 vccd1 _20450_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_69 _09501_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19109_ _20273_/CLK _19109_/D vssd1 vssd1 vccd1 vccd1 _19109_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20381_ _20573_/CLK _20381_/D vssd1 vssd1 vccd1 vccd1 _20381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_99_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20763_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_28_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20667_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21002_ _21010_/CLK _21002_/D vssd1 vssd1 vccd1 vccd1 _21002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09626_ _14668_/B _09689_/C vssd1 vssd1 vccd1 vccd1 _09630_/C sky130_fd_sc_hd__xnor2_1
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_270_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09557_ _19179_/Q _11367_/A _12519_/A vssd1 vssd1 vccd1 vccd1 _09561_/C sky130_fd_sc_hd__or3_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09488_ _09488_/A vssd1 vssd1 vccd1 vccd1 _09488_/Y sky130_fd_sc_hd__inv_4
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20717_ _20717_/CLK _20717_/D vssd1 vssd1 vccd1 vccd1 _20717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11450_ _12144_/C1 _11439_/X _11442_/X _11449_/X _12152_/A1 vssd1 vssd1 vccd1 vccd1
+ _11450_/X sky130_fd_sc_hd__a311o_2
X_20648_ _20717_/CLK _20648_/D vssd1 vssd1 vccd1 vccd1 _20648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ _10399_/X _10400_/X _12426_/S vssd1 vssd1 vccd1 vccd1 _10401_/X sky130_fd_sc_hd__mux2_1
X_11381_ _12427_/A1 _20373_/Q _20437_/Q _12428_/S vssd1 vssd1 vccd1 vccd1 _11381_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20579_ _20579_/CLK _20579_/D vssd1 vssd1 vccd1 vccd1 _20579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _13009_/Y _13120_/B vssd1 vssd1 vccd1 vccd1 _13121_/B sky130_fd_sc_hd__nand2b_1
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10332_ _19879_/Q _10345_/S vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__or2_1
XFILLER_164_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13051_ _20952_/Q _20886_/Q vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__and2_1
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _19813_/Q _11192_/A2 _10261_/X _15129_/A0 _10262_/X vssd1 vssd1 vccd1 vccd1
+ _10263_/X sky130_fd_sc_hd__o221a_1
Xfanout2003 _16866_/B2 vssd1 vssd1 vccd1 vccd1 _16886_/B2 sky130_fd_sc_hd__buf_4
XFILLER_279_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12002_ _09834_/A _19924_/Q _10622_/S _20049_/Q vssd1 vssd1 vccd1 vccd1 _12002_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_87_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1302 _16982_/B1 vssd1 vssd1 vccd1 vccd1 _16932_/B1 sky130_fd_sc_hd__buf_6
XFILLER_105_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10194_ _12277_/A1 _17899_/A1 _10193_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _15528_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1313 _14853_/S vssd1 vssd1 vccd1 vccd1 _15983_/A sky130_fd_sc_hd__buf_6
Xfanout1324 _12463_/B vssd1 vssd1 vccd1 vccd1 _15258_/A sky130_fd_sc_hd__buf_4
XFILLER_120_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1335 _11392_/A2 vssd1 vssd1 vccd1 vccd1 _12412_/A2 sky130_fd_sc_hd__buf_8
X_16810_ _16846_/A input77/X vssd1 vssd1 vccd1 vccd1 _16810_/Y sky130_fd_sc_hd__nand2_1
Xfanout1346 _17321_/A2 vssd1 vssd1 vccd1 vccd1 _17327_/A2 sky130_fd_sc_hd__buf_2
XFILLER_238_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17790_ _20567_/Q _17930_/A1 _17794_/S vssd1 vssd1 vccd1 vccd1 _20567_/D sky130_fd_sc_hd__mux2_1
Xfanout1357 _16567_/A vssd1 vssd1 vccd1 vccd1 _16551_/A sky130_fd_sc_hd__buf_2
Xfanout1368 _12921_/X vssd1 vssd1 vccd1 vccd1 _14330_/A2 sky130_fd_sc_hd__buf_8
XFILLER_19_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1379 _11947_/S vssd1 vssd1 vccd1 vccd1 _11944_/S sky130_fd_sc_hd__buf_6
XFILLER_47_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16741_ _16822_/A _16741_/B vssd1 vssd1 vccd1 vccd1 _16741_/Y sky130_fd_sc_hd__nor2_1
XFILLER_235_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13953_ _19151_/Q _13953_/A2 _14004_/B1 _13952_/X _16159_/C1 vssd1 vssd1 vccd1 vccd1
+ _19151_/D sky130_fd_sc_hd__o221a_1
XFILLER_281_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19460_ _20719_/CLK _19460_/D vssd1 vssd1 vccd1 vccd1 _19460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12904_ _19522_/Q _12916_/A2 _12903_/X _12916_/B2 vssd1 vssd1 vccd1 vccd1 _12906_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16672_ _16672_/A _17812_/A vssd1 vssd1 vccd1 vccd1 _16673_/C sky130_fd_sc_hd__nor2_1
XFILLER_59_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ _19102_/Q _14738_/B _13889_/B1 _19168_/Q _16171_/A vssd1 vssd1 vccd1 vccd1
+ _19102_/D sky130_fd_sc_hd__o221a_1
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18411_ _20860_/Q _18210_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18412_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ _19542_/Q _16036_/A2 _15621_/X _15622_/X _16167_/C1 vssd1 vssd1 vccd1 vccd1
+ _19542_/D sky130_fd_sc_hd__o221a_1
XFILLER_185_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19391_ _20682_/CLK _19391_/D vssd1 vssd1 vccd1 vccd1 _19391_/Q sky130_fd_sc_hd__dfxtp_1
X_12835_ _12835_/A _12835_/B vssd1 vssd1 vccd1 vccd1 _12835_/Y sky130_fd_sc_hd__nor2_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _20826_/Q _18343_/B _18341_/Y _18708_/A vssd1 vssd1 vccd1 vccd1 _20826_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _14815_/S _15548_/Y _15553_/X vssd1 vssd1 vccd1 vccd1 _15554_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _19504_/Q _12786_/B vssd1 vssd1 vccd1 vccd1 _12767_/B sky130_fd_sc_hd__and2_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14505_ _19283_/Q _17202_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19283_/D sky130_fd_sc_hd__mux2_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _19550_/Q _18308_/B vssd1 vssd1 vccd1 vccd1 _18273_/Y sky130_fd_sc_hd__nand2b_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _09834_/A _19816_/Q _19320_/Q _10622_/S vssd1 vssd1 vccd1 vccd1 _11717_/X
+ sky130_fd_sc_hd__a22o_1
X_15485_ _19713_/Q _15454_/S _15484_/X vssd1 vssd1 vccd1 vccd1 _15485_/X sky130_fd_sc_hd__o21a_1
X_12697_ _12698_/C _12698_/D vssd1 vssd1 vccd1 vccd1 _13544_/B sky130_fd_sc_hd__nor2_2
X_17224_ _18134_/A _17224_/B vssd1 vssd1 vccd1 vccd1 _17224_/X sky130_fd_sc_hd__or2_1
X_14436_ _09488_/A _14435_/Y _13100_/A vssd1 vssd1 vccd1 vccd1 _14437_/C sky130_fd_sc_hd__o21a_1
X_11648_ _15713_/A vssd1 vssd1 vccd1 vccd1 _11648_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 core_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_4
Xinput23 core_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_4
Xinput34 core_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_4
X_17155_ _20121_/Q _17189_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20121_/D sky130_fd_sc_hd__mux2_1
Xinput45 dout0[11] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_2
X_14367_ _14427_/A _14367_/B vssd1 vssd1 vccd1 vccd1 _14367_/Y sky130_fd_sc_hd__nor2_1
X_11579_ _12051_/A1 _19481_/Q _19449_/Q _11978_/S _12123_/C1 vssd1 vssd1 vccd1 vccd1
+ _11579_/X sky130_fd_sc_hd__a221o_1
Xinput56 dout0[21] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_2
Xinput67 dout0[31] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_2
X_16106_ _10463_/X _16106_/A2 _16105_/X vssd1 vssd1 vccd1 vccd1 _19577_/D sky130_fd_sc_hd__o21a_1
Xinput78 dout0[41] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_2
Xinput89 dout0[51] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_2
X_13318_ _20958_/Q _13607_/B _13316_/X _13317_/Y _18462_/A vssd1 vssd1 vccd1 vccd1
+ _13318_/Y sky130_fd_sc_hd__a221oi_4
X_17086_ _20056_/Q _17679_/A1 _17114_/S vssd1 vssd1 vccd1 vccd1 _20056_/D sky130_fd_sc_hd__mux2_1
X_14298_ _20284_/Q _14330_/A2 _14330_/B1 input224/X vssd1 vssd1 vccd1 vccd1 _14300_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16037_ _16037_/A _16037_/B vssd1 vssd1 vccd1 vccd1 _16037_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13249_ _13362_/B _13362_/C _13362_/A vssd1 vssd1 vccd1 vccd1 _13249_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_254_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17988_ _20734_/Q _17991_/C vssd1 vssd1 vccd1 vccd1 _17989_/B sky130_fd_sc_hd__and2_1
XFILLER_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19727_ _19970_/CLK _19727_/D vssd1 vssd1 vccd1 vccd1 _19727_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_284_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1880 _19163_/Q vssd1 vssd1 vccd1 vccd1 _12464_/A sky130_fd_sc_hd__buf_12
X_16939_ _16981_/A1 _15834_/X _16879_/X _16938_/X vssd1 vssd1 vccd1 vccd1 _16939_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_266_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1891 _16185_/A vssd1 vssd1 vccd1 vccd1 _16187_/A sky130_fd_sc_hd__buf_4
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19658_ _20410_/CLK _19658_/D vssd1 vssd1 vccd1 vccd1 _19658_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_146_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19511_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_281_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18609_ _18499_/X _18621_/A2 _18607_/Y _18608_/Y vssd1 vssd1 vccd1 vccd1 _18610_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_53_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19589_ _19589_/CLK _19589_/D vssd1 vssd1 vccd1 vccd1 _19589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20502_ _20675_/CLK _20502_/D vssd1 vssd1 vccd1 vccd1 _20502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20433_ _20465_/CLK _20433_/D vssd1 vssd1 vccd1 vccd1 _20433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20364_ _20688_/CLK _20364_/D vssd1 vssd1 vccd1 vccd1 _20364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20295_ _20296_/CLK _20295_/D vssd1 vssd1 vccd1 vccd1 _20295_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_103_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10950_ _12514_/C _10950_/B vssd1 vssd1 vccd1 vccd1 _10950_/Y sky130_fd_sc_hd__nor2_1
XFILLER_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09609_ _09609_/A _19098_/Q _19096_/Q _12967_/B vssd1 vssd1 vccd1 vccd1 _09610_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10881_ _12277_/A1 _17925_/A1 _10880_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _15267_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _14803_/A1 _12582_/C _12752_/B vssd1 vssd1 vccd1 vccd1 _12786_/B sky130_fd_sc_hd__a21o_4
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12551_ _12551_/A _12551_/B _12551_/C _12551_/D vssd1 vssd1 vccd1 vccd1 _12554_/A
+ sky130_fd_sc_hd__or4_2
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11502_ _20573_/Q _11897_/B _11501_/X _12123_/C1 vssd1 vssd1 vccd1 vccd1 _11502_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15270_ input6/X _15334_/B vssd1 vssd1 vccd1 vccd1 _15270_/X sky130_fd_sc_hd__or2_1
X_12482_ _12579_/D _15220_/B vssd1 vssd1 vccd1 vccd1 _12482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11433_ _11418_/X _11419_/X _12134_/S vssd1 vssd1 vccd1 vccd1 _11433_/X sky130_fd_sc_hd__mux2_1
X_14221_ _14221_/A _14221_/B vssd1 vssd1 vccd1 vccd1 _14221_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14152_ _14148_/B _14151_/Y _14202_/S vssd1 vssd1 vccd1 vccd1 _14152_/X sky130_fd_sc_hd__mux2_1
X_11364_ _12392_/C1 _11353_/X _11356_/X _11363_/X _12400_/A1 vssd1 vssd1 vccd1 vccd1
+ _11364_/X sky130_fd_sc_hd__a311o_1
XFILLER_98_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10315_ _11250_/S _10314_/X _10313_/X _11274_/B2 vssd1 vssd1 vccd1 vccd1 _10315_/X
+ sky130_fd_sc_hd__a211o_1
X_13103_ _13091_/X _13397_/B _13101_/Y _13102_/Y _18651_/B vssd1 vssd1 vccd1 vccd1
+ _13103_/X sky130_fd_sc_hd__o311a_1
X_14083_ _14099_/A _14099_/B _14083_/C vssd1 vssd1 vccd1 vccd1 _14083_/X sky130_fd_sc_hd__or3_1
X_18960_ _18960_/A _18960_/B vssd1 vssd1 vccd1 vccd1 _21008_/D sky130_fd_sc_hd__nor2_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11295_ _20118_/Q _20086_/Q _11295_/S vssd1 vssd1 vccd1 vccd1 _11295_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17911_ _20682_/Q _17911_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20682_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13034_ _20961_/Q _20895_/Q vssd1 vssd1 vccd1 vccd1 _13034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_279_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10246_ _10262_/A _19349_/Q _20704_/Q _11042_/B _11378_/S vssd1 vssd1 vccd1 vccd1
+ _10246_/X sky130_fd_sc_hd__a221o_1
X_18891_ _18891_/A _18891_/B vssd1 vssd1 vccd1 vccd1 _20998_/D sky130_fd_sc_hd__nor2_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1110 _17877_/A1 vssd1 vssd1 vccd1 vccd1 _17805_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_152_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1121 _17871_/A1 vssd1 vssd1 vccd1 vccd1 _17939_/A1 sky130_fd_sc_hd__buf_4
Xfanout1132 _17859_/A1 vssd1 vssd1 vccd1 vccd1 _17684_/A1 sky130_fd_sc_hd__buf_4
XFILLER_154_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17842_ _20617_/Q _17914_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20617_/D sky130_fd_sc_hd__mux2_1
X_10177_ _20474_/Q _11303_/S _09730_/A vssd1 vssd1 vccd1 vccd1 _10177_/X sky130_fd_sc_hd__o21a_1
XFILLER_267_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1143 _09936_/A2 vssd1 vssd1 vccd1 vccd1 _17907_/A1 sky130_fd_sc_hd__buf_2
XFILLER_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1154 _09632_/Y vssd1 vssd1 vccd1 vccd1 _13670_/A1 sky130_fd_sc_hd__buf_8
XFILLER_267_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1165 _15096_/Y vssd1 vssd1 vccd1 vccd1 _15673_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1176 _12558_/Y vssd1 vssd1 vccd1 vccd1 _13730_/B sky130_fd_sc_hd__buf_4
XFILLER_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17773_ _20552_/Q _17913_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20552_/D sky130_fd_sc_hd__mux2_1
XFILLER_248_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14985_ _14988_/B vssd1 vssd1 vccd1 vccd1 _14986_/C sky130_fd_sc_hd__inv_2
Xfanout1187 _09686_/Y vssd1 vssd1 vccd1 vccd1 _11246_/A1 sky130_fd_sc_hd__buf_6
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1198 _17234_/X vssd1 vssd1 vccd1 vccd1 _17302_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_281_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19512_ _20913_/CLK _19512_/D vssd1 vssd1 vccd1 vccd1 _19512_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_281_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16724_ _16708_/Y _17219_/B _16722_/X _12952_/X vssd1 vssd1 vccd1 vccd1 _16724_/X
+ sky130_fd_sc_hd__a31o_1
X_13936_ _19140_/Q _13941_/B _13946_/B1 _13412_/A vssd1 vssd1 vccd1 vccd1 _19140_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_75_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19443_ _20570_/CLK _19443_/D vssd1 vssd1 vccd1 vccd1 _19443_/Q sky130_fd_sc_hd__dfxtp_1
X_16655_ _19912_/Q _17099_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19912_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13867_ _13867_/A _13902_/B vssd1 vssd1 vccd1 vccd1 _13867_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15606_ _15606_/A1 _15595_/X _15605_/X vssd1 vssd1 vccd1 vccd1 _16869_/B sky130_fd_sc_hd__a21oi_4
XFILLER_250_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19374_ _20658_/CLK _19374_/D vssd1 vssd1 vccd1 vccd1 _19374_/Q sky130_fd_sc_hd__dfxtp_1
X_12818_ _12483_/Y _12817_/X _15822_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12818_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16586_ _19859_/Q _16592_/A2 _16592_/B1 input30/X vssd1 vssd1 vccd1 vccd1 _16587_/B
+ sky130_fd_sc_hd__o22a_1
X_13798_ _13798_/A1 _13826_/A1 _13735_/B _13826_/B1 input244/X vssd1 vssd1 vccd1 vccd1
+ _13798_/X sky130_fd_sc_hd__a32o_1
X_18325_ _18459_/B _18341_/B vssd1 vssd1 vccd1 vccd1 _18325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15537_ input268/X _15013_/Y _15531_/X _15606_/A1 vssd1 vssd1 vccd1 vccd1 _15537_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12749_ _12749_/A _12749_/B _12749_/C _12748_/B vssd1 vssd1 vccd1 vccd1 _12791_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18256_ _20805_/Q _18255_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18257_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15468_ _15468_/A _15468_/B vssd1 vssd1 vccd1 vccd1 _15468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17207_ _20171_/Q _17801_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20171_/D sky130_fd_sc_hd__mux2_1
XFILLER_200_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14419_ _14437_/A _14437_/B _14419_/C vssd1 vssd1 vccd1 vccd1 _14419_/X sky130_fd_sc_hd__or3_1
X_18187_ _18708_/A _18187_/B vssd1 vssd1 vccd1 vccd1 _20791_/D sky130_fd_sc_hd__and2_1
X_15399_ _16133_/C _15397_/Y _15398_/X _15369_/A _15442_/A vssd1 vssd1 vccd1 vccd1
+ _15399_/X sky130_fd_sc_hd__a32o_1
XFILLER_265_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17138_ _20106_/Q _17800_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20106_/D sky130_fd_sc_hd__mux2_1
XFILLER_171_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09960_ _20138_/Q _20106_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__mux2_1
X_17069_ _20041_/Q _17871_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20041_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20080_ _20647_/CLK _20080_/D vssd1 vssd1 vccd1 vccd1 _20080_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _20646_/Q _20610_/Q _12146_/S vssd1 vssd1 vccd1 vccd1 _09891_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_281_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20982_ _20982_/CLK _20982_/D vssd1 vssd1 vccd1 vccd1 _20982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_43_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20570_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_194_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20416_ _20706_/CLK _20416_/D vssd1 vssd1 vccd1 vccd1 _20416_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20347_ _20635_/CLK _20347_/D vssd1 vssd1 vccd1 vccd1 _20347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10100_ _10098_/X _10099_/X _12082_/S vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__mux2_1
XFILLER_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11080_ _12310_/C1 _11079_/X _11076_/X _12385_/C1 vssd1 vssd1 vccd1 vccd1 _11080_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_89_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20278_ _21016_/CLK _20278_/D vssd1 vssd1 vccd1 vccd1 _20278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput202 localMemory_wb_adr_i[20] vssd1 vssd1 vccd1 vccd1 _12928_/B sky130_fd_sc_hd__clkbuf_2
X_10031_ _09643_/A _09636_/B _11236_/A _10029_/Y vssd1 vssd1 vccd1 vccd1 _10465_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput213 localMemory_wb_adr_i[9] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__clkbuf_2
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput224 localMemory_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_hd__buf_12
XFILLER_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput235 localMemory_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_hd__buf_12
XFILLER_237_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput246 localMemory_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_hd__buf_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput257 manufacturerID[3] vssd1 vssd1 vccd1 vccd1 _17248_/A sky130_fd_sc_hd__buf_2
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput268 partID[13] vssd1 vssd1 vccd1 vccd1 input268/X sky130_fd_sc_hd__clkbuf_2
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput279 partID[9] vssd1 vssd1 vccd1 vccd1 _17299_/A sky130_fd_sc_hd__clkbuf_2
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_263_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ _19132_/Q _14774_/A2 _14769_/X _14772_/C1 vssd1 vssd1 vccd1 vccd1 _19509_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11982_ _12137_/A1 _11973_/X _11981_/X _12137_/C1 vssd1 vssd1 vccd1 vccd1 _11982_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_91_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13721_ _13780_/A _13721_/B vssd1 vssd1 vccd1 vccd1 _13721_/X sky130_fd_sc_hd__and2_1
XFILLER_260_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10933_ _10931_/X _10932_/Y _11313_/B vssd1 vssd1 vccd1 vccd1 _10933_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_56_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16440_ _19760_/Q _16442_/C _16439_/Y vssd1 vssd1 vccd1 vccd1 _19760_/D sky130_fd_sc_hd__o21a_1
X_10864_ _20466_/Q _20306_/Q _12352_/S vssd1 vssd1 vccd1 vccd1 _10864_/X sky130_fd_sc_hd__mux2_1
X_13652_ _13663_/A _13663_/B _13685_/B vssd1 vssd1 vccd1 vccd1 _13652_/X sky130_fd_sc_hd__and3_4
XFILLER_260_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _19506_/Q _12754_/A vssd1 vssd1 vccd1 vccd1 _12740_/B sky130_fd_sc_hd__and2_2
X_16371_ _18126_/A _16371_/B _16372_/B vssd1 vssd1 vccd1 vccd1 _19734_/D sky130_fd_sc_hd__nor3_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10785_/X _10794_/Y _11201_/A _10777_/X vssd1 vssd1 vccd1 vccd1 _10795_/X
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_223_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13583_ _13581_/Y _13582_/Y _18598_/A vssd1 vssd1 vccd1 vccd1 _13583_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18110_ _18112_/A _18110_/B _18111_/B vssd1 vssd1 vccd1 vccd1 _20778_/D sky130_fd_sc_hd__nor3_1
X_15322_ _15322_/A _15322_/B _15322_/C vssd1 vssd1 vccd1 vccd1 _15322_/X sky130_fd_sc_hd__or3_2
XFILLER_158_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _20721_/CLK _19090_/D vssd1 vssd1 vccd1 vccd1 _19090_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _20870_/Q _12549_/B _12534_/C vssd1 vssd1 vccd1 vccd1 _12550_/A sky130_fd_sc_hd__and3_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18041_ _20752_/Q _18039_/B _18040_/Y vssd1 vssd1 vccd1 vccd1 _20752_/D sky130_fd_sc_hd__o21a_1
XFILLER_200_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15253_ _15545_/A _15545_/B vssd1 vssd1 vccd1 vccd1 _15253_/X sky130_fd_sc_hd__or2_1
XFILLER_149_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12465_ _14895_/A _15026_/A vssd1 vssd1 vccd1 vccd1 _12465_/X sky130_fd_sc_hd__and2_4
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14204_ _14204_/A _14204_/B _14204_/C vssd1 vssd1 vccd1 vccd1 _14204_/X sky130_fd_sc_hd__or3_1
X_11416_ _10277_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _11416_/Y sky130_fd_sc_hd__nand2b_1
X_12396_ _12396_/A1 _19927_/Q _12395_/S _12379_/X vssd1 vssd1 vccd1 vccd1 _12396_/X
+ sky130_fd_sc_hd__o211a_1
X_15184_ _15179_/X _15184_/B _15220_/A vssd1 vssd1 vccd1 vccd1 _15187_/B sky130_fd_sc_hd__and3b_1
XFILLER_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11347_ _09502_/A _11345_/X _11346_/X _12311_/C1 vssd1 vssd1 vccd1 vccd1 _11347_/X
+ sky130_fd_sc_hd__a211o_1
X_14135_ _19216_/Q _14256_/A2 _14134_/X _18698_/A vssd1 vssd1 vccd1 vccd1 _19216_/D
+ sky130_fd_sc_hd__o211a_1
X_19992_ _19992_/CLK _19992_/D vssd1 vssd1 vccd1 vccd1 _19992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14066_ _19192_/Q _14082_/A2 _14065_/X _16087_/B1 vssd1 vssd1 vccd1 vccd1 _19192_/D
+ sky130_fd_sc_hd__o211a_1
X_11278_ _12402_/A1 _17852_/A1 _11277_/X _13675_/A vssd1 vssd1 vccd1 vccd1 _13641_/B
+ sky130_fd_sc_hd__o211a_1
X_18943_ _18667_/Y _18970_/A2 _18941_/Y _18942_/Y vssd1 vssd1 vccd1 vccd1 _18943_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10229_ _20412_/Q _20348_/Q _10986_/B vssd1 vssd1 vccd1 vccd1 _10229_/X sky130_fd_sc_hd__mux2_1
X_13017_ _20970_/Q _20904_/Q vssd1 vssd1 vccd1 vccd1 _13017_/Y sky130_fd_sc_hd__nor2_2
XFILLER_140_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18874_ _18628_/Y _18977_/A2 _18872_/Y _18873_/Y vssd1 vssd1 vccd1 vccd1 _18874_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17825_ _20600_/Q split4/X _17840_/S vssd1 vssd1 vccd1 vccd1 _20600_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17756_ _20535_/Q _17896_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20535_/D sky130_fd_sc_hd__mux2_1
X_14968_ _15314_/D _14987_/A vssd1 vssd1 vccd1 vccd1 _14972_/B sky130_fd_sc_hd__nor2_2
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16707_ _20020_/Q _16706_/X _13466_/B vssd1 vssd1 vccd1 vccd1 _16707_/X sky130_fd_sc_hd__o21ba_4
XFILLER_251_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13919_ _19125_/Q _13583_/Y _13919_/S vssd1 vssd1 vccd1 vccd1 _13920_/B sky130_fd_sc_hd__mux2_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17687_ _20471_/Q _17687_/A1 _17706_/S vssd1 vssd1 vccd1 vccd1 _20471_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14899_ _16720_/A _14899_/B vssd1 vssd1 vccd1 vccd1 _18136_/B sky130_fd_sc_hd__nand2_1
X_19426_ _20585_/CLK _19426_/D vssd1 vssd1 vccd1 vccd1 _19426_/Q sky130_fd_sc_hd__dfxtp_1
X_16638_ _17082_/A _17918_/A vssd1 vssd1 vccd1 vccd1 _16639_/C sky130_fd_sc_hd__nor2_1
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19357_ _20712_/CLK _19357_/D vssd1 vssd1 vccd1 vccd1 _19357_/Q sky130_fd_sc_hd__dfxtp_1
X_16569_ _16593_/A _16569_/B vssd1 vssd1 vccd1 vccd1 _19850_/D sky130_fd_sc_hd__or2_1
XFILLER_204_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18308_ _19557_/Q _18308_/B vssd1 vssd1 vccd1 vccd1 _18308_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19288_ _20641_/CLK _19288_/D vssd1 vssd1 vccd1 vccd1 _19288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18239_ _18248_/B _14281_/B _18238_/Y vssd1 vssd1 vccd1 vccd1 _18514_/B sky130_fd_sc_hd__o21ai_4
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20201_ _20727_/CLK _20201_/D vssd1 vssd1 vccd1 vccd1 _20201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20132_ _20703_/CLK _20132_/D vssd1 vssd1 vccd1 vccd1 _20132_/Q sky130_fd_sc_hd__dfxtp_1
X_09943_ input119/X input154/X _11241_/S vssd1 vssd1 vccd1 vccd1 _09943_/X sky130_fd_sc_hd__mux2_8
Xfanout903 _15939_/A2 vssd1 vssd1 vccd1 vccd1 _16045_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout914 _16041_/B1 vssd1 vssd1 vccd1 vccd1 _15445_/B1 sky130_fd_sc_hd__buf_4
XFILLER_225_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout925 _15595_/B1 vssd1 vssd1 vccd1 vccd1 _15475_/B1 sky130_fd_sc_hd__buf_6
XFILLER_86_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout936 _11223_/A vssd1 vssd1 vccd1 vccd1 _15170_/A sky130_fd_sc_hd__clkbuf_4
X_20063_ _20706_/CLK _20063_/D vssd1 vssd1 vccd1 vccd1 _20063_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout947 _15118_/S vssd1 vssd1 vccd1 vccd1 _15578_/S sky130_fd_sc_hd__buf_6
X_09874_ _20578_/Q _11897_/B vssd1 vssd1 vccd1 vccd1 _09874_/X sky130_fd_sc_hd__or2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_161_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21027_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout958 _11397_/A2 vssd1 vssd1 vccd1 vccd1 _17788_/A1 sky130_fd_sc_hd__buf_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout969 _10474_/X vssd1 vssd1 vccd1 vccd1 _17896_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_307 input234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_318 _13613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_329 _20259_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20965_ _21011_/CLK _20965_/D vssd1 vssd1 vccd1 vccd1 _20965_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _21024_/CLK _20896_/D vssd1 vssd1 vccd1 vccd1 _20896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10580_ _20406_/Q _20342_/Q _11676_/S vssd1 vssd1 vccd1 vccd1 _10580_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12250_ _19827_/Q _12255_/A2 _12248_/X _09738_/A _12249_/X vssd1 vssd1 vccd1 vccd1
+ _12250_/X sky130_fd_sc_hd__o221a_1
XFILLER_166_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11201_/X sky130_fd_sc_hd__or2_2
XFILLER_135_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _12186_/S _12181_/B vssd1 vssd1 vccd1 vccd1 _12181_/X sky130_fd_sc_hd__or2_1
XFILLER_253_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11132_ _11201_/A _11114_/X _11122_/X _11131_/Y vssd1 vssd1 vccd1 vccd1 _11132_/X
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ _10127_/A _11058_/Y _11062_/X _11056_/X vssd1 vssd1 vccd1 vccd1 _11063_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15940_ _16017_/C1 _15939_/X _15935_/X vssd1 vssd1 vccd1 vccd1 _15940_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _19514_/Q _15741_/A _11649_/S vssd1 vssd1 vccd1 vccd1 _11742_/B sky130_fd_sc_hd__mux2_8
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15871_ _19727_/Q _15961_/A2 _15961_/B1 _19759_/Q vssd1 vssd1 vccd1 vccd1 _15871_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ _20366_/Q _17678_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20366_/D sky130_fd_sc_hd__mux2_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14822_ _10016_/B _10641_/B _14822_/S vssd1 vssd1 vccd1 vccd1 _14822_/X sky130_fd_sc_hd__mux2_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _18483_/X _18621_/A2 _18588_/Y _18589_/Y vssd1 vssd1 vccd1 vccd1 _18591_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _20301_/Q _17780_/A1 _17570_/S vssd1 vssd1 vccd1 vccd1 _20301_/D sky130_fd_sc_hd__mux2_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14753_ _19501_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14753_/X sky130_fd_sc_hd__or2_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _20552_/Q _11965_/B vssd1 vssd1 vccd1 vccd1 _11965_/X sky130_fd_sc_hd__or2_1
XFILLER_251_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13704_ _13740_/A _13666_/B _13665_/A _15076_/A vssd1 vssd1 vccd1 vccd1 _13704_/X
+ sky130_fd_sc_hd__a22o_1
X_10916_ _19666_/Q _11342_/S _10915_/X _11338_/A1 vssd1 vssd1 vccd1 vccd1 _10916_/X
+ sky130_fd_sc_hd__o211a_1
X_17472_ _20271_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17472_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14684_ _19443_/Q _17933_/A1 _14702_/S vssd1 vssd1 vccd1 vccd1 _19443_/D sky130_fd_sc_hd__mux2_1
X_11896_ _20550_/Q _11915_/S vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__or2_1
X_19211_ _20426_/CLK _19211_/D vssd1 vssd1 vccd1 vccd1 _19211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16423_ _19754_/Q _16426_/C _18104_/A vssd1 vssd1 vccd1 vccd1 _16423_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_204_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13635_ _13635_/A _13740_/B vssd1 vssd1 vccd1 vccd1 _13637_/C sky130_fd_sc_hd__or2_1
X_10847_ _10832_/X _10846_/X _12401_/A1 vssd1 vssd1 vccd1 vccd1 _10847_/X sky130_fd_sc_hd__a21o_2
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19142_ _19520_/CLK _19142_/D vssd1 vssd1 vccd1 vccd1 _19142_/Q sky130_fd_sc_hd__dfxtp_1
X_16354_ _19727_/Q _19728_/Q _16354_/C vssd1 vssd1 vccd1 vccd1 _16356_/B sky130_fd_sc_hd__and3_1
XFILLER_201_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13566_ _13556_/Y _13565_/X _17952_/A vssd1 vssd1 vccd1 vccd1 _13566_/Y sky130_fd_sc_hd__a21oi_4
X_10778_ _20371_/Q _20435_/Q _12268_/S vssd1 vssd1 vccd1 vccd1 _10778_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15305_ _19708_/Q _15475_/A2 _15475_/B1 _19740_/Q vssd1 vssd1 vccd1 vccd1 _15305_/X
+ sky130_fd_sc_hd__a22o_1
X_12517_ _13897_/A _12517_/B _12517_/C vssd1 vssd1 vccd1 vccd1 _12518_/C sky130_fd_sc_hd__or3_1
X_19073_ _20418_/Q vssd1 vssd1 vccd1 vccd1 _20418_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16285_ _18054_/A _19702_/Q vssd1 vssd1 vccd1 vccd1 _19702_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13497_ _13631_/B _15185_/A vssd1 vssd1 vccd1 vccd1 _13497_/Y sky130_fd_sc_hd__nor2_2
X_18024_ _20747_/Q _20746_/Q _18024_/C vssd1 vssd1 vccd1 vccd1 _18030_/C sky130_fd_sc_hd__and3_1
X_15236_ _20950_/Q _15322_/C _15568_/B1 _20822_/Q _15235_/X vssd1 vssd1 vccd1 vccd1
+ _15236_/X sky130_fd_sc_hd__a221o_1
XFILLER_173_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ _12450_/A _12449_/C _12447_/A vssd1 vssd1 vccd1 vccd1 _12469_/S sky130_fd_sc_hd__a21o_1
XFILLER_154_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15167_ _15043_/X _15059_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15168_/A sky130_fd_sc_hd__mux2_1
X_12379_ _20052_/Q _12397_/S vssd1 vssd1 vccd1 vccd1 _12379_/X sky130_fd_sc_hd__or2_1
XFILLER_181_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14118_ _20266_/Q _14237_/A2 _14216_/B1 input215/X vssd1 vssd1 vccd1 vccd1 _14123_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_141_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19975_ _19978_/CLK _19975_/D vssd1 vssd1 vccd1 vccd1 _19975_/Q sky130_fd_sc_hd__dfxtp_1
X_15098_ _16133_/C _15094_/Y _15097_/X _12562_/A _15442_/A vssd1 vssd1 vccd1 vccd1
+ _15098_/X sky130_fd_sc_hd__a32o_1
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14049_ _14081_/A _14069_/B _14049_/C vssd1 vssd1 vccd1 vccd1 _14049_/X sky130_fd_sc_hd__or3_1
X_18926_ _19108_/Q _18954_/A2 _18967_/B1 _15843_/A vssd1 vssd1 vccd1 vccd1 _18927_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18857_ _19098_/Q _18864_/A2 _18864_/B1 _13426_/B vssd1 vssd1 vccd1 vccd1 _18858_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09590_ _19098_/Q _12967_/B _09609_/A vssd1 vssd1 vccd1 vccd1 _09592_/C sky130_fd_sc_hd__o21bai_4
X_17808_ _20585_/Q _17948_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20585_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18788_ _18470_/Y _20983_/Q _18819_/B vssd1 vssd1 vccd1 vccd1 _18788_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17739_ _20520_/Q _17913_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20520_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20750_ _20751_/CLK _20750_/D vssd1 vssd1 vccd1 vccd1 _20750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19409_ _20568_/CLK _19409_/D vssd1 vssd1 vccd1 vccd1 _19409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20681_ _20681_/CLK _20681_/D vssd1 vssd1 vccd1 vccd1 _20681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout700 _13855_/Y vssd1 vssd1 vccd1 vccd1 _14107_/A sky130_fd_sc_hd__buf_4
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20115_ _20179_/CLK _20115_/D vssd1 vssd1 vccd1 vccd1 _20115_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1709 _11378_/S vssd1 vssd1 vccd1 vccd1 _12419_/C1 sky130_fd_sc_hd__buf_6
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout711 _16279_/B vssd1 vssd1 vccd1 vccd1 _13822_/A1 sky130_fd_sc_hd__buf_4
XFILLER_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09926_ _09776_/S _09921_/Y _09925_/Y _12020_/C1 vssd1 vssd1 vccd1 vccd1 _09926_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout722 _13480_/Y vssd1 vssd1 vccd1 vccd1 _13775_/A sky130_fd_sc_hd__buf_8
Xfanout733 _18997_/B vssd1 vssd1 vccd1 vccd1 _19015_/B sky130_fd_sc_hd__buf_6
XFILLER_120_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout744 _18818_/A2 vssd1 vssd1 vccd1 vccd1 _18977_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_277_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout755 _18937_/B vssd1 vssd1 vccd1 vccd1 _18964_/B sky130_fd_sc_hd__buf_6
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20046_ _20681_/CLK _20046_/D vssd1 vssd1 vccd1 vccd1 _20046_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout766 _18593_/A2 vssd1 vssd1 vccd1 vccd1 _18767_/A sky130_fd_sc_hd__buf_6
XFILLER_219_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09857_ _12107_/A1 _09790_/X _09856_/X _11397_/B2 vssd1 vssd1 vccd1 vccd1 _15795_/A
+ sky130_fd_sc_hd__a22o_4
Xfanout777 _18616_/B vssd1 vssd1 vccd1 vccd1 _18612_/B sky130_fd_sc_hd__buf_4
XFILLER_246_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout788 _12525_/Y vssd1 vssd1 vccd1 vccd1 _13323_/C sky130_fd_sc_hd__buf_6
XFILLER_86_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout799 _12479_/A vssd1 vssd1 vccd1 vccd1 split8/A sky130_fd_sc_hd__buf_12
XFILLER_273_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09788_ _19581_/Q _09787_/X _11229_/S vssd1 vssd1 vccd1 vccd1 _10285_/A sky130_fd_sc_hd__mux2_2
XFILLER_234_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_104 _12978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_115 _16235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _13656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_137 _13687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _13750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11794_/B _11794_/C _13420_/A vssd1 vssd1 vccd1 vccd1 _15652_/A sky130_fd_sc_hd__a21o_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20949_/CLK _20948_/D vssd1 vssd1 vccd1 vccd1 _20948_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _13780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10701_ _19872_/Q _19773_/Q _12268_/S vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11681_ _20040_/Q _19915_/Q _11682_/S vssd1 vssd1 vccd1 vccd1 _11681_/X sky130_fd_sc_hd__mux2_1
X_20879_ _21041_/CLK _20879_/D vssd1 vssd1 vccd1 vccd1 _20879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13420_ _13420_/A _13420_/B vssd1 vssd1 vccd1 vccd1 _13427_/B sky130_fd_sc_hd__xnor2_4
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10632_ _10409_/A _10624_/X _10627_/X _10631_/X vssd1 vssd1 vccd1 vccd1 _10632_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_197_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10563_ _20470_/Q _20310_/Q _11994_/S vssd1 vssd1 vccd1 vccd1 _10563_/X sky130_fd_sc_hd__mux2_1
X_13351_ _20930_/Q _13350_/B _18628_/B vssd1 vssd1 vccd1 vccd1 _13352_/C sky130_fd_sc_hd__a21oi_1
XFILLER_167_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12302_ _12298_/X _12301_/X _12302_/S vssd1 vssd1 vccd1 vccd1 _12302_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16070_ _11239_/X _16106_/A2 _16069_/X vssd1 vssd1 vccd1 vccd1 _19559_/D sky130_fd_sc_hd__o21a_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10494_ _11266_/A1 _20667_/Q _09623_/B _10152_/S vssd1 vssd1 vccd1 vccd1 _10494_/X
+ sky130_fd_sc_hd__o31a_1
X_13282_ _12748_/X _13281_/Y _13107_/A vssd1 vssd1 vccd1 vccd1 _13282_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15021_ _15021_/A _15021_/B _15021_/C vssd1 vssd1 vccd1 vccd1 _15021_/X sky130_fd_sc_hd__and3_4
X_12233_ _20426_/Q _12313_/S _12211_/X _12324_/S vssd1 vssd1 vccd1 vccd1 _12233_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12164_ _19394_/Q _20685_/Q _12165_/S vssd1 vssd1 vccd1 vccd1 _12164_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11115_ _20367_/Q _20431_/Q _11116_/S vssd1 vssd1 vccd1 vccd1 _11115_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16972_ _19242_/Q _16980_/A2 _16980_/B1 _19111_/Q _16971_/X vssd1 vssd1 vccd1 vccd1
+ _16972_/X sky130_fd_sc_hd__o221a_2
X_12095_ _12828_/A _12095_/B vssd1 vssd1 vccd1 vccd1 _12095_/Y sky130_fd_sc_hd__nand2_1
X_19760_ _19970_/CLK _19760_/D vssd1 vssd1 vccd1 vccd1 _19760_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11046_ _11375_/S _11041_/X _11045_/X _11384_/S vssd1 vssd1 vccd1 vccd1 _11047_/B
+ sky130_fd_sc_hd__o211a_1
X_18711_ _20956_/Q _18210_/Y _18719_/S vssd1 vssd1 vccd1 vccd1 _18712_/B sky130_fd_sc_hd__mux2_1
X_15923_ _15923_/A _15923_/B _15814_/A vssd1 vssd1 vccd1 vccd1 _15923_/X sky130_fd_sc_hd__or3b_1
XFILLER_265_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19691_ _20179_/CLK _19691_/D vssd1 vssd1 vccd1 vccd1 _19691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18642_ _18891_/A _18642_/B vssd1 vssd1 vccd1 vccd1 _20933_/D sky130_fd_sc_hd__nor2_1
XFILLER_92_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _21036_/Q _21004_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _15854_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _15220_/A _15095_/B vssd1 vssd1 vccd1 vccd1 _15096_/A sky130_fd_sc_hd__and2_2
XFILLER_218_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _20916_/Q _18592_/B vssd1 vssd1 vccd1 vccd1 _18573_/Y sky130_fd_sc_hd__nand2_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _15948_/A1 _12800_/X _15784_/X _15921_/B2 vssd1 vssd1 vccd1 vccd1 _15787_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_224_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12997_ _19242_/Q _19241_/Q _19240_/Q _13231_/B vssd1 vssd1 vccd1 vccd1 _13114_/B
+ sky130_fd_sc_hd__and4_2
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ _20297_/Q _17524_/B vssd1 vssd1 vccd1 vccd1 _17524_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14736_ _19493_/Q _17708_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19493_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11948_ _11948_/A1 _11947_/X _11946_/X vssd1 vssd1 vccd1 vccd1 _11948_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17455_ _17460_/A2 _20264_/Q _16191_/A _17454_/X vssd1 vssd1 vccd1 vccd1 _20264_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _19429_/Q _17951_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19429_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11879_ _13434_/A vssd1 vssd1 vccd1 vccd1 _11880_/B sky130_fd_sc_hd__inv_2
XFILLER_232_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16406_ _19747_/Q _16404_/B _16405_/Y vssd1 vssd1 vccd1 vccd1 _19747_/D sky130_fd_sc_hd__o21a_1
XFILLER_220_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13618_ _13626_/A1 _13411_/B _13426_/A _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13618_/X
+ sky130_fd_sc_hd__a22o_2
X_17386_ _20241_/Q _17337_/B _17530_/A2 _20290_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17386_/X sky130_fd_sc_hd__a221o_1
X_14598_ _19364_/Q _17950_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19364_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19125_ _21021_/CLK _19125_/D vssd1 vssd1 vccd1 vccd1 _19125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16337_ _19721_/Q _16338_/C _19722_/Q vssd1 vssd1 vccd1 vccd1 _16339_/B sky130_fd_sc_hd__a21oi_1
XFILLER_119_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ _13064_/A _13064_/B _13064_/C _13064_/D vssd1 vssd1 vccd1 vccd1 _13549_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19056_ _20401_/Q vssd1 vssd1 vccd1 vccd1 _20401_/D sky130_fd_sc_hd__clkbuf_2
X_16268_ _19684_/Q _17942_/A1 _16272_/S vssd1 vssd1 vccd1 vccd1 _19684_/D sky130_fd_sc_hd__mux2_1
X_18007_ _20740_/Q _18005_/B _18006_/Y vssd1 vssd1 vccd1 vccd1 _20740_/D sky130_fd_sc_hd__o21a_1
Xoutput303 _21046_/X vssd1 vssd1 vccd1 vccd1 clk0 sky130_fd_sc_hd__clkbuf_2
X_15219_ _15220_/A _15220_/B vssd1 vssd1 vccd1 vccd1 _15219_/Y sky130_fd_sc_hd__nor2_8
XFILLER_127_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput314 _13621_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[18] sky130_fd_sc_hd__buf_4
X_16199_ _16605_/A _17574_/B _16199_/C vssd1 vssd1 vccd1 vccd1 _16199_/X sky130_fd_sc_hd__and3_4
XFILLER_173_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput325 _13494_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[2] sky130_fd_sc_hd__buf_4
XFILLER_99_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput336 _13683_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[11] sky130_fd_sc_hd__buf_4
XFILLER_99_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput347 _13729_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[21] sky130_fd_sc_hd__buf_4
Xoutput358 _13780_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[31] sky130_fd_sc_hd__buf_4
Xoutput369 _13640_/X vssd1 vssd1 vccd1 vccd1 core_wb_sel_o[3] sky130_fd_sc_hd__buf_4
XFILLER_259_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19958_ _20662_/CLK _19958_/D vssd1 vssd1 vccd1 vccd1 _19958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09711_ _20648_/Q _20612_/Q _11965_/B vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__mux2_1
X_18909_ _18647_/Y _18970_/A2 _18907_/Y _18908_/Y vssd1 vssd1 vccd1 vccd1 _18909_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_274_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19889_ _20713_/CLK _19889_/D vssd1 vssd1 vccd1 vccd1 _19889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_255_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09642_ _11234_/A _09684_/A _09638_/Y _09641_/X vssd1 vssd1 vccd1 vccd1 _09686_/D
+ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_271_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09573_ _12708_/A _11922_/A1 _16063_/B2 vssd1 vssd1 vccd1 vccd1 _09573_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20802_ _20990_/CLK _20802_/D vssd1 vssd1 vccd1 vccd1 _20802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20733_ _20766_/CLK _20733_/D vssd1 vssd1 vccd1 vccd1 _20733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20664_ _20664_/CLK _20664_/D vssd1 vssd1 vccd1 vccd1 _20664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20595_ _20663_/CLK _20595_/D vssd1 vssd1 vccd1 vccd1 _20595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1506 _11916_/S vssd1 vssd1 vccd1 vccd1 _11527_/S sky130_fd_sc_hd__buf_6
XFILLER_238_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1517 _12139_/S vssd1 vssd1 vccd1 vccd1 _12146_/S sky130_fd_sc_hd__buf_6
XFILLER_132_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout530 _17574_/X vssd1 vssd1 vccd1 vccd1 _17590_/S sky130_fd_sc_hd__buf_12
Xfanout1528 _10428_/S vssd1 vssd1 vccd1 vccd1 _10426_/S sky130_fd_sc_hd__buf_6
Xfanout1539 _10137_/C vssd1 vssd1 vccd1 vccd1 _10217_/S sky130_fd_sc_hd__buf_6
Xfanout541 _17166_/S vssd1 vssd1 vccd1 vccd1 _17183_/S sky130_fd_sc_hd__buf_12
X_09909_ _11851_/A _19323_/Q _11851_/C vssd1 vssd1 vccd1 vccd1 _09909_/X sky130_fd_sc_hd__or3_1
Xfanout552 _17076_/S vssd1 vssd1 vccd1 vccd1 _17078_/S sky130_fd_sc_hd__clkbuf_16
Xfanout563 _16639_/X vssd1 vssd1 vccd1 vccd1 _16670_/S sky130_fd_sc_hd__buf_6
Xfanout574 _16471_/S vssd1 vssd1 vccd1 vccd1 _16488_/S sky130_fd_sc_hd__buf_12
Xfanout585 _16106_/A2 vssd1 vssd1 vccd1 vccd1 _16126_/A2 sky130_fd_sc_hd__buf_4
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20029_ _20467_/CLK _20029_/D vssd1 vssd1 vccd1 vccd1 _20029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout596 _14670_/X vssd1 vssd1 vccd1 vccd1 _14699_/S sky130_fd_sc_hd__buf_12
X_12920_ _12918_/Y _12919_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _12920_/X sky130_fd_sc_hd__o21a_1
XFILLER_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9__f_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_9__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_62_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12851_ _12852_/A _12852_/B _12852_/C vssd1 vssd1 vccd1 vccd1 _12851_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11802_ _11761_/A _11761_/B _09859_/X vssd1 vssd1 vccd1 vccd1 _11802_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ input269/X _15013_/Y _15564_/X _15606_/A1 vssd1 vssd1 vccd1 vccd1 _15570_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12782_/A _12782_/B vssd1 vssd1 vccd1 vccd1 _12782_/X sky130_fd_sc_hd__or2_1
XFILLER_215_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _13612_/A _16133_/B _19299_/Q vssd1 vssd1 vccd1 vccd1 _14522_/B sky130_fd_sc_hd__a21oi_1
XFILLER_187_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11729_/A _11733_/B vssd1 vssd1 vccd1 vccd1 _11733_/Y sky130_fd_sc_hd__nand2b_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _20185_/Q _17235_/Y _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17240_/X sky130_fd_sc_hd__a21o_1
XFILLER_186_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _18694_/A _14452_/B vssd1 vssd1 vccd1 vccd1 _19250_/D sky130_fd_sc_hd__and2_1
XFILLER_186_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _19680_/Q _20168_/Q _11665_/S vssd1 vssd1 vccd1 vccd1 _11664_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13403_ _19230_/Q _13403_/B vssd1 vssd1 vccd1 vccd1 _13403_/X sky130_fd_sc_hd__xor2_1
XFILLER_186_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17171_ _20137_/Q _17696_/A1 _17178_/S vssd1 vssd1 vccd1 vccd1 _20137_/D sky130_fd_sc_hd__mux2_1
X_10615_ _19375_/Q _10603_/B _10613_/X _11718_/S _10614_/X vssd1 vssd1 vccd1 vccd1
+ _10615_/X sky130_fd_sc_hd__o221a_1
X_14383_ _19520_/Q _14383_/B vssd1 vssd1 vccd1 vccd1 _14384_/B sky130_fd_sc_hd__nand2_1
XFILLER_259_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11595_ _12138_/A1 _20512_/Q _11980_/S _11585_/X vssd1 vssd1 vccd1 vccd1 _11595_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_259_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16122_ _10468_/X _16132_/A2 _16121_/X vssd1 vssd1 vccd1 vccd1 _19585_/D sky130_fd_sc_hd__o21a_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13334_ _13334_/A _13334_/B _13334_/C vssd1 vssd1 vccd1 vccd1 _13334_/X sky130_fd_sc_hd__or3_1
X_10546_ _11239_/A1 _13978_/A2 _10545_/X _11239_/B1 _19840_/Q vssd1 vssd1 vccd1 vccd1
+ _10546_/X sky130_fd_sc_hd__o32a_1
XFILLER_109_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16053_ _16053_/A _16053_/B vssd1 vssd1 vccd1 vccd1 _16053_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _13264_/B _13264_/C _13264_/A vssd1 vssd1 vccd1 vccd1 _13265_/Y sky130_fd_sc_hd__a21oi_1
X_10477_ _19672_/Q _20160_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _10477_/X sky130_fd_sc_hd__mux2_1
X_15004_ _20786_/Q _14987_/Y _14989_/X _15003_/X vssd1 vssd1 vccd1 vccd1 _15004_/X
+ sky130_fd_sc_hd__a211o_1
X_12216_ _09503_/A _12371_/A1 _19363_/Q _12377_/S vssd1 vssd1 vccd1 vccd1 _12216_/X
+ sky130_fd_sc_hd__a31o_1
X_13196_ _13195_/A _13195_/B _13195_/Y _13397_/B vssd1 vssd1 vccd1 vccd1 _13196_/X
+ sky130_fd_sc_hd__a211o_1
X_19812_ _20539_/CLK _19812_/D vssd1 vssd1 vccd1 vccd1 _19812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12147_ _12134_/S _12146_/X _12145_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _12147_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_2_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19743_ _20763_/CLK _19743_/D vssd1 vssd1 vccd1 vccd1 _19743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16955_ _20422_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16955_/X sky130_fd_sc_hd__a21o_1
X_12078_ _12084_/A _19923_/Q _12081_/S0 _20048_/Q vssd1 vssd1 vccd1 vccd1 _12078_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_249_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11029_ _11027_/X _11028_/X _11033_/S vssd1 vssd1 vccd1 vccd1 _11029_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15906_ _19728_/Q _15933_/B vssd1 vssd1 vccd1 vccd1 _15906_/X sky130_fd_sc_hd__or2_1
X_16886_ _16932_/B1 _16882_/X _16885_/Y _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16887_/B
+ sky130_fd_sc_hd__o2bb2a_4
X_19674_ _20711_/CLK _19674_/D vssd1 vssd1 vccd1 vccd1 _19674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_265_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15837_ _16024_/A1 _15835_/X _15836_/Y _15816_/A _15975_/B2 vssd1 vssd1 vccd1 vccd1
+ _15837_/X sky130_fd_sc_hd__a32o_1
X_18625_ _18511_/X _18688_/A2 _18623_/Y _18624_/Y vssd1 vssd1 vccd1 vccd1 _18626_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18556_ _18651_/B _18556_/B vssd1 vssd1 vccd1 vccd1 _18556_/X sky130_fd_sc_hd__or2_2
X_15768_ _15768_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15768_/X sky130_fd_sc_hd__and2_1
XFILLER_52_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14719_ _19476_/Q _17657_/A1 _14719_/S vssd1 vssd1 vccd1 vccd1 _19476_/D sky130_fd_sc_hd__mux2_1
X_17507_ _17525_/A1 _17506_/Y _18932_/A vssd1 vssd1 vccd1 vccd1 _20288_/D sky130_fd_sc_hd__a21oi_1
X_18487_ _18604_/B _18487_/B vssd1 vssd1 vccd1 vccd1 _18487_/X sky130_fd_sc_hd__or2_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15699_ _16050_/A1 _15698_/X _15686_/Y vssd1 vssd1 vccd1 vccd1 _15699_/X sky130_fd_sc_hd__a21o_1
XFILLER_268_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_490 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17438_ _17452_/A _17438_/B vssd1 vssd1 vccd1 vccd1 _17438_/X sky130_fd_sc_hd__or2_1
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 _15480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_26 _15689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_37 _16728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_48 _16887_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ _20233_/Q _17371_/A2 _17368_/X _18720_/A vssd1 vssd1 vccd1 vccd1 _20233_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_59 _17336_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19108_ _20273_/CLK _19108_/D vssd1 vssd1 vccd1 vccd1 _19108_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20380_ _20702_/CLK _20380_/D vssd1 vssd1 vccd1 vccd1 _20380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19039_ _21038_/Q _19049_/A2 _19038_/X _18746_/A vssd1 vssd1 vccd1 vccd1 _21038_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21001_ _21010_/CLK _21001_/D vssd1 vssd1 vccd1 vccd1 _21001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_68_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20659_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09625_ _11345_/S _10979_/C vssd1 vssd1 vccd1 vccd1 _09625_/Y sky130_fd_sc_hd__nand2_8
XFILLER_216_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09556_ _09556_/A _12574_/A vssd1 vssd1 vccd1 vccd1 _09556_/X sky130_fd_sc_hd__or2_2
XFILLER_270_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09487_ _11234_/A vssd1 vssd1 vccd1 vccd1 _18163_/B sky130_fd_sc_hd__inv_4
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20716_ _20716_/CLK _20716_/D vssd1 vssd1 vccd1 vccd1 _20716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20647_ _20647_/CLK _20647_/D vssd1 vssd1 vccd1 vccd1 _20647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10400_ _20129_/Q _20097_/Q _10400_/S vssd1 vssd1 vccd1 vccd1 _10400_/X sky130_fd_sc_hd__mux2_1
X_11380_ _20469_/Q _11377_/S _12419_/C1 vssd1 vssd1 vccd1 vccd1 _11380_/X sky130_fd_sc_hd__o21a_1
X_20578_ _20714_/CLK _20578_/D vssd1 vssd1 vccd1 vccd1 _20578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10331_ _14894_/A _15922_/B2 _10330_/X vssd1 vssd1 vccd1 vccd1 _10365_/A sky130_fd_sc_hd__a21oi_4
XFILLER_124_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10262_ _10262_/A _19317_/Q _11021_/C vssd1 vssd1 vccd1 vccd1 _10262_/X sky130_fd_sc_hd__or3_1
XFILLER_180_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ _20953_/Q _20887_/Q vssd1 vssd1 vccd1 vccd1 _13050_/X sky130_fd_sc_hd__or2_1
XFILLER_152_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout2004 _16866_/B2 vssd1 vssd1 vccd1 vccd1 _16740_/B2 sky130_fd_sc_hd__buf_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _12519_/A _11649_/S _12000_/Y vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__o21a_1
XFILLER_87_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10193_ _10181_/X _10192_/X _12275_/A vssd1 vssd1 vccd1 vccd1 _10193_/X sky130_fd_sc_hd__mux2_2
XFILLER_278_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1303 _13468_/B vssd1 vssd1 vccd1 vccd1 _16982_/B1 sky130_fd_sc_hd__buf_6
XFILLER_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1314 _14822_/S vssd1 vssd1 vccd1 vccd1 _14870_/S sky130_fd_sc_hd__buf_6
XFILLER_79_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1325 _12462_/Y vssd1 vssd1 vccd1 vccd1 _12463_/B sky130_fd_sc_hd__buf_4
XFILLER_120_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1336 _11392_/A2 vssd1 vssd1 vccd1 vccd1 _12255_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_266_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1347 _17356_/A2 vssd1 vssd1 vccd1 vccd1 _17321_/A2 sky130_fd_sc_hd__buf_6
XFILLER_238_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1358 _16525_/X vssd1 vssd1 vccd1 vccd1 _16567_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_219_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1369 _14267_/A2 vssd1 vssd1 vccd1 vccd1 _14237_/A2 sky130_fd_sc_hd__buf_8
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16740_ _16982_/B1 _16737_/X _16739_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16741_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_13952_ _19183_/Q _14047_/C _14003_/S vssd1 vssd1 vccd1 vccd1 _13952_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _15960_/A _12486_/B _12484_/X _12902_/Y vssd1 vssd1 vccd1 vccd1 _12903_/X
+ sky130_fd_sc_hd__o22a_1
X_16671_ _19928_/Q _17674_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19928_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13883_ _19101_/Q _14738_/B _13889_/B1 _15678_/A1 _16189_/A vssd1 vssd1 vccd1 vccd1
+ _19101_/D sky130_fd_sc_hd__o221a_1
XFILLER_262_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18410_ _18414_/A _18410_/B vssd1 vssd1 vccd1 vccd1 _20859_/D sky130_fd_sc_hd__and2_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15622_ _19165_/Q _16063_/A2 _16036_/A2 vssd1 vssd1 vccd1 vccd1 _15622_/X sky130_fd_sc_hd__a21bo_1
X_19390_ _20678_/CLK _19390_/D vssd1 vssd1 vccd1 vccd1 _19390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _19512_/Q _12845_/A vssd1 vssd1 vccd1 vccd1 _12835_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18341_ _18490_/B _18341_/B vssd1 vssd1 vccd1 vccd1 _18341_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _16053_/A _15547_/X _15550_/Y _15365_/A vssd1 vssd1 vccd1 vccd1 _15553_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12763_/X _12764_/Y _12752_/B vssd1 vssd1 vccd1 vccd1 _12767_/A sky130_fd_sc_hd__a21oi_4
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14504_ _19282_/Q _17099_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19282_/D sky130_fd_sc_hd__mux2_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _18724_/A _18272_/B vssd1 vssd1 vccd1 vccd1 _20808_/D sky130_fd_sc_hd__and2_1
X_11716_ _09834_/A _20040_/Q _19915_/Q _10621_/S vssd1 vssd1 vccd1 vccd1 _11716_/X
+ sky130_fd_sc_hd__a22o_1
X_15484_ _19745_/Q _15604_/A2 _15483_/X _16048_/C1 vssd1 vssd1 vccd1 vccd1 _15484_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12696_ _12698_/A _12698_/B vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17223_ _14130_/B _17219_/Y _17222_/X _18698_/A vssd1 vssd1 vccd1 vccd1 _20183_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14435_ _14435_/A _14435_/B vssd1 vssd1 vccd1 vccd1 _14435_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_174_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ _12194_/A1 _17905_/A1 _11646_/Y _09750_/Y vssd1 vssd1 vccd1 vccd1 _15713_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_238_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 core_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_4
XFILLER_156_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17154_ _20120_/Q _17922_/A1 _17166_/S vssd1 vssd1 vccd1 vccd1 _20120_/D sky130_fd_sc_hd__mux2_1
Xinput24 core_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_4
XFILLER_167_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14366_ _14366_/A _14366_/B vssd1 vssd1 vccd1 vccd1 _14367_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput35 core_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_4
X_11578_ _19884_/Q _19785_/Q _11978_/S vssd1 vssd1 vccd1 vccd1 _11578_/X sky130_fd_sc_hd__mux2_1
Xinput46 dout0[12] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput57 dout0[22] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_2
X_16105_ _19577_/Q _16067_/X _16143_/A vssd1 vssd1 vccd1 vccd1 _16105_/X sky130_fd_sc_hd__o21a_1
Xinput68 dout0[32] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13317_ _13316_/A _13316_/B _13607_/B vssd1 vssd1 vccd1 vccd1 _13317_/Y sky130_fd_sc_hd__a21oi_2
X_17085_ _20055_/Q _17678_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20055_/D sky130_fd_sc_hd__mux2_1
X_10529_ _19633_/Q _19939_/Q _19277_/Q _20064_/Q _11292_/S0 _11026_/C vssd1 vssd1
+ vccd1 vccd1 _10529_/X sky130_fd_sc_hd__mux4_1
Xinput79 dout0[42] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14297_ _19232_/Q _14398_/A2 _14295_/X _14296_/X _14776_/C1 vssd1 vssd1 vccd1 vccd1
+ _19232_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16036_ _19557_/Q _16036_/A2 _16034_/X _16035_/X _16171_/A vssd1 vssd1 vccd1 vccd1
+ _19557_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13248_ _13248_/A _13321_/C vssd1 vssd1 vccd1 vccd1 _13362_/C sky130_fd_sc_hd__or2_2
XFILLER_269_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13179_ _12438_/Y _13178_/B _16026_/S vssd1 vssd1 vccd1 vccd1 _13180_/B sky130_fd_sc_hd__o21bai_4
XFILLER_285_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17987_ _20733_/Q _17984_/A _17986_/Y vssd1 vssd1 vccd1 vccd1 _20733_/D sky130_fd_sc_hd__o21a_1
XFILLER_284_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19726_ _19759_/CLK _19726_/D vssd1 vssd1 vccd1 vccd1 _19726_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1870 _15649_/A1 vssd1 vssd1 vccd1 vccd1 _12103_/A1 sky130_fd_sc_hd__buf_6
X_16938_ _19238_/Q _16980_/A2 _16980_/B1 _19107_/Q _16937_/X vssd1 vssd1 vccd1 vccd1
+ _16938_/X sky130_fd_sc_hd__o221a_1
XFILLER_226_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1881 _12510_/C vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__buf_8
XFILLER_284_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1892 _13887_/C1 vssd1 vssd1 vccd1 vccd1 _16185_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_203_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19657_ _20410_/CLK _19657_/D vssd1 vssd1 vccd1 vccd1 _19657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ _16869_/A _16869_/B vssd1 vssd1 vccd1 vccd1 _16869_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18608_ _19505_/Q _18612_/B vssd1 vssd1 vccd1 vccd1 _18608_/Y sky130_fd_sc_hd__nand2_1
XFILLER_252_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19588_ _19590_/CLK _19588_/D vssd1 vssd1 vccd1 vccd1 _19588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18539_ _20906_/Q fanout750/X _18538_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18540_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xclkbuf_leaf_186_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20263_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_279_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_115_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20863_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20501_ _20633_/CLK _20501_/D vssd1 vssd1 vccd1 vccd1 _20501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_194_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20432_ _20565_/CLK _20432_/D vssd1 vssd1 vccd1 vccd1 _20432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20363_ _20630_/CLK _20363_/D vssd1 vssd1 vccd1 vccd1 _20363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20294_ _20296_/CLK _20294_/D vssd1 vssd1 vccd1 vccd1 _20294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _19090_/Q _19089_/Q _19088_/Q _09610_/A vssd1 vssd1 vccd1 vccd1 _12976_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_113_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10880_ _10870_/X _10879_/Y _11201_/A _10862_/X vssd1 vssd1 vccd1 vccd1 _10880_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _19153_/Q _12480_/B vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__and2_2
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ _12550_/A _12550_/B _12550_/C _12550_/D vssd1 vssd1 vccd1 vccd1 _12555_/A
+ sky130_fd_sc_hd__or4_4
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11501_ _19414_/Q _11916_/S vssd1 vssd1 vccd1 vccd1 _11501_/X sky130_fd_sc_hd__or2_1
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12481_ _12579_/D _15220_/B vssd1 vssd1 vccd1 vccd1 _12493_/A sky130_fd_sc_hd__and2_4
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14220_ _14209_/A _14211_/B _14209_/B vssd1 vssd1 vccd1 vccd1 _14221_/B sky130_fd_sc_hd__a21bo_1
XFILLER_138_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11432_ _11423_/X _11425_/X _11431_/X _12058_/S _12137_/A1 vssd1 vssd1 vccd1 vccd1
+ _11432_/X sky130_fd_sc_hd__o221a_1
XFILLER_22_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14151_ _14151_/A _14160_/B vssd1 vssd1 vccd1 vccd1 _14151_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11363_ _11363_/A1 _11359_/X _11362_/X _12399_/C1 vssd1 vssd1 vccd1 vccd1 _11363_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _20976_/Q _13397_/B vssd1 vssd1 vccd1 vccd1 _13102_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10314_ _20639_/Q _20603_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14082_ _19200_/Q _14082_/A2 _14081_/X _16087_/B1 vssd1 vssd1 vccd1 vccd1 _19200_/D
+ sky130_fd_sc_hd__o211a_1
X_11294_ _11288_/X _11293_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _11294_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17910_ _20681_/Q _17910_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20681_/D sky130_fd_sc_hd__mux2_1
X_13033_ _20961_/Q _20895_/Q vssd1 vssd1 vccd1 vccd1 _13033_/X sky130_fd_sc_hd__or2_4
X_10245_ _19413_/Q _20572_/Q _11042_/B vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__mux2_1
X_18890_ _18520_/X _18978_/B _18888_/X _18889_/Y vssd1 vssd1 vccd1 vccd1 _18891_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_133_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1100 _17946_/A1 vssd1 vssd1 vccd1 vccd1 _17806_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_239_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1111 _11886_/X vssd1 vssd1 vccd1 vccd1 _17877_/A1 sky130_fd_sc_hd__buf_6
XFILLER_121_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10176_ _20314_/Q _11305_/B vssd1 vssd1 vccd1 vccd1 _10176_/X sky130_fd_sc_hd__or2_1
X_17841_ _20616_/Q _17913_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20616_/D sky130_fd_sc_hd__mux2_1
Xfanout1122 _17905_/A1 vssd1 vssd1 vccd1 vccd1 _17871_/A1 sky130_fd_sc_hd__buf_4
Xfanout1133 _17927_/A1 vssd1 vssd1 vccd1 vccd1 _17859_/A1 sky130_fd_sc_hd__buf_4
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1144 _09870_/X vssd1 vssd1 vccd1 vccd1 _09936_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1155 _12402_/A1 vssd1 vssd1 vccd1 vccd1 _12245_/A1 sky130_fd_sc_hd__buf_12
XFILLER_78_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1166 _14930_/X vssd1 vssd1 vccd1 vccd1 _15133_/B sky130_fd_sc_hd__buf_6
XFILLER_78_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14984_ _15314_/B _14987_/B vssd1 vssd1 vccd1 vccd1 _14988_/B sky130_fd_sc_hd__or2_2
Xfanout1177 _13350_/B vssd1 vssd1 vccd1 vccd1 _13363_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17772_ _20551_/Q _17878_/A1 _17772_/S vssd1 vssd1 vccd1 vccd1 _20551_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1188 _10561_/A vssd1 vssd1 vccd1 vccd1 _12156_/A1 sky130_fd_sc_hd__buf_6
Xfanout1199 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17279_/C1 sky130_fd_sc_hd__buf_4
XFILLER_266_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19511_ _19511_/CLK _19511_/D vssd1 vssd1 vccd1 vccd1 _19511_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_263_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16723_ _18198_/B _17219_/B _16717_/X vssd1 vssd1 vccd1 vccd1 _16723_/X sky130_fd_sc_hd__a21o_1
X_13935_ _19139_/Q _13941_/B _13946_/B1 _13411_/A vssd1 vssd1 vccd1 vccd1 _19139_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16654_ _19911_/Q _17934_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19911_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19442_ _20451_/CLK _19442_/D vssd1 vssd1 vccd1 vccd1 _19442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13866_ _19086_/Q _13953_/A2 _13900_/A2 _19152_/Q _16197_/A vssd1 vssd1 vccd1 vccd1
+ _19086_/D sky130_fd_sc_hd__o221a_1
X_15605_ _19717_/Q _15395_/S _15604_/X vssd1 vssd1 vccd1 vccd1 _15605_/X sky130_fd_sc_hd__o21a_1
XFILLER_223_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12817_ _12872_/B _12817_/B vssd1 vssd1 vccd1 vccd1 _12817_/X sky130_fd_sc_hd__or2_1
X_19373_ _20664_/CLK _19373_/D vssd1 vssd1 vccd1 vccd1 _19373_/Q sky130_fd_sc_hd__dfxtp_1
X_16585_ _16591_/A _16585_/B vssd1 vssd1 vccd1 vccd1 _19858_/D sky130_fd_sc_hd__or2_1
XFILLER_234_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13797_ _13826_/A1 _13660_/B _13826_/B1 input243/X vssd1 vssd1 vccd1 vccd1 _13797_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15536_ _20863_/Q _15535_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15536_/X sky130_fd_sc_hd__mux2_1
X_18324_ _18981_/C _18324_/B vssd1 vssd1 vccd1 vccd1 _18324_/Y sky130_fd_sc_hd__nor2_8
XFILLER_188_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12749_/C _12748_/B vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__and2b_1
XFILLER_176_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18255_ _18523_/B vssd1 vssd1 vccd1 vccd1 _18255_/Y sky130_fd_sc_hd__clkinv_2
X_15467_ _15223_/X _15466_/X _15612_/S vssd1 vssd1 vccd1 vccd1 _15468_/B sky130_fd_sc_hd__mux2_4
X_12679_ _19161_/Q _12479_/X _15348_/B2 _10308_/S vssd1 vssd1 vccd1 vccd1 _12686_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17206_ _20170_/Q _17800_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20170_/D sky130_fd_sc_hd__mux2_1
X_14418_ _13139_/A _14417_/X _13138_/X vssd1 vssd1 vccd1 vccd1 _14419_/C sky130_fd_sc_hd__a21o_1
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18186_ _20791_/Q _18185_/Y _18311_/S vssd1 vssd1 vccd1 vccd1 _18187_/B sky130_fd_sc_hd__mux2_1
X_15398_ _15283_/A _15380_/Y _15457_/B1 vssd1 vssd1 vccd1 vccd1 _15398_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17137_ _20105_/Q _17696_/A1 _17144_/S vssd1 vssd1 vccd1 vccd1 _20105_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14349_ _19237_/Q _14438_/A2 _14348_/X _16191_/A vssd1 vssd1 vccd1 vccd1 _19237_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17068_ _20040_/Q _17870_/A1 _17076_/S vssd1 vssd1 vccd1 vccd1 _20040_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16019_ _20816_/Q _15016_/Y _15384_/Y _16018_/X vssd1 vssd1 vccd1 vccd1 _16019_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _12138_/A1 _20514_/Q _12143_/S _09872_/X vssd1 vssd1 vccd1 vccd1 _09890_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_258_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19709_ _20757_/CLK _19709_/D vssd1 vssd1 vccd1 vccd1 _19709_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_214_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20981_ _21013_/CLK _20981_/D vssd1 vssd1 vccd1 vccd1 _20981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_272_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_253_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20415_ _20666_/CLK _20415_/D vssd1 vssd1 vccd1 vccd1 _20415_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_147_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_83_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _19621_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20346_ _20638_/CLK _20346_/D vssd1 vssd1 vccd1 vccd1 _20346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20451_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20277_ _21016_/CLK _20277_/D vssd1 vssd1 vccd1 vccd1 _20277_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ _11234_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10553_/C sky130_fd_sc_hd__or2_1
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput203 localMemory_wb_adr_i[21] vssd1 vssd1 vccd1 vccd1 _12928_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput214 localMemory_wb_cyc_i vssd1 vssd1 vccd1 vccd1 _17014_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput225 localMemory_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_hd__buf_12
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput236 localMemory_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_hd__buf_12
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput247 localMemory_wb_sel_i[0] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput258 manufacturerID[4] vssd1 vssd1 vccd1 vccd1 _17251_/A sky130_fd_sc_hd__buf_2
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput269 partID[14] vssd1 vssd1 vccd1 vccd1 input269/X sky130_fd_sc_hd__clkbuf_2
XFILLER_236_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ _11975_/X _11977_/X _11980_/X _12135_/A _11981_/C1 vssd1 vssd1 vccd1 vccd1
+ _11981_/X sky130_fd_sc_hd__o221a_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13720_ _13663_/A _13757_/B _13719_/X vssd1 vssd1 vccd1 vccd1 _13721_/B sky130_fd_sc_hd__a21oi_4
X_10932_ _12513_/C _11281_/B vssd1 vssd1 vccd1 vccd1 _10932_/Y sky130_fd_sc_hd__nand2_2
XFILLER_204_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13651_ _13685_/A _13685_/B vssd1 vssd1 vccd1 vccd1 _13651_/Y sky130_fd_sc_hd__nand2_1
X_10863_ _20370_/Q _20434_/Q _12352_/S vssd1 vssd1 vccd1 vccd1 _10863_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _19505_/Q _19504_/Q _12782_/A vssd1 vssd1 vccd1 vccd1 _12754_/A sky130_fd_sc_hd__and3_1
X_16370_ _19734_/Q _19733_/Q _16370_/C vssd1 vssd1 vccd1 vccd1 _16372_/B sky130_fd_sc_hd__and3_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A _19223_/Q vssd1 vssd1 vccd1 vccd1 _13582_/Y sky130_fd_sc_hd__nand2_1
X_10794_ _12275_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10794_/Y sky130_fd_sc_hd__nor2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15396_/A1 _15305_/X _15320_/X vssd1 vssd1 vccd1 vccd1 _16784_/B sky130_fd_sc_hd__a21oi_4
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12533_ _12533_/A _12533_/B vssd1 vssd1 vccd1 vccd1 _12587_/A sky130_fd_sc_hd__or2_2
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18040_ _18126_/A _18045_/C vssd1 vssd1 vccd1 vccd1 _18040_/Y sky130_fd_sc_hd__nor2_1
X_15252_ _15060_/X _15045_/X _15292_/S vssd1 vssd1 vccd1 vccd1 _15545_/B sky130_fd_sc_hd__mux2_1
X_12464_ _12464_/A _12468_/B _12464_/C vssd1 vssd1 vccd1 vccd1 _15026_/A sky130_fd_sc_hd__and3_4
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14203_ _13582_/A _14202_/X _13581_/Y vssd1 vssd1 vccd1 vccd1 _14204_/C sky130_fd_sc_hd__a21bo_1
X_11415_ _11415_/A _11415_/B vssd1 vssd1 vccd1 vccd1 _11415_/X sky130_fd_sc_hd__or2_1
X_15183_ _12463_/B _15177_/X _15182_/Y _14882_/B vssd1 vssd1 vccd1 vccd1 _15184_/B
+ sky130_fd_sc_hd__o22a_1
X_12395_ _12393_/X _12394_/X _12395_/S vssd1 vssd1 vccd1 vccd1 _12395_/X sky130_fd_sc_hd__mux2_1
X_14134_ _14255_/A _14204_/B _14134_/C vssd1 vssd1 vccd1 vccd1 _14134_/X sky130_fd_sc_hd__or3_1
X_11346_ _11345_/S _11334_/X _11338_/X _12310_/C1 vssd1 vssd1 vccd1 vccd1 _11346_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19991_ _19992_/CLK _19991_/D vssd1 vssd1 vccd1 vccd1 _19991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ _14081_/A _16133_/B _14065_/C vssd1 vssd1 vccd1 vccd1 _14065_/X sky130_fd_sc_hd__or3_1
X_18942_ _19143_/Q _18976_/A2 _18949_/B1 vssd1 vssd1 vccd1 vccd1 _18942_/Y sky130_fd_sc_hd__a21oi_1
X_11277_ _09689_/A _11260_/X _11276_/X _11012_/A vssd1 vssd1 vccd1 vccd1 _11277_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13016_ _20971_/Q _20905_/Q vssd1 vssd1 vccd1 vccd1 _13016_/Y sky130_fd_sc_hd__nand2_2
XFILLER_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10228_ _11250_/S _10227_/X _10226_/X _11009_/B2 vssd1 vssd1 vccd1 vccd1 _10228_/X
+ sky130_fd_sc_hd__a211o_1
X_18873_ _19133_/Q _12533_/B _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18873_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17824_ _20599_/Q _17896_/A1 _17845_/S vssd1 vssd1 vccd1 vccd1 _20599_/D sky130_fd_sc_hd__mux2_1
XFILLER_255_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10159_ _12301_/S _10158_/X _10157_/X _11353_/C1 vssd1 vssd1 vccd1 vccd1 _10159_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_121_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14967_ _14967_/A _15014_/D vssd1 vssd1 vccd1 vccd1 _14987_/A sky130_fd_sc_hd__nand2_2
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17755_ _20534_/Q _17861_/A1 _17772_/S vssd1 vssd1 vccd1 vccd1 _20534_/D sky130_fd_sc_hd__mux2_1
XFILLER_270_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16706_ _12962_/S _12930_/B _16279_/B _13473_/B _13472_/Y vssd1 vssd1 vccd1 vccd1
+ _16706_/X sky130_fd_sc_hd__a221o_4
X_13918_ _18710_/A _13918_/B vssd1 vssd1 vccd1 vccd1 _19124_/D sky130_fd_sc_hd__and2_1
X_14898_ _14898_/A _15096_/A vssd1 vssd1 vccd1 vccd1 _14898_/Y sky130_fd_sc_hd__nand2_1
X_17686_ _20470_/Q _17686_/A1 _17703_/S vssd1 vssd1 vccd1 vccd1 _20470_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19425_ _20716_/CLK _19425_/D vssd1 vssd1 vccd1 vccd1 _19425_/Q sky130_fd_sc_hd__dfxtp_1
X_16637_ _19896_/Q _17674_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19896_/D sky130_fd_sc_hd__mux2_1
X_13849_ _20265_/Q _20264_/Q vssd1 vssd1 vccd1 vccd1 _17451_/B sky130_fd_sc_hd__nand2b_2
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19356_ _20711_/CLK _19356_/D vssd1 vssd1 vccd1 vccd1 _19356_/Q sky130_fd_sc_hd__dfxtp_1
X_16568_ _19850_/Q _16576_/A2 _16576_/B1 input20/X vssd1 vssd1 vccd1 vccd1 _16569_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_222_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18307_ _18718_/A _18307_/B vssd1 vssd1 vccd1 vccd1 _20815_/D sky130_fd_sc_hd__and2_1
X_15519_ _16052_/A1 _15505_/X _15518_/Y _15494_/A _15442_/A vssd1 vssd1 vccd1 vccd1
+ _15519_/X sky130_fd_sc_hd__a32o_1
X_16499_ _19806_/Q _17058_/A1 _16521_/S vssd1 vssd1 vccd1 vccd1 _19806_/D sky130_fd_sc_hd__mux2_1
X_19287_ _20717_/CLK _19287_/D vssd1 vssd1 vccd1 vccd1 _19287_/Q sky130_fd_sc_hd__dfxtp_1
X_18238_ _19543_/Q _18248_/B vssd1 vssd1 vccd1 vccd1 _18238_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18169_ _18213_/B _14139_/B _18168_/Y vssd1 vssd1 vccd1 vccd1 _18466_/B sky130_fd_sc_hd__o21ai_4
XFILLER_172_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20200_ _20727_/CLK _20200_/D vssd1 vssd1 vccd1 vccd1 _20200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20131_ _20718_/CLK _20131_/D vssd1 vssd1 vccd1 vccd1 _20131_/Q sky130_fd_sc_hd__dfxtp_1
X_09942_ _19547_/Q _12155_/A2 _12155_/B1 _19611_/Q vssd1 vssd1 vccd1 vccd1 _09942_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout904 _15322_/C vssd1 vssd1 vccd1 vccd1 _15939_/A2 sky130_fd_sc_hd__buf_6
Xfanout915 _16011_/B1 vssd1 vssd1 vccd1 vccd1 _16041_/B1 sky130_fd_sc_hd__buf_8
Xfanout926 _14935_/Y vssd1 vssd1 vccd1 vccd1 _15595_/B1 sky130_fd_sc_hd__buf_4
X_20062_ _20181_/CLK _20062_/D vssd1 vssd1 vccd1 vccd1 _20062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout937 _11223_/A vssd1 vssd1 vccd1 vccd1 _15155_/S sky130_fd_sc_hd__buf_4
X_09873_ _19950_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _09873_/X sky130_fd_sc_hd__or2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout948 _15118_/S vssd1 vssd1 vccd1 vccd1 _15612_/S sky130_fd_sc_hd__buf_6
XFILLER_85_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout959 _11397_/A2 vssd1 vssd1 vccd1 vccd1 _17894_/A1 sky130_fd_sc_hd__clkbuf_4
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_261_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_308 input235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_130_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21021_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_319 _13614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20964_ _20998_/CLK _20964_/D vssd1 vssd1 vccd1 vccd1 _20964_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20895_ _21025_/CLK _20895_/D vssd1 vssd1 vccd1 vccd1 _20895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11200_ _11194_/X _11199_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12180_ _19651_/Q _19957_/Q _12182_/S vssd1 vssd1 vccd1 vccd1 _12181_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11131_ _11396_/S _11131_/B vssd1 vssd1 vccd1 vccd1 _11131_/Y sky130_fd_sc_hd__nor2_1
XFILLER_268_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20329_ _20641_/CLK _20329_/D vssd1 vssd1 vccd1 vccd1 _20329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ _19561_/Q _11061_/A _09659_/X _11061_/Y vssd1 vssd1 vccd1 vccd1 _11062_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10013_ _12194_/A1 _17906_/A1 _10012_/X _12194_/B2 vssd1 vssd1 vccd1 vccd1 _15741_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ _15870_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15870_/X sky130_fd_sc_hd__and2_1
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_218_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _21046_/A
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ _11742_/B _10640_/B _14822_/S vssd1 vssd1 vccd1 vccd1 _14821_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_251_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _17745_/A _17676_/B _17540_/C vssd1 vssd1 vccd1 vccd1 _17540_/X sky130_fd_sc_hd__and3_4
X_14752_ _19123_/Q _14764_/A2 _14751_/X _18476_/A vssd1 vssd1 vccd1 vccd1 _19500_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _12156_/A1 _11963_/X _11962_/X vssd1 vssd1 vccd1 vccd1 _11964_/X sky130_fd_sc_hd__a21o_1
XFILLER_251_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13742_/A _13730_/B vssd1 vssd1 vccd1 vccd1 _13703_/Y sky130_fd_sc_hd__nor2_1
X_10915_ _20154_/Q _12213_/B vssd1 vssd1 vccd1 vccd1 _10915_/X sky130_fd_sc_hd__or2_1
X_17471_ _17495_/A1 _17470_/Y _18704_/A vssd1 vssd1 vccd1 vccd1 _20270_/D sky130_fd_sc_hd__a21oi_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14683_ _19442_/Q _17689_/A1 _14699_/S vssd1 vssd1 vccd1 vccd1 _19442_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11895_ _20358_/Q _11895_/B vssd1 vssd1 vccd1 vccd1 _11895_/X sky130_fd_sc_hd__or2_1
X_19210_ _19704_/CLK _19210_/D vssd1 vssd1 vccd1 vccd1 _19210_/Q sky130_fd_sc_hd__dfxtp_1
X_13634_ _15954_/A _13189_/B _16235_/B _13478_/B vssd1 vssd1 vccd1 vccd1 _13634_/X
+ sky130_fd_sc_hd__a31o_2
X_16422_ _19753_/Q _16420_/B _16421_/Y vssd1 vssd1 vccd1 vccd1 _19753_/D sky130_fd_sc_hd__o21a_1
X_10846_ _12392_/C1 _10835_/X _10838_/X _10845_/X _12400_/A1 vssd1 vssd1 vccd1 vccd1
+ _10846_/X sky130_fd_sc_hd__a311o_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19141_ _20291_/CLK _19141_/D vssd1 vssd1 vccd1 vccd1 _19141_/Q sky130_fd_sc_hd__dfxtp_1
X_16353_ _19727_/Q _16354_/C _19728_/Q vssd1 vssd1 vccd1 vccd1 _16355_/B sky130_fd_sc_hd__a21oi_1
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ _18589_/B _13563_/X _13564_/Y _13561_/Y _13582_/A vssd1 vssd1 vccd1 vccd1
+ _13565_/X sky130_fd_sc_hd__a311o_4
XFILLER_9_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10777_ _10771_/X _10776_/X _12415_/S vssd1 vssd1 vccd1 vccd1 _10777_/X sky130_fd_sc_hd__mux2_2
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15304_ _15304_/A _16009_/B vssd1 vssd1 vccd1 vccd1 _15304_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12516_ _12516_/A _12588_/B _12516_/C vssd1 vssd1 vccd1 vccd1 _12516_/Y sky130_fd_sc_hd__nor3_4
X_19072_ _20417_/Q vssd1 vssd1 vccd1 vccd1 _20417_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_200_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16284_ _20006_/Q split1/X _19701_/D vssd1 vssd1 vccd1 vccd1 _19700_/D sky130_fd_sc_hd__and3_1
XFILLER_200_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13496_ _15185_/A vssd1 vssd1 vccd1 vccd1 _13496_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15235_ _20918_/Q _15567_/A2 _15234_/X vssd1 vssd1 vccd1 vccd1 _15235_/X sky130_fd_sc_hd__o21a_1
XFILLER_185_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18023_ _20746_/Q _18024_/C _18022_/Y vssd1 vssd1 vccd1 vccd1 _20746_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12447_ _12447_/A _12447_/B vssd1 vssd1 vccd1 vccd1 _16054_/A sky130_fd_sc_hd__nor2_4
XFILLER_246_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15166_ _15166_/A vssd1 vssd1 vccd1 vccd1 _15166_/Y sky130_fd_sc_hd__inv_2
X_12378_ _20555_/Q _12397_/S vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__or2_1
XFILLER_5_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14117_ _14117_/A _14117_/B _16716_/B vssd1 vssd1 vccd1 vccd1 _14117_/Y sky130_fd_sc_hd__nor3_4
X_11329_ _09638_/Y _11327_/Y _11328_/X _10035_/Y vssd1 vssd1 vccd1 vccd1 _11329_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_259_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19974_ _21016_/CLK _19974_/D vssd1 vssd1 vccd1 vccd1 _19974_/Q sky130_fd_sc_hd__dfxtp_1
X_15097_ _15283_/A _15078_/X _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__a21o_1
X_14048_ _19183_/Q _14082_/A2 _14047_/X _16087_/B1 vssd1 vssd1 vccd1 vccd1 _19183_/D
+ sky130_fd_sc_hd__o211a_1
X_18925_ _18932_/A _18925_/B vssd1 vssd1 vccd1 vccd1 _21003_/D sky130_fd_sc_hd__nor2_1
X_18856_ _18856_/A _18856_/B vssd1 vssd1 vccd1 vccd1 _20993_/D sky130_fd_sc_hd__nor2_1
XFILLER_121_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17807_ _20584_/Q _17947_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20584_/D sky130_fd_sc_hd__mux2_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18787_ _19497_/Q _18901_/S _18786_/X _18589_/B vssd1 vssd1 vccd1 vccd1 _18787_/X
+ sky130_fd_sc_hd__o211a_1
X_15999_ _19763_/Q _15999_/A2 _15998_/X _15999_/C1 vssd1 vssd1 vccd1 vccd1 _15999_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_282_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17738_ _20519_/Q _17878_/A1 _17738_/S vssd1 vssd1 vccd1 vccd1 _20519_/D sky130_fd_sc_hd__mux2_1
XFILLER_270_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17669_ _20455_/Q _17806_/A1 _17669_/S vssd1 vssd1 vccd1 vccd1 _20455_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_250_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19408_ _20701_/CLK _19408_/D vssd1 vssd1 vccd1 vccd1 _19408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20680_ _20706_/CLK _20680_/D vssd1 vssd1 vccd1 vccd1 _20680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19339_ _20694_/CLK _19339_/D vssd1 vssd1 vccd1 vccd1 _19339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout701 _13855_/Y vssd1 vssd1 vccd1 vccd1 _14081_/A sky130_fd_sc_hd__buf_6
XFILLER_160_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09925_ _09922_/X _09924_/X _11949_/S vssd1 vssd1 vccd1 vccd1 _09925_/Y sky130_fd_sc_hd__a21oi_1
X_20114_ _20641_/CLK _20114_/D vssd1 vssd1 vccd1 vccd1 _20114_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout712 _16279_/B vssd1 vssd1 vccd1 vccd1 split2/A sky130_fd_sc_hd__buf_12
XFILLER_277_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout723 _13480_/Y vssd1 vssd1 vccd1 vccd1 _13663_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_259_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout734 _18997_/B vssd1 vssd1 vccd1 vccd1 _19013_/B sky130_fd_sc_hd__buf_6
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout745 _18818_/A2 vssd1 vssd1 vccd1 vccd1 _18867_/A2 sky130_fd_sc_hd__buf_6
X_20045_ _20077_/CLK _20045_/D vssd1 vssd1 vccd1 vccd1 _20045_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout756 _18937_/B vssd1 vssd1 vccd1 vccd1 _18978_/B sky130_fd_sc_hd__buf_4
X_09856_ _12105_/A _09847_/X _09855_/X _09839_/X vssd1 vssd1 vccd1 vccd1 _09856_/X
+ sky130_fd_sc_hd__o31a_4
Xfanout767 _18593_/A2 vssd1 vssd1 vccd1 vccd1 _18462_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_219_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout778 _18616_/B vssd1 vssd1 vccd1 vccd1 _18604_/B sky130_fd_sc_hd__buf_4
XFILLER_218_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout789 _12786_/B vssd1 vssd1 vccd1 vccd1 _12758_/B sky130_fd_sc_hd__buf_6
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09787_ _09672_/A _14011_/A2 _09786_/X _11239_/B1 _19853_/Q vssd1 vssd1 vccd1 vccd1
+ _09787_/X sky130_fd_sc_hd__o32a_1
Xclkbuf_4_8__f_wb_clk_i clkbuf_3_4_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_8__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_105 _12963_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 _16235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_127 _13660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_138 _13711_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _21013_/CLK _20947_/D vssd1 vssd1 vccd1 vccd1 _20947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _13750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10700_ _12265_/A _10700_/B vssd1 vssd1 vccd1 vccd1 _10700_/Y sky130_fd_sc_hd__nor2_1
XFILLER_199_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _09806_/S _11679_/X _11678_/X _11680_/C1 vssd1 vssd1 vccd1 vccd1 _11680_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_186_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20878_ _21040_/CLK _20878_/D vssd1 vssd1 vccd1 vccd1 _20878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10631_ _10260_/S _10629_/X _10630_/X _12088_/S vssd1 vssd1 vccd1 vccd1 _10631_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_22_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13350_ _13350_/A _13350_/B _13350_/C _13349_/X vssd1 vssd1 vccd1 vccd1 _13352_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_128_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10562_ _19536_/Q _09596_/B _10543_/X _10561_/Y vssd1 vssd1 vccd1 vccd1 _10562_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12301_ _12299_/X _12300_/X _12301_/S vssd1 vssd1 vccd1 vccd1 _12301_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ _13281_/A _13281_/B vssd1 vssd1 vccd1 vccd1 _13281_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10493_ _11266_/A1 _20503_/Q _10316_/S _20535_/Q vssd1 vssd1 vccd1 vccd1 _10493_/X
+ sky130_fd_sc_hd__o22a_1
X_15020_ _15020_/A _15134_/B vssd1 vssd1 vccd1 vccd1 _15020_/Y sky130_fd_sc_hd__nor2_1
X_12232_ _12241_/S _12231_/X _12230_/X _12314_/C1 vssd1 vssd1 vccd1 vccd1 _12232_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _12161_/X _12162_/X _12189_/A vssd1 vssd1 vccd1 vccd1 _12163_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11114_ _11108_/X _11113_/X _12415_/S vssd1 vssd1 vccd1 vccd1 _11114_/X sky130_fd_sc_hd__mux2_2
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16971_ _20424_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16971_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12094_ _12103_/A1 _12092_/X _12093_/X vssd1 vssd1 vccd1 vccd1 _12095_/B sky130_fd_sc_hd__o21ai_1
XFILLER_122_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18710_ _18710_/A _18710_/B vssd1 vssd1 vccd1 vccd1 _20955_/D sky130_fd_sc_hd__and2_1
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11045_ _11042_/X _11043_/X _11044_/X _12429_/A1 _12430_/S vssd1 vssd1 vccd1 vccd1
+ _11045_/X sky130_fd_sc_hd__a221o_1
X_15922_ _12513_/A _16063_/A2 _15898_/A _15922_/B2 vssd1 vssd1 vccd1 vccd1 _15923_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19690_ _20641_/CLK _19690_/D vssd1 vssd1 vccd1 vccd1 _19690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18641_ _18523_/X _18688_/A2 _18639_/Y _18640_/Y vssd1 vssd1 vccd1 vccd1 _18642_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _20874_/Q _16018_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15853_/X sky130_fd_sc_hd__o21ba_1
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14804_ _19526_/Q _13609_/A _16167_/C1 _14803_/Y vssd1 vssd1 vccd1 vccd1 _19526_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_206_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18572_ _18783_/A _18572_/B vssd1 vssd1 vccd1 vccd1 _20915_/D sky130_fd_sc_hd__nor2_1
XFILLER_149_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _19241_/Q _19240_/Q _13231_/B vssd1 vssd1 vccd1 vccd1 _12996_/Y sky130_fd_sc_hd__nand3_1
X_15784_ _15526_/B _15767_/X _15783_/X _15976_/B2 vssd1 vssd1 vccd1 vccd1 _15784_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_92_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _17525_/A1 _17522_/Y _17430_/A vssd1 vssd1 vccd1 vccd1 _20296_/D sky130_fd_sc_hd__a21oi_1
X_14735_ _19492_/Q _17707_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19492_/D sky130_fd_sc_hd__mux2_1
XFILLER_217_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11947_ _19423_/Q _20582_/Q _11947_/S vssd1 vssd1 vccd1 vccd1 _11947_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_650 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _19428_/Q _17950_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19428_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17454_ _17454_/A _17454_/B _17454_/C _17454_/D vssd1 vssd1 vccd1 vccd1 _17454_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11878_ _11878_/A _11878_/B vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__nor2_4
XFILLER_205_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16405_ _18086_/A _16410_/C vssd1 vssd1 vccd1 vccd1 _16405_/Y sky130_fd_sc_hd__nor2_1
X_13617_ _13626_/A1 _13388_/D _13426_/B _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13617_/X
+ sky130_fd_sc_hd__a22o_2
X_10829_ _10814_/X _10815_/X _12309_/S vssd1 vssd1 vccd1 vccd1 _10829_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14597_ _19363_/Q _17949_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19363_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17385_ _20241_/Q _17401_/A2 _17384_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _20241_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19124_ _19698_/CLK _19124_/D vssd1 vssd1 vccd1 vccd1 _19124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13548_ _12652_/B _13543_/X _13544_/Y _13547_/X vssd1 vssd1 vccd1 vccd1 _13552_/B
+ sky130_fd_sc_hd__a31o_1
X_16336_ _19721_/Q _16338_/C _16335_/Y vssd1 vssd1 vccd1 vccd1 _19721_/D sky130_fd_sc_hd__o21a_1
XFILLER_158_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19055_ _20400_/Q vssd1 vssd1 vccd1 vccd1 _20400_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16267_ _19683_/Q _17801_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19683_/D sky130_fd_sc_hd__mux2_1
X_13479_ _13479_/A _13481_/A vssd1 vssd1 vccd1 vccd1 _13479_/X sky130_fd_sc_hd__and2_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18006_ _18094_/A _18011_/C vssd1 vssd1 vccd1 vccd1 _18006_/Y sky130_fd_sc_hd__nor2_1
X_15218_ _15258_/A _15218_/B vssd1 vssd1 vccd1 vccd1 _15218_/X sky130_fd_sc_hd__or2_1
X_16198_ _17850_/A _16672_/A vssd1 vssd1 vccd1 vccd1 _16199_/C sky130_fd_sc_hd__nor2_1
Xoutput304 _21047_/X vssd1 vssd1 vccd1 vccd1 clk1 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput315 _13622_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[19] sky130_fd_sc_hd__buf_4
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput326 _13510_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[3] sky130_fd_sc_hd__buf_4
XFILLER_160_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput337 _13687_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[12] sky130_fd_sc_hd__buf_4
XFILLER_113_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15149_ _15283_/A _15129_/X _15457_/B1 vssd1 vssd1 vccd1 vccd1 _15149_/X sky130_fd_sc_hd__a21o_1
XFILLER_5_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput348 _13733_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[22] sky130_fd_sc_hd__buf_4
Xoutput359 _13649_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[3] sky130_fd_sc_hd__buf_4
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19957_ _20075_/CLK _19957_/D vssd1 vssd1 vccd1 vccd1 _19957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09710_ _11983_/A1 _20516_/Q _11513_/S _09691_/X vssd1 vssd1 vccd1 vccd1 _09710_/X
+ sky130_fd_sc_hd__o211a_1
X_18908_ _19138_/Q _18976_/A2 _18767_/B vssd1 vssd1 vccd1 vccd1 _18908_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19888_ _20712_/CLK _19888_/D vssd1 vssd1 vccd1 vccd1 _19888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09641_ _09612_/X _09636_/B _09640_/Y vssd1 vssd1 vccd1 vccd1 _09641_/X sky130_fd_sc_hd__a21o_1
XFILLER_283_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18839_ _18608_/Y _18867_/A2 _18837_/Y _18838_/Y vssd1 vssd1 vccd1 vccd1 _18839_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09572_ _12577_/A _13653_/A vssd1 vssd1 vccd1 vccd1 _09572_/X sky130_fd_sc_hd__or2_1
XFILLER_282_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20801_ _21020_/CLK _20801_/D vssd1 vssd1 vccd1 vccd1 _20801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20732_ _20795_/CLK _20732_/D vssd1 vssd1 vccd1 vccd1 _20732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20663_ _20663_/CLK _20663_/D vssd1 vssd1 vccd1 vccd1 _20663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20594_ _20630_/CLK _20594_/D vssd1 vssd1 vccd1 vccd1 _20594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1507 _11818_/B2 vssd1 vssd1 vccd1 vccd1 _11916_/S sky130_fd_sc_hd__buf_6
XFILLER_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout520 _17642_/X vssd1 vssd1 vccd1 vccd1 _17671_/S sky130_fd_sc_hd__clkbuf_16
Xfanout1518 fanout1522/X vssd1 vssd1 vccd1 vccd1 _12139_/S sky130_fd_sc_hd__buf_6
Xfanout531 _17574_/X vssd1 vssd1 vccd1 vccd1 _17606_/S sky130_fd_sc_hd__clkbuf_8
Xfanout1529 _10425_/S vssd1 vssd1 vccd1 vccd1 _10428_/S sky130_fd_sc_hd__buf_6
Xfanout542 _17178_/S vssd1 vssd1 vccd1 vccd1 _17166_/S sky130_fd_sc_hd__buf_12
XFILLER_265_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09908_ _11851_/A _19918_/Q _12188_/S _20043_/Q vssd1 vssd1 vccd1 vccd1 _09908_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_76_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout553 _17049_/X vssd1 vssd1 vccd1 vccd1 _17076_/S sky130_fd_sc_hd__buf_6
Xfanout564 _16605_/X vssd1 vssd1 vccd1 vccd1 _16634_/S sky130_fd_sc_hd__buf_12
XFILLER_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout575 _16456_/X vssd1 vssd1 vccd1 vccd1 _16471_/S sky130_fd_sc_hd__buf_12
Xfanout586 _16068_/Y vssd1 vssd1 vccd1 vccd1 _16106_/A2 sky130_fd_sc_hd__buf_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20028_ _20061_/CLK _20028_/D vssd1 vssd1 vccd1 vccd1 _20028_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout597 _14685_/S vssd1 vssd1 vccd1 vccd1 _14702_/S sky130_fd_sc_hd__buf_12
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09839_ _09839_/A _09839_/B vssd1 vssd1 vccd1 vccd1 _09839_/X sky130_fd_sc_hd__or2_1
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12850_ _12850_/A1 _12832_/B _13350_/A _12710_/B vssd1 vssd1 vccd1 vccd1 _12852_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _11795_/A _11795_/B _11800_/X vssd1 vssd1 vccd1 vccd1 _11804_/A sky130_fd_sc_hd__a21o_1
XFILLER_262_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_wb_clk_i ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _19503_/Q _12781_/B vssd1 vssd1 vccd1 vccd1 _12782_/B sky130_fd_sc_hd__nor2_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _19298_/Q _17674_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19298_/D sky130_fd_sc_hd__mux2_1
XFILLER_214_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11791_/A _11791_/B _11731_/X vssd1 vssd1 vccd1 vccd1 _11795_/A sky130_fd_sc_hd__a21o_2
XFILLER_215_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _20221_/Q _19250_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14452_/B sky130_fd_sc_hd__mux2_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _12051_/A1 _19480_/Q _19448_/Q _11978_/S _12051_/C1 vssd1 vssd1 vccd1 vccd1
+ _11663_/X sky130_fd_sc_hd__a221o_1
XFILLER_230_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _12715_/Y _12726_/C _13377_/Y split6/X vssd1 vssd1 vccd1 vccd1 _13402_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17170_ _20136_/Q _17695_/A1 _17178_/S vssd1 vssd1 vccd1 vccd1 _20136_/D sky130_fd_sc_hd__mux2_1
X_10614_ _12711_/A _20666_/Q _10405_/C _10629_/A vssd1 vssd1 vccd1 vccd1 _10614_/X
+ sky130_fd_sc_hd__o31a_1
X_14382_ _19520_/Q _14383_/B vssd1 vssd1 vccd1 vccd1 _14382_/Y sky130_fd_sc_hd__nor2_1
X_11594_ _11981_/C1 _11593_/X _11590_/X _12137_/C1 vssd1 vssd1 vccd1 vccd1 _11594_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_128_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16121_ _19585_/Q _16127_/A2 _16131_/B1 vssd1 vssd1 vccd1 vccd1 _16121_/X sky130_fd_sc_hd__o21a_1
X_13333_ _13332_/B _13347_/A _13332_/A vssd1 vssd1 vccd1 vccd1 _13334_/C sky130_fd_sc_hd__a21oi_1
X_10545_ input170/X input142/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10545_/X sky130_fd_sc_hd__mux2_8
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16052_ _16052_/A1 _16050_/X _16051_/Y _13181_/B _16052_/B2 vssd1 vssd1 vccd1 vccd1
+ _16052_/X sky130_fd_sc_hd__a32o_1
XFILLER_155_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ _13264_/A _13264_/B _13264_/C vssd1 vssd1 vccd1 vccd1 _13264_/X sky130_fd_sc_hd__and3_1
XFILLER_109_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10476_ _20128_/Q _20096_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _10476_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15003_ _20850_/Q _15601_/S _14998_/X _14993_/X _15002_/X vssd1 vssd1 vccd1 vccd1
+ _15003_/X sky130_fd_sc_hd__o221a_1
XFILLER_68_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12215_ _20586_/Q _12213_/B _12214_/X _12371_/C1 vssd1 vssd1 vccd1 vccd1 _12215_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13195_ _13195_/A _13195_/B vssd1 vssd1 vccd1 vccd1 _13195_/Y sky130_fd_sc_hd__nor2_1
XFILLER_269_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19811_ _20341_/CLK _19811_/D vssd1 vssd1 vccd1 vccd1 _19811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_269_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12146_ _19826_/Q _19330_/Q _12146_/S vssd1 vssd1 vccd1 vccd1 _12146_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19742_ _20763_/CLK _19742_/D vssd1 vssd1 vccd1 vccd1 _19742_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16954_ _19985_/Q _17012_/A2 _16953_/Y _17012_/C1 vssd1 vssd1 vccd1 vccd1 _19985_/D
+ sky130_fd_sc_hd__a211o_1
X_12077_ _12513_/A _11649_/S _12076_/Y vssd1 vssd1 vccd1 vccd1 _12110_/A sky130_fd_sc_hd__o21a_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11028_ _20400_/Q _20336_/Q _20628_/Q _20592_/Q _11035_/S _11021_/C vssd1 vssd1 vccd1
+ vccd1 _11028_/X sky130_fd_sc_hd__mux4_1
X_15905_ _19728_/Q _15961_/A2 _15961_/B1 _19760_/Q vssd1 vssd1 vccd1 vccd1 _15905_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_238_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19673_ _20711_/CLK _19673_/D vssd1 vssd1 vccd1 vccd1 _19673_/Q sky130_fd_sc_hd__dfxtp_1
X_16885_ _16885_/A _16885_/B vssd1 vssd1 vccd1 vccd1 _16885_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18624_ _19509_/Q _18628_/B vssd1 vssd1 vccd1 vccd1 _18624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_266_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _16051_/A1 _15822_/X _16051_/B1 vssd1 vssd1 vccd1 vccd1 _15836_/Y sky130_fd_sc_hd__o21ai_1
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18555_ _18966_/A _18555_/B vssd1 vssd1 vccd1 vccd1 _20911_/D sky130_fd_sc_hd__nor2_1
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12979_ _12979_/A vssd1 vssd1 vccd1 vccd1 _14110_/C sky130_fd_sc_hd__inv_2
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _15219_/Y _15762_/Y _15763_/Y _15766_/X vssd1 vssd1 vccd1 vccd1 _15767_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17506_ _20288_/Q _17522_/B vssd1 vssd1 vccd1 vccd1 _17506_/Y sky130_fd_sc_hd__nand2_1
X_14718_ _19475_/Q _17933_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19475_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18486_ _18589_/B _18487_/B vssd1 vssd1 vccd1 vccd1 _18486_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_480 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15698_ _15941_/B2 _15687_/X _15688_/X _15697_/X vssd1 vssd1 vccd1 vccd1 _15698_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_491 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_268_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17437_ _17441_/C _17457_/C _17423_/X _14440_/Y vssd1 vssd1 vccd1 vccd1 _17437_/X
+ sky130_fd_sc_hd__a211o_1
X_14649_ _19411_/Q _17933_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19411_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_16 _16833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_27 _15725_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_38 _16739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 _16895_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17368_ _20232_/Q _17378_/A2 _17370_/B1 _20281_/Q _17370_/C1 vssd1 vssd1 vccd1 vccd1
+ _17368_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19107_ _19523_/CLK _19107_/D vssd1 vssd1 vccd1 vccd1 _19107_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16319_ _19715_/Q _16322_/C _18086_/A vssd1 vssd1 vccd1 vccd1 _16319_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17299_ _17299_/A _17329_/S _17305_/C vssd1 vssd1 vccd1 vccd1 _17299_/X sky130_fd_sc_hd__and3_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19038_ _18290_/Y _19046_/A2 _19048_/B1 _12550_/D _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19038_/X sky130_fd_sc_hd__a221o_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21000_ _21000_/CLK _21000_/D vssd1 vssd1 vccd1 vccd1 _21000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09624_ _10308_/S _14112_/B vssd1 vssd1 vccd1 vccd1 _09624_/Y sky130_fd_sc_hd__nor2_8
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09555_ _14895_/A _19156_/Q _09555_/C _09567_/A vssd1 vssd1 vccd1 vccd1 _12569_/A
+ sky130_fd_sc_hd__or4_4
Xclkbuf_leaf_37_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20703_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _19993_/Q vssd1 vssd1 vccd1 vccd1 _09486_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20715_ _20715_/CLK _20715_/D vssd1 vssd1 vccd1 vccd1 _20715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20646_ _20646_/CLK _20646_/D vssd1 vssd1 vccd1 vccd1 _20646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20577_ _20714_/CLK _20577_/D vssd1 vssd1 vccd1 vccd1 _20577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10330_ _12403_/A1 _13693_/A _12403_/B1 vssd1 vssd1 vccd1 vccd1 _10330_/X sky130_fd_sc_hd__o21a_1
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10261_ _10262_/A _19912_/Q _11303_/S _20037_/Q vssd1 vssd1 vccd1 vccd1 _10261_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout2005 _16875_/B2 vssd1 vssd1 vccd1 vccd1 _16866_/B2 sky130_fd_sc_hd__clkbuf_4
X_12000_ _12403_/A1 _11999_/Y _12403_/B1 vssd1 vssd1 vccd1 vccd1 _12000_/Y sky130_fd_sc_hd__o21ai_1
X_10192_ _10186_/X _10191_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _10192_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1304 _13468_/B vssd1 vssd1 vccd1 vccd1 _17008_/B1 sky130_fd_sc_hd__buf_6
Xfanout1315 _14853_/S vssd1 vssd1 vccd1 vccd1 _14822_/S sky130_fd_sc_hd__clkbuf_4
Xfanout1326 _15365_/A vssd1 vssd1 vccd1 vccd1 _15220_/A sky130_fd_sc_hd__buf_8
Xfanout1337 _11192_/A2 vssd1 vssd1 vccd1 vccd1 _11392_/A2 sky130_fd_sc_hd__buf_4
Xfanout1348 _17364_/A2 vssd1 vssd1 vccd1 vccd1 _17356_/A2 sky130_fd_sc_hd__buf_6
XFILLER_143_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1359 _14038_/B1 vssd1 vssd1 vccd1 vccd1 _14035_/B1 sky130_fd_sc_hd__buf_4
XFILLER_247_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13951_ _13853_/B _13960_/A2 _11141_/X _13853_/Y _19832_/Q vssd1 vssd1 vccd1 vccd1
+ _14047_/C sky130_fd_sc_hd__o32a_1
XFILLER_98_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12902_ _12902_/A vssd1 vssd1 vccd1 vccd1 _12902_/Y sky130_fd_sc_hd__inv_2
X_16670_ _19927_/Q _17114_/A1 _16670_/S vssd1 vssd1 vccd1 vccd1 _19927_/D sky130_fd_sc_hd__mux2_1
X_13882_ _19100_/Q _14738_/B _13889_/B1 _15649_/A1 _16171_/A vssd1 vssd1 vccd1 vccd1
+ _19100_/D sky130_fd_sc_hd__o221a_1
XFILLER_98_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_261_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ _15686_/A _15526_/A vssd1 vssd1 vccd1 vccd1 _12833_/Y sky130_fd_sc_hd__nand2_2
X_15621_ _13426_/A _15620_/Y _16034_/S vssd1 vssd1 vccd1 vccd1 _15621_/X sky130_fd_sc_hd__mux2_1
XFILLER_262_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18340_ _20825_/Q _18349_/B _18339_/Y _18710_/A vssd1 vssd1 vccd1 vccd1 _20825_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _13426_/C _15259_/B _16056_/B1 _15551_/X vssd1 vssd1 vccd1 vccd1 _15552_/X
+ sky130_fd_sc_hd__a211o_1
X_12764_ _15443_/A _12784_/B vssd1 vssd1 vccd1 vccd1 _12764_/Y sky130_fd_sc_hd__nand2_2
XFILLER_226_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14503_ _19281_/Q _17934_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19281_/D sky130_fd_sc_hd__mux2_1
X_11715_ _11718_/S _11712_/X _11714_/X vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__a21o_1
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15483_ _20797_/Q _16047_/A2 _15481_/X _15482_/X vssd1 vssd1 vccd1 vccd1 _15483_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_188_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18271_ _20808_/Q _18270_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18272_/B sky130_fd_sc_hd__mux2_1
X_12695_ _12513_/A _13589_/A1 _12642_/Y _12643_/X vssd1 vssd1 vccd1 vccd1 _12698_/D
+ sky130_fd_sc_hd__a211oi_2
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17222_ _20183_/Q _17224_/B vssd1 vssd1 vccd1 vccd1 _17222_/X sky130_fd_sc_hd__or2_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14434_ _14433_/A _14433_/B _14433_/Y _14427_/A vssd1 vssd1 vccd1 vccd1 _14435_/B
+ sky130_fd_sc_hd__a211o_1
X_11646_ _11646_/A _11646_/B vssd1 vssd1 vccd1 vccd1 _11646_/Y sky130_fd_sc_hd__nand2_2
XFILLER_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 core_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_4
X_17153_ _20119_/Q _17678_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20119_/D sky130_fd_sc_hd__mux2_1
X_14365_ _14363_/Y _14365_/B vssd1 vssd1 vccd1 vccd1 _14366_/B sky130_fd_sc_hd__nand2b_1
XFILLER_11_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput25 core_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_4
Xinput36 core_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_6
X_11577_ _20384_/Q _20448_/Q _11979_/S vssd1 vssd1 vccd1 vccd1 _11577_/X sky130_fd_sc_hd__mux2_1
Xinput47 dout0[13] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_2
X_16104_ _10551_/X _16132_/A2 _16103_/X vssd1 vssd1 vccd1 vccd1 _19576_/D sky130_fd_sc_hd__o21a_1
Xinput58 dout0[23] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
X_13316_ _13316_/A _13316_/B vssd1 vssd1 vccd1 vccd1 _13316_/X sky130_fd_sc_hd__or2_2
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17084_ _20054_/Q _17852_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20054_/D sky130_fd_sc_hd__mux2_1
X_10528_ _19808_/Q _11291_/A2 _10526_/X _11291_/B2 _10527_/X vssd1 vssd1 vccd1 vccd1
+ _10528_/X sky130_fd_sc_hd__o221a_1
XFILLER_128_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput69 dout0[33] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_2
X_14296_ _14296_/A _14397_/A _14397_/B vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__or3_1
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ _13346_/A _13346_/B _13332_/A _13346_/C vssd1 vssd1 vccd1 vccd1 _13321_/C
+ sky130_fd_sc_hd__a211o_1
X_16035_ _12517_/B _16063_/A2 _16007_/A vssd1 vssd1 vccd1 vccd1 _16035_/X sky130_fd_sc_hd__a21bo_1
XFILLER_108_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10459_ _11228_/A1 _13978_/A2 _10458_/X _11239_/B1 _19841_/Q vssd1 vssd1 vccd1 vccd1
+ _10459_/X sky130_fd_sc_hd__o32a_1
XFILLER_254_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13178_ _13178_/A _13178_/B vssd1 vssd1 vccd1 vccd1 _13181_/A sky130_fd_sc_hd__xnor2_4
XFILLER_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12129_ _12125_/X _12128_/X _12129_/S vssd1 vssd1 vccd1 vccd1 _12129_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17986_ _18080_/A _17991_/C vssd1 vssd1 vccd1 vccd1 _17986_/Y sky130_fd_sc_hd__nor2_1
XFILLER_257_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19725_ _19970_/CLK _19725_/D vssd1 vssd1 vccd1 vccd1 _19725_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1860 _18765_/B vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16937_ _20420_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16937_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1871 _19166_/Q vssd1 vssd1 vccd1 vccd1 _15649_/A1 sky130_fd_sc_hd__buf_6
XFILLER_272_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1882 _19162_/Q vssd1 vssd1 vccd1 vccd1 _12510_/C sky130_fd_sc_hd__buf_8
Xfanout1893 _18752_/A vssd1 vssd1 vccd1 vccd1 _17393_/C1 sky130_fd_sc_hd__buf_4
XFILLER_38_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19656_ _20410_/CLK _19656_/D vssd1 vssd1 vccd1 vccd1 _19656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16868_ _19975_/Q _16887_/A _16867_/Y _16896_/C1 vssd1 vssd1 vccd1 vccd1 _19975_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18607_ _20925_/Q _18619_/B vssd1 vssd1 vccd1 vccd1 _18607_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15819_ _13413_/A _12565_/B _15818_/X vssd1 vssd1 vccd1 vccd1 _15819_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19587_ _19589_/CLK _19587_/D vssd1 vssd1 vccd1 vccd1 _19587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16799_ input104/X input75/X _16799_/S vssd1 vssd1 vccd1 vccd1 _16800_/A sky130_fd_sc_hd__mux2_2
XFILLER_252_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18538_ _18651_/B _18538_/B vssd1 vssd1 vccd1 vccd1 _18538_/X sky130_fd_sc_hd__or2_1
XFILLER_280_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18469_ _18467_/Y _18468_/X _18476_/A vssd1 vssd1 vccd1 vccd1 _20884_/D sky130_fd_sc_hd__o21a_1
X_20500_ _20664_/CLK _20500_/D vssd1 vssd1 vccd1 vccd1 _20500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20431_ _20463_/CLK _20431_/D vssd1 vssd1 vccd1 vccd1 _20431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_155_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19759_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20362_ _20686_/CLK _20362_/D vssd1 vssd1 vccd1 vccd1 _20362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20293_ _20296_/CLK _20293_/D vssd1 vssd1 vccd1 vccd1 _20293_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_161_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09607_ _12975_/A _09607_/B _12976_/A vssd1 vssd1 vccd1 vccd1 _09607_/X sky130_fd_sc_hd__and3b_4
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09538_ _19152_/Q _19151_/Q _19150_/Q vssd1 vssd1 vccd1 vccd1 _12480_/B sky130_fd_sc_hd__and3_2
XFILLER_231_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11500_ _19945_/Q _11897_/B vssd1 vssd1 vccd1 vccd1 _11500_/X sky130_fd_sc_hd__or2_1
XFILLER_269_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12480_ _12480_/A _12480_/B _13867_/A vssd1 vssd1 vccd1 vccd1 _15220_/B sky130_fd_sc_hd__and3_4
XFILLER_40_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _11429_/X _11430_/X _12134_/S vssd1 vssd1 vccd1 vccd1 _11431_/X sky130_fd_sc_hd__mux2_2
XFILLER_184_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20629_ _20667_/CLK _20629_/D vssd1 vssd1 vccd1 vccd1 _20629_/Q sky130_fd_sc_hd__dfxtp_1
X_14150_ _14141_/A _14138_/Y _14140_/B vssd1 vssd1 vccd1 vccd1 _14160_/B sky130_fd_sc_hd__o21ai_2
XFILLER_138_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ _12301_/S _11361_/X _11360_/X _12314_/C1 vssd1 vssd1 vccd1 vccd1 _11362_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ _13091_/A _13091_/B _13091_/C vssd1 vssd1 vccd1 vccd1 _13101_/Y sky130_fd_sc_hd__a21oi_1
X_10313_ _11266_/A1 _20507_/Q _11256_/S _10312_/X vssd1 vssd1 vccd1 vccd1 _10313_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14081_ _14081_/A _16133_/B _14081_/C vssd1 vssd1 vccd1 vccd1 _14081_/X sky130_fd_sc_hd__or3_1
XFILLER_3_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11293_ _11291_/X _11292_/X _11297_/S vssd1 vssd1 vccd1 vccd1 _11293_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13032_ _20962_/Q _20896_/Q vssd1 vssd1 vccd1 vccd1 _13353_/B sky130_fd_sc_hd__nand2_1
X_10244_ _12711_/A _15922_/B2 _10243_/X vssd1 vssd1 vccd1 vccd1 _10277_/A sky130_fd_sc_hd__a21oi_4
XFILLER_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1101 _17178_/A1 vssd1 vssd1 vccd1 vccd1 _17946_/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout1112 _17944_/A1 vssd1 vssd1 vccd1 vccd1 _17804_/A1 sky130_fd_sc_hd__clkbuf_4
X_17840_ _20615_/Q _17878_/A1 _17840_/S vssd1 vssd1 vccd1 vccd1 _20615_/D sky130_fd_sc_hd__mux2_1
XFILLER_239_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10175_ _10173_/X _10174_/X _11378_/S vssd1 vssd1 vccd1 vccd1 _10175_/X sky130_fd_sc_hd__mux2_1
XFILLER_267_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1123 _11612_/X vssd1 vssd1 vccd1 vccd1 _17905_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_239_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1134 _17893_/A1 vssd1 vssd1 vccd1 vccd1 _17927_/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1145 _17908_/A1 vssd1 vssd1 vccd1 vccd1 _17802_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1156 _09632_/Y vssd1 vssd1 vccd1 vccd1 _12402_/A1 sky130_fd_sc_hd__buf_12
XFILLER_120_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17771_ _20550_/Q _17911_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20550_/D sky130_fd_sc_hd__mux2_1
Xfanout1167 _16050_/A1 vssd1 vssd1 vccd1 vccd1 _15973_/A1 sky130_fd_sc_hd__buf_4
X_14983_ _14983_/A _14987_/B vssd1 vssd1 vccd1 vccd1 _14983_/Y sky130_fd_sc_hd__nor2_1
Xfanout1178 _13350_/B vssd1 vssd1 vccd1 vccd1 _13366_/C1 sky130_fd_sc_hd__buf_2
XFILLER_282_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1189 _10385_/A vssd1 vssd1 vccd1 vccd1 _10127_/A sky130_fd_sc_hd__buf_6
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19510_ _19511_/CLK _19510_/D vssd1 vssd1 vccd1 vccd1 _19510_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_235_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16722_ _19215_/Q _16996_/A2 _16996_/B1 _19084_/Q _16721_/X vssd1 vssd1 vccd1 vccd1
+ _16722_/X sky130_fd_sc_hd__o221a_1
X_13934_ _19138_/Q _13941_/B _13946_/B1 _13412_/B vssd1 vssd1 vccd1 vccd1 _19138_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_263_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19441_ _20711_/CLK _19441_/D vssd1 vssd1 vccd1 vccd1 _19441_/Q sky130_fd_sc_hd__dfxtp_1
X_16653_ _19910_/Q _17097_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19910_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13865_ _19085_/Q _13863_/B _13881_/B1 _19151_/Q _15288_/C1 vssd1 vssd1 vccd1 vccd1
+ _19085_/D sky130_fd_sc_hd__o221a_1
XFILLER_263_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15604_ _19749_/Q _15604_/A2 _15603_/X _16048_/C1 vssd1 vssd1 vccd1 vccd1 _15604_/X
+ sky130_fd_sc_hd__a211o_1
X_19372_ _20663_/CLK _19372_/D vssd1 vssd1 vccd1 vccd1 _19372_/Q sky130_fd_sc_hd__dfxtp_1
X_12816_ _19516_/Q _12804_/B _19517_/Q vssd1 vssd1 vccd1 vccd1 _12817_/B sky130_fd_sc_hd__a21oi_1
X_16584_ _19858_/Q _16592_/A2 _16592_/B1 input29/X vssd1 vssd1 vccd1 vccd1 _16585_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13796_ _13802_/A1 _13656_/B _13805_/B1 input242/X vssd1 vssd1 vccd1 vccd1 _13796_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18323_ _18981_/B _18323_/B _18154_/B vssd1 vssd1 vccd1 vccd1 _18324_/B sky130_fd_sc_hd__or3b_4
XFILLER_72_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15535_ _20959_/Q _15939_/A2 _15996_/B1 _20831_/Q _15534_/X vssd1 vssd1 vccd1 vccd1
+ _15535_/X sky130_fd_sc_hd__a221o_4
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12747_/A _12747_/B _12747_/C vssd1 vssd1 vccd1 vccd1 _12748_/B sky130_fd_sc_hd__nand3_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18254_ _18313_/B _14312_/B _18253_/Y vssd1 vssd1 vccd1 vccd1 _18523_/B sky130_fd_sc_hd__o21ai_4
X_12678_ _13501_/B _12678_/B vssd1 vssd1 vccd1 vccd1 _13511_/A sky130_fd_sc_hd__and2b_1
X_15466_ _15163_/Y _15175_/B _15611_/S vssd1 vssd1 vccd1 vccd1 _15466_/X sky130_fd_sc_hd__mux2_1
X_17205_ _20169_/Q _17696_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20169_/D sky130_fd_sc_hd__mux2_1
X_14417_ _14413_/B _14416_/Y _14417_/S vssd1 vssd1 vccd1 vccd1 _14417_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11629_ _11872_/A _12023_/S _11626_/X _11628_/X vssd1 vssd1 vccd1 vccd1 _11629_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18185_ _18480_/B vssd1 vssd1 vccd1 vccd1 _18185_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15397_ _15282_/A _16804_/B _15380_/Y vssd1 vssd1 vccd1 vccd1 _15397_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_156_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17136_ _20104_/Q _17695_/A1 _17144_/S vssd1 vssd1 vccd1 vccd1 _20104_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14348_ _14437_/A _14437_/B _14348_/C vssd1 vssd1 vccd1 vccd1 _14348_/X sky130_fd_sc_hd__or3_1
XFILLER_265_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17067_ _20039_/Q _17903_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20039_/D sky130_fd_sc_hd__mux2_1
X_14279_ _20282_/Q _14330_/A2 _14330_/B1 input222/X vssd1 vssd1 vccd1 vccd1 _14281_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_171_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16018_ _20880_/Q _16018_/A2 _16017_/X vssd1 vssd1 vccd1 vccd1 _16018_/X sky130_fd_sc_hd__o21a_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _20727_/Q _17971_/C _17968_/Y vssd1 vssd1 vccd1 vccd1 _20727_/D sky130_fd_sc_hd__o21a_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19708_ _20757_/CLK _19708_/D vssd1 vssd1 vccd1 vccd1 _19708_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1690 _10937_/A vssd1 vssd1 vccd1 vccd1 _10356_/A sky130_fd_sc_hd__buf_6
XFILLER_66_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20980_ _20980_/CLK _20980_/D vssd1 vssd1 vccd1 vccd1 _20980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19639_ _20673_/CLK _19639_/D vssd1 vssd1 vccd1 vccd1 _19639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20414_ _20425_/CLK _20414_/D vssd1 vssd1 vccd1 vccd1 _20414_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20345_ _20683_/CLK _20345_/D vssd1 vssd1 vccd1 vccd1 _20345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20276_ _21013_/CLK _20276_/D vssd1 vssd1 vccd1 vccd1 _20276_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_161_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput204 localMemory_wb_adr_i[22] vssd1 vssd1 vccd1 vccd1 _12928_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_49_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput215 localMemory_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_hd__buf_12
XFILLER_103_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput226 localMemory_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_hd__buf_12
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput237 localMemory_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_hd__buf_12
XFILLER_102_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20491_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 localMemory_wb_sel_i[1] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput259 manufacturerID[5] vssd1 vssd1 vccd1 vccd1 _17254_/A sky130_fd_sc_hd__buf_2
XFILLER_276_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ _11978_/X _11979_/X _11980_/S vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__mux2_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10931_ _12569_/A _13650_/B _10930_/Y _11281_/B vssd1 vssd1 vccd1 vccd1 _10931_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_95_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10862_ _10856_/X _10861_/X _12415_/S vssd1 vssd1 vccd1 vccd1 _10862_/X sky130_fd_sc_hd__mux2_1
XFILLER_231_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13650_ _13657_/A _13650_/B vssd1 vssd1 vccd1 vccd1 _13685_/B sky130_fd_sc_hd__nor2_8
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _19503_/Q _12781_/B vssd1 vssd1 vccd1 vccd1 _12782_/A sky130_fd_sc_hd__and2_2
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13581_ _18462_/A _13579_/X _13580_/X vssd1 vssd1 vccd1 vccd1 _13581_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _11375_/S _10792_/X _10789_/X _12431_/A1 vssd1 vssd1 vccd1 vccd1 _10794_/B
+ sky130_fd_sc_hd__o211a_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15320_ _19708_/Q _15454_/S _15307_/X _15319_/X _14941_/X vssd1 vssd1 vccd1 vccd1
+ _15320_/X sky130_fd_sc_hd__o221a_2
XFILLER_213_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12532_ _19118_/Q _19117_/Q vssd1 vssd1 vccd1 vccd1 _12532_/X sky130_fd_sc_hd__or2_1
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15251_ _15048_/X _15037_/X _15254_/S vssd1 vssd1 vccd1 vccd1 _15251_/X sky130_fd_sc_hd__mux2_1
X_12463_ _12463_/A _12463_/B vssd1 vssd1 vccd1 vccd1 _12463_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14202_ _14198_/B _14201_/Y _14202_/S vssd1 vssd1 vccd1 vccd1 _14202_/X sky130_fd_sc_hd__mux2_1
X_11414_ _10365_/A _11414_/B vssd1 vssd1 vccd1 vccd1 _11415_/B sky130_fd_sc_hd__nand2b_1
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15182_ _15610_/A1 _15181_/X _15610_/B1 vssd1 vssd1 vccd1 vccd1 _15182_/Y sky130_fd_sc_hd__o21ai_1
X_12394_ _19828_/Q _19332_/Q _12397_/S vssd1 vssd1 vccd1 vccd1 _12394_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14133_ _18152_/B _14132_/X _12523_/X vssd1 vssd1 vccd1 vccd1 _14134_/C sky130_fd_sc_hd__o21ba_1
X_11345_ _11343_/X _11344_/X _11345_/S vssd1 vssd1 vccd1 vccd1 _11345_/X sky130_fd_sc_hd__mux2_1
X_19990_ _20860_/CLK _19990_/D vssd1 vssd1 vccd1 vccd1 _19990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14064_ _19191_/Q _14082_/A2 _14063_/X _16087_/B1 vssd1 vssd1 vccd1 vccd1 _19191_/D
+ sky130_fd_sc_hd__o211a_1
X_18941_ _18975_/A _18941_/B vssd1 vssd1 vccd1 vccd1 _18941_/Y sky130_fd_sc_hd__nand2_1
X_11276_ _09689_/C _11264_/X _11267_/X _11275_/X _12311_/C1 vssd1 vssd1 vccd1 vccd1
+ _11276_/X sky130_fd_sc_hd__o311a_1
XFILLER_134_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13015_ _20971_/Q _20905_/Q vssd1 vssd1 vccd1 vccd1 _13015_/X sky130_fd_sc_hd__or2_4
X_10227_ _20640_/Q _20604_/Q _10986_/B vssd1 vssd1 vccd1 vccd1 _10227_/X sky130_fd_sc_hd__mux2_1
X_18872_ _18968_/A _18872_/B vssd1 vssd1 vccd1 vccd1 _18872_/Y sky130_fd_sc_hd__nand2_1
XFILLER_279_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17823_ _20598_/Q _17861_/A1 _17840_/S vssd1 vssd1 vccd1 vccd1 _20598_/D sky130_fd_sc_hd__mux2_1
X_10158_ _19280_/Q _20067_/Q _12296_/S vssd1 vssd1 vccd1 vccd1 _10158_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17754_ _20533_/Q _17894_/A1 _17776_/S vssd1 vssd1 vccd1 vccd1 _20533_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14966_ _14973_/A _14973_/B _14966_/C vssd1 vssd1 vccd1 vccd1 _15314_/D sky130_fd_sc_hd__or3_4
X_10089_ _19410_/Q _20569_/Q _10518_/S vssd1 vssd1 vccd1 vccd1 _10089_/X sky130_fd_sc_hd__mux2_1
X_16705_ _19960_/Q _17674_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19960_/D sky130_fd_sc_hd__mux2_1
XFILLER_207_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13917_ _19124_/Q _13566_/Y _13919_/S vssd1 vssd1 vccd1 vccd1 _13918_/B sky130_fd_sc_hd__mux2_1
X_17685_ _20469_/Q _17928_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20469_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14897_ _14897_/A _14897_/B vssd1 vssd1 vccd1 vccd1 _14897_/Y sky130_fd_sc_hd__nor2_2
XFILLER_223_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19424_ _20583_/CLK _19424_/D vssd1 vssd1 vccd1 vccd1 _19424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16636_ _19895_/Q _17707_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19895_/D sky130_fd_sc_hd__mux2_1
X_13848_ _17441_/A _17423_/D vssd1 vssd1 vccd1 vccd1 _17421_/A sky130_fd_sc_hd__or2_1
XFILLER_63_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19355_ _20710_/CLK _19355_/D vssd1 vssd1 vccd1 vccd1 _19355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16567_ _16567_/A _16567_/B vssd1 vssd1 vccd1 vccd1 _19849_/D sky130_fd_sc_hd__or2_1
XFILLER_149_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13779_ _13779_/A _13779_/B vssd1 vssd1 vccd1 vccd1 _13780_/B sky130_fd_sc_hd__nor2_8
XFILLER_149_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18306_ _20815_/Q _18305_/Y _18316_/S vssd1 vssd1 vccd1 vccd1 _18307_/B sky130_fd_sc_hd__mux2_1
XFILLER_176_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15518_ _15644_/A1 _16842_/B _15504_/Y vssd1 vssd1 vccd1 vccd1 _15518_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_188_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19286_ _20480_/CLK _19286_/D vssd1 vssd1 vccd1 vccd1 _19286_/Q sky130_fd_sc_hd__dfxtp_1
X_16498_ _19805_/Q _17859_/A1 _16521_/S vssd1 vssd1 vccd1 vccd1 _19805_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18237_ _18422_/A _18237_/B vssd1 vssd1 vccd1 vccd1 _20801_/D sky130_fd_sc_hd__and2_1
X_15449_ _20956_/Q _15568_/A2 _15568_/B1 _20828_/Q _15448_/X vssd1 vssd1 vccd1 vccd1
+ _15449_/X sky130_fd_sc_hd__a221o_4
XFILLER_209_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18168_ _19529_/Q _18213_/B vssd1 vssd1 vccd1 vccd1 _18168_/Y sky130_fd_sc_hd__nand2b_4
XFILLER_144_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17119_ _20087_/Q _17678_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20087_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18099_ _20774_/Q _18101_/C _18098_/Y vssd1 vssd1 vccd1 vccd1 _20774_/D sky130_fd_sc_hd__o21a_1
XFILLER_172_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20130_ _20711_/CLK _20130_/D vssd1 vssd1 vccd1 vccd1 _20130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09941_ _09941_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _13415_/A sky130_fd_sc_hd__and2_4
XFILLER_277_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout905 _15322_/C vssd1 vssd1 vccd1 vccd1 _15568_/A2 sky130_fd_sc_hd__clkbuf_16
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout916 _15934_/B1 vssd1 vssd1 vccd1 vccd1 _16011_/B1 sky130_fd_sc_hd__buf_6
X_20061_ _20061_/CLK _20061_/D vssd1 vssd1 vccd1 vccd1 _20061_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout927 _15989_/A2 vssd1 vssd1 vccd1 vccd1 _15961_/A2 sky130_fd_sc_hd__buf_4
XFILLER_258_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09872_ _20546_/Q _12146_/S vssd1 vssd1 vccd1 vccd1 _09872_/X sky130_fd_sc_hd__or2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout938 _11187_/X vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__buf_4
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout949 _10933_/Y vssd1 vssd1 vccd1 vccd1 _15066_/S sky130_fd_sc_hd__buf_8
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_7__f_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_7__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_227_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_309 input236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20963_ _21030_/CLK _20963_/D vssd1 vssd1 vccd1 vccd1 _20963_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ _20959_/CLK _20894_/D vssd1 vssd1 vccd1 vccd1 _20894_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_213_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_170_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21042_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ _11309_/A1 _11125_/X _11129_/X _12431_/A1 vssd1 vssd1 vccd1 vccd1 _11131_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20328_ _20716_/CLK _20328_/D vssd1 vssd1 vccd1 vccd1 _20328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11061_ _11061_/A _16073_/A vssd1 vssd1 vccd1 vccd1 _11061_/Y sky130_fd_sc_hd__nor2_1
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20259_ _20425_/CLK _20259_/D vssd1 vssd1 vccd1 vccd1 _20259_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_49_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ _10003_/X _10011_/Y _12192_/A1 _09995_/X vssd1 vssd1 vccd1 vccd1 _10012_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _14818_/X _14819_/X _15039_/A vssd1 vssd1 vccd1 vccd1 _14820_/X sky130_fd_sc_hd__mux2_1
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _19500_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14751_/X sky130_fd_sc_hd__or2_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ _12039_/A1 _10382_/B _10037_/B vssd1 vssd1 vccd1 vccd1 _11963_/X sky130_fd_sc_hd__a21o_4
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _16598_/C _13702_/B vssd1 vssd1 vccd1 vccd1 _13702_/Y sky130_fd_sc_hd__nor2_1
X_10914_ _09618_/A _20693_/Q _12296_/S _10912_/X _10913_/X vssd1 vssd1 vccd1 vccd1
+ _10914_/X sky130_fd_sc_hd__a311o_1
X_17470_ _20270_/Q _17494_/B vssd1 vssd1 vccd1 vccd1 _17470_/Y sky130_fd_sc_hd__nand2_1
XFILLER_244_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _19441_/Q _17163_/A1 _14699_/S vssd1 vssd1 vccd1 vccd1 _19441_/D sky130_fd_sc_hd__mux2_1
X_11894_ _11977_/A1 _20714_/Q _11891_/B _11893_/X vssd1 vssd1 vccd1 vccd1 _11894_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16421_ _18104_/A _16426_/C vssd1 vssd1 vccd1 vccd1 _16421_/Y sky130_fd_sc_hd__nor2_1
X_10845_ _12314_/C1 _10844_/X _10841_/X _12399_/C1 vssd1 vssd1 vccd1 vccd1 _10845_/X
+ sky130_fd_sc_hd__o211a_1
X_13633_ _13658_/A _16054_/B _15076_/A _14525_/B vssd1 vssd1 vccd1 vccd1 _16235_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_232_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19140_ _20291_/CLK _19140_/D vssd1 vssd1 vccd1 vccd1 _19140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16352_ _19727_/Q _16354_/C _16351_/Y vssd1 vssd1 vccd1 vccd1 _19727_/D sky130_fd_sc_hd__o21a_1
X_10776_ _10774_/X _10775_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _10776_/X sky130_fd_sc_hd__mux2_2
XFILLER_157_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13564_ _20953_/Q _13564_/B vssd1 vssd1 vccd1 vccd1 _13564_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15303_ _15303_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15303_/Y sky130_fd_sc_hd__nand2_1
X_12515_ _12519_/A _12515_/B _12515_/C _11367_/A vssd1 vssd1 vccd1 vccd1 _12516_/C
+ sky130_fd_sc_hd__or4b_2
X_19071_ _20416_/Q vssd1 vssd1 vccd1 vccd1 _20416_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_201_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13495_ _13495_/A _13495_/B vssd1 vssd1 vccd1 vccd1 _15185_/A sky130_fd_sc_hd__xnor2_4
X_16283_ _20624_/Q _17015_/B _19701_/D vssd1 vssd1 vccd1 vccd1 _19699_/D sky130_fd_sc_hd__and3_1
XFILLER_157_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18022_ _18112_/A _18022_/B vssd1 vssd1 vccd1 vccd1 _18022_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15234_ _20886_/Q _15322_/A _15323_/B _15233_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15234_/X sky130_fd_sc_hd__a221o_1
X_12446_ _12446_/A vssd1 vssd1 vccd1 vccd1 _12449_/C sky130_fd_sc_hd__inv_2
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12377_ _12373_/X _12376_/X _12377_/S vssd1 vssd1 vccd1 vccd1 _12377_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15165_ _15044_/X _15046_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _15166_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11328_ _10037_/Y _11230_/Y _09669_/X vssd1 vssd1 vccd1 vccd1 _11328_/X sky130_fd_sc_hd__a21o_1
X_14116_ _14397_/A _14397_/B vssd1 vssd1 vccd1 vccd1 _14116_/Y sky130_fd_sc_hd__nor2_1
X_19973_ _20004_/CLK _19973_/D vssd1 vssd1 vccd1 vccd1 _19973_/Q sky130_fd_sc_hd__dfxtp_1
X_15096_ _15096_/A _15096_/B vssd1 vssd1 vccd1 vccd1 _15096_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18924_ _18535_/X _18971_/B _18922_/X _18923_/Y vssd1 vssd1 vccd1 vccd1 _18925_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_268_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11259_ _11257_/X _11258_/X _11259_/S vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__mux2_1
X_14047_ _14081_/A _16133_/B _14047_/C vssd1 vssd1 vccd1 vccd1 _14047_/X sky130_fd_sc_hd__or3_1
XFILLER_262_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18855_ _18505_/X _18861_/B _18853_/X _18854_/Y vssd1 vssd1 vccd1 vccd1 _18856_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_255_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17806_ _20583_/Q _17806_/A1 _17806_/S vssd1 vssd1 vccd1 vccd1 _20583_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18786_ _18784_/X _18785_/X _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18786_/X sky130_fd_sc_hd__a21o_1
XFILLER_83_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15998_ _20815_/Q _15998_/A2 _15991_/X _16000_/A1 _15997_/X vssd1 vssd1 vccd1 vccd1
+ _15998_/X sky130_fd_sc_hd__a221o_1
X_17737_ _20518_/Q _17911_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20518_/D sky130_fd_sc_hd__mux2_1
XFILLER_78_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ _15019_/A _14947_/X _15453_/A2 _19734_/Q _16048_/C1 vssd1 vssd1 vccd1 vccd1
+ _14949_/X sky130_fd_sc_hd__a221o_2
XFILLER_36_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17668_ _20454_/Q _17805_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20454_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19407_ _20698_/CLK _19407_/D vssd1 vssd1 vccd1 vccd1 _19407_/Q sky130_fd_sc_hd__dfxtp_1
X_16619_ _19878_/Q _17199_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19878_/D sky130_fd_sc_hd__mux2_1
XFILLER_211_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17599_ _20357_/Q _17910_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20357_/D sky130_fd_sc_hd__mux2_1
X_19338_ _20720_/CLK _19338_/D vssd1 vssd1 vccd1 vccd1 _19338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19269_ _20061_/CLK _19269_/D vssd1 vssd1 vccd1 vccd1 _19269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20113_ _20716_/CLK _20113_/D vssd1 vssd1 vccd1 vccd1 _20113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_259_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09924_ _20322_/Q _09928_/S _09923_/X vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__a21o_1
Xfanout702 _13473_/X vssd1 vssd1 vccd1 vccd1 split1/A sky130_fd_sc_hd__buf_8
Xfanout713 _13463_/X vssd1 vssd1 vccd1 vccd1 _16279_/B sky130_fd_sc_hd__buf_12
XFILLER_277_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout724 _13438_/Y vssd1 vssd1 vccd1 vccd1 split3/A sky130_fd_sc_hd__buf_8
XFILLER_258_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout735 _18983_/Y vssd1 vssd1 vccd1 vccd1 _18997_/B sky130_fd_sc_hd__buf_6
XFILLER_59_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout746 _18767_/X vssd1 vssd1 vccd1 vccd1 _18818_/A2 sky130_fd_sc_hd__buf_6
XFILLER_259_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20044_ _20479_/CLK _20044_/D vssd1 vssd1 vccd1 vccd1 _20044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout757 _18769_/Y vssd1 vssd1 vccd1 vccd1 _18937_/B sky130_fd_sc_hd__buf_4
X_09855_ _10516_/S _09850_/X _09854_/X _10260_/S vssd1 vssd1 vccd1 vccd1 _09855_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_259_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout768 _09530_/Y vssd1 vssd1 vccd1 vccd1 _18593_/A2 sky130_fd_sc_hd__buf_6
XFILLER_285_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout779 _18490_/A vssd1 vssd1 vccd1 vccd1 _18616_/B sky130_fd_sc_hd__clkbuf_4
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ input121/X input156/X _11241_/S vssd1 vssd1 vccd1 vccd1 _09786_/X sky130_fd_sc_hd__mux2_8
XFILLER_218_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_106 _12975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_117 _16237_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 _13660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20946_ _21018_/CLK _20946_/D vssd1 vssd1 vccd1 vccd1 _20946_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20877_ _21041_/CLK _20877_/D vssd1 vssd1 vccd1 vccd1 _20877_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10630_ _12711_/A _19471_/Q _19439_/Q _10628_/S _10630_/C1 vssd1 vssd1 vccd1 vccd1
+ _10630_/X sky130_fd_sc_hd__a221o_1
XFILLER_139_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10561_ _10561_/A _10561_/B vssd1 vssd1 vccd1 vccd1 _10561_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12300_ _19693_/Q _20181_/Q _12300_/S vssd1 vssd1 vccd1 vccd1 _12300_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13280_ _13309_/A _13309_/B vssd1 vssd1 vccd1 vccd1 _13281_/B sky130_fd_sc_hd__nand2_1
XFILLER_212_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10492_ _20407_/Q _10502_/A2 _10489_/X _10490_/X _10491_/X vssd1 vssd1 vccd1 vccd1
+ _10492_/X sky130_fd_sc_hd__o221a_1
XFILLER_10_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ _20654_/Q _20618_/Q _12313_/S vssd1 vssd1 vccd1 vccd1 _12231_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12162_ _20553_/Q _20521_/Q _12182_/S vssd1 vssd1 vccd1 vccd1 _12162_/X sky130_fd_sc_hd__mux2_1
XFILLER_269_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11113_ _11111_/X _11112_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _11113_/X sky130_fd_sc_hd__mux2_2
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16970_ _19987_/Q _17012_/A2 _16969_/Y _17012_/C1 vssd1 vssd1 vccd1 vccd1 _19987_/D
+ sky130_fd_sc_hd__a211o_1
X_12093_ _12102_/A1 _19360_/Q _20715_/Q _12097_/S _12100_/B1 vssd1 vssd1 vccd1 vccd1
+ _12093_/X sky130_fd_sc_hd__a221o_1
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ _11021_/A _20121_/Q _20089_/Q _11039_/S vssd1 vssd1 vccd1 vccd1 _11044_/X
+ sky130_fd_sc_hd__a22o_1
X_15921_ _15948_/A1 _12889_/X _15920_/X _15921_/B2 vssd1 vssd1 vccd1 vccd1 _15923_/A
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18640_ _19513_/Q _18671_/B vssd1 vssd1 vccd1 vccd1 _18640_/Y sky130_fd_sc_hd__nand2_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15852_ _20746_/Q _15934_/A2 _15934_/B1 _20778_/Q vssd1 vssd1 vccd1 vccd1 _15852_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_276_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14803_ _14803_/A1 _12478_/Y _13609_/A vssd1 vssd1 vccd1 vccd1 _14803_/Y sky130_fd_sc_hd__o21ai_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _18463_/X _18564_/A _18569_/Y _18570_/Y vssd1 vssd1 vccd1 vccd1 _18572_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _16024_/A1 _15781_/X _15782_/Y _15762_/A _15975_/B2 vssd1 vssd1 vccd1 vccd1
+ _15783_/X sky130_fd_sc_hd__a32o_1
XFILLER_64_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12995_ _19239_/Q _19238_/Q _19237_/Q _13390_/B vssd1 vssd1 vccd1 vccd1 _13231_/B
+ sky130_fd_sc_hd__and4_2
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17522_ _20296_/Q _17522_/B vssd1 vssd1 vccd1 vccd1 _17522_/Y sky130_fd_sc_hd__nand2_1
X_14734_ _19491_/Q _17706_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19491_/D sky130_fd_sc_hd__mux2_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _11946_/A1 _19359_/Q _20714_/Q _11947_/S _11946_/C1 vssd1 vssd1 vccd1 vccd1
+ _11946_/X sky130_fd_sc_hd__a221o_1
XFILLER_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_640 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_651 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _17446_/A _17446_/B _17460_/A2 vssd1 vssd1 vccd1 vccd1 _17454_/D sky130_fd_sc_hd__o21ai_1
X_14665_ _19427_/Q _17949_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19427_/D sky130_fd_sc_hd__mux2_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11877_ _11877_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11878_/B sky130_fd_sc_hd__and2_2
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ _19747_/Q _16404_/B vssd1 vssd1 vccd1 vccd1 _16410_/C sky130_fd_sc_hd__and2_2
X_13616_ _13626_/A1 _13388_/A _13426_/C _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13616_/X
+ sky130_fd_sc_hd__a22o_2
X_10828_ _10819_/X _10821_/X _10827_/X _10831_/S _12311_/A1 vssd1 vssd1 vccd1 vccd1
+ _10828_/X sky130_fd_sc_hd__o221a_1
X_17384_ _20240_/Q _17390_/A2 _17530_/A2 _20289_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17384_/X sky130_fd_sc_hd__a221o_1
XFILLER_198_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14596_ _19362_/Q _17112_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19362_/D sky130_fd_sc_hd__mux2_1
X_19123_ _19223_/CLK _19123_/D vssd1 vssd1 vccd1 vccd1 _19123_/Q sky130_fd_sc_hd__dfxtp_1
X_16335_ _19721_/Q _16338_/C _18863_/A vssd1 vssd1 vccd1 vccd1 _16335_/Y sky130_fd_sc_hd__a21oi_1
X_13547_ _13575_/C _13559_/B _13545_/X _13546_/X vssd1 vssd1 vccd1 vccd1 _13547_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ _11094_/S _10758_/X _10757_/X _12398_/C1 vssd1 vssd1 vccd1 vccd1 _10759_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_158_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19054_ _20399_/Q vssd1 vssd1 vccd1 vccd1 _20399_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_187_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16266_ _19682_/Q _17800_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19682_/D sky130_fd_sc_hd__mux2_1
XFILLER_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13478_ _13478_/A _13478_/B vssd1 vssd1 vccd1 vccd1 _13478_/X sky130_fd_sc_hd__and2_2
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18005_ _20740_/Q _18005_/B vssd1 vssd1 vccd1 vccd1 _18011_/C sky130_fd_sc_hd__and2_4
XFILLER_161_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15217_ _15610_/A1 _15212_/X _15216_/X vssd1 vssd1 vccd1 vccd1 _15218_/B sky130_fd_sc_hd__a21oi_4
X_12429_ _12429_/A1 _12428_/X _12427_/X vssd1 vssd1 vccd1 vccd1 _12429_/X sky130_fd_sc_hd__o21a_1
XFILLER_195_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16197_ _16197_/A _16197_/B vssd1 vssd1 vccd1 vccd1 _19622_/D sky130_fd_sc_hd__and2_1
XFILLER_173_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput305 _13478_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[0] sky130_fd_sc_hd__buf_4
XFILLER_142_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput316 _13479_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[1] sky130_fd_sc_hd__buf_4
Xoutput327 _13525_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[4] sky130_fd_sc_hd__buf_4
X_15148_ _15282_/A _16743_/B _15129_/X vssd1 vssd1 vccd1 vccd1 _15148_/Y sky130_fd_sc_hd__o21ai_2
Xoutput338 _13692_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[13] sky130_fd_sc_hd__buf_4
XFILLER_141_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput349 _13738_/X vssd1 vssd1 vccd1 vccd1 core_wb_data_o[23] sky130_fd_sc_hd__buf_4
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15079_ _19703_/Q _15595_/A2 _15595_/B1 _19735_/Q vssd1 vssd1 vccd1 vccd1 _15079_/X
+ sky130_fd_sc_hd__a22o_1
X_19956_ _19956_/CLK _19956_/D vssd1 vssd1 vccd1 vccd1 _19956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18907_ _18975_/A _18907_/B vssd1 vssd1 vccd1 vccd1 _18907_/Y sky130_fd_sc_hd__nand2_2
X_19887_ _20451_/CLK _19887_/D vssd1 vssd1 vccd1 vccd1 _19887_/Q sky130_fd_sc_hd__dfxtp_1
X_09640_ _11234_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _09640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18838_ _19128_/Q _12533_/B _18949_/B1 vssd1 vssd1 vccd1 vccd1 _18838_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_109_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20860_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ _12577_/A _13653_/A vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__nor2_8
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18769_ _18320_/A _18457_/B _18457_/C _18570_/B vssd1 vssd1 vccd1 vccd1 _18769_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_255_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20800_ _20863_/CLK _20800_/D vssd1 vssd1 vccd1 vccd1 _20800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20731_ _20795_/CLK _20731_/D vssd1 vssd1 vccd1 vccd1 _20731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20662_ _20662_/CLK _20662_/D vssd1 vssd1 vccd1 vccd1 _20662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20593_ _20667_/CLK _20593_/D vssd1 vssd1 vccd1 vccd1 _20593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout510 _17745_/X vssd1 vssd1 vccd1 vccd1 _17777_/S sky130_fd_sc_hd__buf_12
XFILLER_160_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1508 fanout1534/X vssd1 vssd1 vccd1 vccd1 _11818_/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout1519 fanout1522/X vssd1 vssd1 vccd1 vccd1 _12148_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_99_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout521 _17642_/X vssd1 vssd1 vccd1 vccd1 _17669_/S sky130_fd_sc_hd__buf_6
Xfanout532 _17540_/X vssd1 vssd1 vccd1 vccd1 _17569_/S sky130_fd_sc_hd__clkbuf_16
X_09907_ _11423_/C1 _16063_/B2 _09906_/X vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__a21oi_2
Xfanout543 _17151_/X vssd1 vssd1 vccd1 vccd1 _17178_/S sky130_fd_sc_hd__buf_12
Xfanout554 _17049_/X vssd1 vssd1 vccd1 vccd1 _17081_/S sky130_fd_sc_hd__buf_12
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout565 _16605_/X vssd1 vssd1 vccd1 vccd1 _16632_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_259_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20027_ _20085_/CLK _20027_/D vssd1 vssd1 vccd1 vccd1 _20027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout576 _16272_/S vssd1 vssd1 vccd1 vccd1 _16274_/S sky130_fd_sc_hd__buf_8
Xfanout587 _14738_/Y vssd1 vssd1 vccd1 vccd1 _14802_/A2 sky130_fd_sc_hd__clkbuf_8
X_09838_ _09832_/X _09837_/X _12088_/S vssd1 vssd1 vccd1 vccd1 _09839_/B sky130_fd_sc_hd__mux2_1
XFILLER_274_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout598 _14670_/X vssd1 vssd1 vccd1 vccd1 _14685_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09769_ _09776_/S _09764_/Y _09768_/Y _12020_/C1 vssd1 vssd1 vccd1 vccd1 _09769_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_246_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _13413_/A _13414_/A _13415_/A _13416_/A vssd1 vssd1 vccd1 vccd1 _11800_/X
+ sky130_fd_sc_hd__or4_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _13586_/A _12790_/B vssd1 vssd1 vccd1 vccd1 _13571_/B sky130_fd_sc_hd__nor2_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11731_ _13420_/A _13421_/A _13418_/A _13419_/A vssd1 vssd1 vccd1 vccd1 _11731_/X
+ sky130_fd_sc_hd__or4_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ _21025_/CLK _20929_/D vssd1 vssd1 vccd1 vccd1 _20929_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_159_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _18700_/A _14450_/B vssd1 vssd1 vccd1 vccd1 _19249_/D sky130_fd_sc_hd__and2_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _19883_/Q _19784_/Q _11994_/S vssd1 vssd1 vccd1 vccd1 _11662_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ _12726_/C _13377_/Y _12715_/Y vssd1 vssd1 vccd1 vccd1 _13401_/Y sky130_fd_sc_hd__o21ai_1
X_10613_ _12711_/A _20502_/Q _10628_/S _20534_/Q vssd1 vssd1 vccd1 vccd1 _10613_/X
+ sky130_fd_sc_hd__o22a_1
X_14381_ _20292_/Q _14431_/A2 _14431_/B1 input233/X vssd1 vssd1 vccd1 vccd1 _14383_/B
+ sky130_fd_sc_hd__a22o_2
X_11593_ _11591_/X _11592_/X _12135_/A vssd1 vssd1 vccd1 vccd1 _11593_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ _10556_/X _16132_/A2 _16119_/X vssd1 vssd1 vccd1 vccd1 _19584_/D sky130_fd_sc_hd__o21a_1
X_10544_ _19568_/Q _11240_/S vssd1 vssd1 vccd1 vccd1 _10544_/X sky130_fd_sc_hd__or2_1
XFILLER_183_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13332_ _13332_/A _13332_/B _13347_/A vssd1 vssd1 vccd1 vccd1 _13334_/B sky130_fd_sc_hd__and3_1
XFILLER_182_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16051_ _16051_/A1 _16037_/Y _16051_/B1 vssd1 vssd1 vccd1 vccd1 _16051_/Y sky130_fd_sc_hd__o21ai_1
X_10475_ _19537_/Q _09596_/B _12245_/A1 _10473_/Y vssd1 vssd1 vccd1 vccd1 _13675_/B
+ sky130_fd_sc_hd__a211o_4
X_13263_ _13205_/A _19238_/Q _18752_/A _13262_/Y vssd1 vssd1 vccd1 vccd1 _13412_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15002_ _15322_/B _15000_/X _15001_/Y _14999_/X vssd1 vssd1 vccd1 vccd1 _15002_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12214_ _19427_/Q _12375_/S vssd1 vssd1 vccd1 vccd1 _12214_/X sky130_fd_sc_hd__or2_1
X_13194_ _13017_/Y _13194_/B vssd1 vssd1 vccd1 vccd1 _13195_/B sky130_fd_sc_hd__nand2b_1
XFILLER_68_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12145_ _19651_/Q _12146_/S _12131_/X _12150_/S vssd1 vssd1 vccd1 vccd1 _12145_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20081_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19810_ _20472_/CLK _19810_/D vssd1 vssd1 vccd1 vccd1 _19810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19741_ _20757_/CLK _19741_/D vssd1 vssd1 vccd1 vccd1 _19741_/Q sky130_fd_sc_hd__dfxtp_1
X_16953_ _16949_/Y _16952_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16953_/Y sky130_fd_sc_hd__a21oi_4
X_12076_ _12403_/A1 _12075_/Y _12403_/B1 vssd1 vssd1 vccd1 vccd1 _12076_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_111_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11027_ _19369_/Q _11291_/A2 _11025_/X _11291_/B2 _11026_/X vssd1 vssd1 vccd1 vccd1
+ _11027_/X sky130_fd_sc_hd__o221a_1
X_15904_ _15904_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15904_/Y sky130_fd_sc_hd__nand2_1
X_19672_ _20703_/CLK _19672_/D vssd1 vssd1 vccd1 vccd1 _19672_/Q sky130_fd_sc_hd__dfxtp_1
X_16884_ input50/X input85/X _16884_/S vssd1 vssd1 vccd1 vccd1 _16885_/B sky130_fd_sc_hd__mux2_8
XFILLER_65_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_202_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20075_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_264_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18623_ _20929_/Q _18686_/B vssd1 vssd1 vccd1 vccd1 _18623_/Y sky130_fd_sc_hd__nand2_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _15973_/A1 _15834_/X _15822_/X vssd1 vssd1 vccd1 vccd1 _15835_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_280_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18554_ _20911_/Q fanout750/X _18553_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18555_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _16053_/A _15438_/Y _15765_/X vssd1 vssd1 vccd1 vccd1 _15766_/X sky130_fd_sc_hd__o21ba_1
X_12978_ _12978_/A _12978_/B _12975_/X vssd1 vssd1 vccd1 vccd1 _12979_/A sky130_fd_sc_hd__or3b_1
XFILLER_45_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17505_/A1 _17504_/Y _18932_/A vssd1 vssd1 vccd1 vccd1 _20287_/D sky130_fd_sc_hd__a21oi_1
XFILLER_75_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14717_ _19474_/Q _17689_/A1 _14733_/S vssd1 vssd1 vccd1 vccd1 _19474_/D sky130_fd_sc_hd__mux2_1
X_18485_ _18783_/A _18485_/B vssd1 vssd1 vccd1 vccd1 _20888_/D sky130_fd_sc_hd__nor2_1
X_11929_ _12003_/A _20518_/Q _11932_/S0 _20550_/Q vssd1 vssd1 vccd1 vccd1 _11929_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_221_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15697_ _19752_/Q _15999_/A2 _15696_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15697_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_470 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_481 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_492 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17436_ _17446_/A _17451_/A vssd1 vssd1 vccd1 vccd1 _17457_/C sky130_fd_sc_hd__nor2_1
XFILLER_220_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14648_ _19410_/Q _17932_/A1 _14650_/S vssd1 vssd1 vccd1 vccd1 _19410_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_17 _16833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_28 _15807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_39 _16739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17367_ _20232_/Q _17371_/A2 _17366_/X _18718_/A vssd1 vssd1 vccd1 vccd1 _20232_/D
+ sky130_fd_sc_hd__o211a_1
X_14579_ _19345_/Q _17931_/A1 _14594_/S vssd1 vssd1 vccd1 vccd1 _19345_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19106_ _20721_/CLK _19106_/D vssd1 vssd1 vccd1 vccd1 _19106_/Q sky130_fd_sc_hd__dfxtp_4
X_16318_ _16322_/C _16318_/B vssd1 vssd1 vccd1 vccd1 _19714_/D sky130_fd_sc_hd__nor2_1
XFILLER_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17298_ _20205_/Q _17328_/A2 _17296_/X _17297_/X _17974_/B1 vssd1 vssd1 vccd1 vccd1
+ _20205_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19037_ _21037_/Q _19049_/A2 _19036_/X _18748_/A vssd1 vssd1 vccd1 vccd1 _21037_/D
+ sky130_fd_sc_hd__o211a_1
X_16249_ _19665_/Q _17923_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19665_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19939_ _20667_/CLK _19939_/D vssd1 vssd1 vccd1 vccd1 _19939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09623_ _17709_/C _09623_/B vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__xnor2_1
XFILLER_256_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09554_ _12510_/A _19156_/Q _09555_/C _09567_/A vssd1 vssd1 vccd1 vccd1 _16066_/A
+ sky130_fd_sc_hd__nor4_4
XFILLER_270_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09485_ _17423_/D vssd1 vssd1 vccd1 vccd1 _17451_/A sky130_fd_sc_hd__inv_2
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20714_ _20714_/CLK _20714_/D vssd1 vssd1 vccd1 vccd1 _20714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_77_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20670_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_168_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20645_ _20645_/CLK _20645_/D vssd1 vssd1 vccd1 vccd1 _20645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20576_ _20716_/CLK _20576_/D vssd1 vssd1 vccd1 vccd1 _20576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _10251_/X _10259_/X _10260_/S vssd1 vssd1 vccd1 vccd1 _10260_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout2006 _13466_/A vssd1 vssd1 vccd1 vccd1 _16875_/B2 sky130_fd_sc_hd__buf_4
XFILLER_79_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10191_ _10189_/X _10190_/X _11033_/S vssd1 vssd1 vccd1 vccd1 _10191_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1305 _13466_/X vssd1 vssd1 vccd1 vccd1 _13468_/B sky130_fd_sc_hd__buf_6
XFILLER_160_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1316 _12470_/Y vssd1 vssd1 vccd1 vccd1 _15264_/B sky130_fd_sc_hd__buf_6
XFILLER_278_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1327 _12459_/Y vssd1 vssd1 vccd1 vccd1 _15365_/A sky130_fd_sc_hd__buf_8
Xfanout1338 _09738_/Y vssd1 vssd1 vccd1 vccd1 _11192_/A2 sky130_fd_sc_hd__buf_8
XFILLER_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1349 _17230_/Y vssd1 vssd1 vccd1 vccd1 _17364_/A2 sky130_fd_sc_hd__buf_6
XFILLER_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13950_ _19150_/Q _13953_/A2 _14004_/B1 _13949_/X _16197_/A vssd1 vssd1 vccd1 vccd1
+ _19150_/D sky130_fd_sc_hd__o221a_1
XFILLER_143_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12901_ _19522_/Q _12901_/B vssd1 vssd1 vccd1 vccd1 _12902_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13881_ _19099_/Q _13953_/A2 _13881_/B1 _19165_/Q _15288_/C1 vssd1 vssd1 vccd1 vccd1
+ _19099_/D sky130_fd_sc_hd__o221a_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _16005_/A1 _12703_/X _15619_/Y vssd1 vssd1 vccd1 vccd1 _15620_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12832_ _19168_/Q _12832_/B vssd1 vssd1 vccd1 vccd1 _12839_/B sky130_fd_sc_hd__nor2_2
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15551_/A _16028_/C vssd1 vssd1 vccd1 vccd1 _15551_/X sky130_fd_sc_hd__and2_1
XFILLER_188_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12763_ _14803_/A1 _12582_/C _12784_/B _12762_/Y vssd1 vssd1 vccd1 vccd1 _12763_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_261_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _19280_/Q _17899_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19280_/D sky130_fd_sc_hd__mux2_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18270_ _18532_/B vssd1 vssd1 vccd1 vccd1 _18270_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _09834_/C _11713_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _11714_/X sky130_fd_sc_hd__a21o_1
X_15482_ _17305_/A _15482_/A2 _15476_/X _15606_/A1 vssd1 vssd1 vccd1 vccd1 _15482_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12694_ _13526_/B _13526_/C _12693_/Y vssd1 vssd1 vccd1 vccd1 _13544_/A sky130_fd_sc_hd__a21o_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _14139_/B _17219_/Y _17220_/X _18698_/A vssd1 vssd1 vccd1 vccd1 _20182_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14433_/A _14433_/B vssd1 vssd1 vccd1 vccd1 _14433_/Y sky130_fd_sc_hd__nor2_1
XFILLER_230_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11645_ _12192_/A1 _11634_/X _11638_/X _11644_/X vssd1 vssd1 vccd1 vccd1 _11646_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17152_ _20118_/Q _17780_/A1 _17166_/S vssd1 vssd1 vccd1 vccd1 _20118_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14364_ _19518_/Q _14364_/B vssd1 vssd1 vccd1 vccd1 _14365_/B sky130_fd_sc_hd__nand2_1
Xinput15 core_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_4
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ _20480_/Q _20320_/Q _11599_/S vssd1 vssd1 vccd1 vccd1 _11576_/X sky130_fd_sc_hd__mux2_1
Xinput26 core_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_4
XFILLER_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput37 core_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_4
X_16103_ _19576_/Q _16127_/A2 _16107_/B1 vssd1 vssd1 vccd1 vccd1 _16103_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 dout0[14] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
Xinput59 dout0[24] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_2
X_13315_ _13039_/Y _13315_/B vssd1 vssd1 vccd1 vccd1 _13316_/B sky130_fd_sc_hd__nand2b_1
X_17083_ _17851_/A _17851_/B _17083_/C vssd1 vssd1 vccd1 vccd1 _17083_/X sky130_fd_sc_hd__and3_4
X_10527_ _11290_/A _19312_/Q _11290_/C vssd1 vssd1 vccd1 vccd1 _10527_/X sky130_fd_sc_hd__or3_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14295_ _14325_/A _14293_/Y _14294_/X _14295_/C1 vssd1 vssd1 vccd1 vccd1 _14295_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16034_ _13181_/A _16033_/X _16034_/S vssd1 vssd1 vccd1 vccd1 _16034_/X sky130_fd_sc_hd__mux2_1
X_10458_ input108/X input143/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__mux2_8
X_13246_ _13346_/A _13346_/B _13346_/C vssd1 vssd1 vccd1 vccd1 _13347_/A sky130_fd_sc_hd__a21o_1
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10389_ _09829_/A _19473_/Q _19441_/Q _10400_/S vssd1 vssd1 vccd1 vccd1 _10389_/X
+ sky130_fd_sc_hd__a22o_1
X_13177_ _12281_/Y _13182_/B _12283_/B vssd1 vssd1 vccd1 vccd1 _13178_/B sky130_fd_sc_hd__a21oi_4
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12128_ _12126_/X _12127_/X _12134_/S vssd1 vssd1 vccd1 vccd1 _12128_/X sky130_fd_sc_hd__mux2_1
X_17985_ _20733_/Q _20732_/Q _17985_/C vssd1 vssd1 vccd1 vccd1 _17991_/C sky130_fd_sc_hd__and3_1
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1850 _13192_/A vssd1 vssd1 vccd1 vccd1 _11268_/A sky130_fd_sc_hd__buf_8
X_16936_ _19983_/Q _17012_/A2 _16935_/Y _18094_/A vssd1 vssd1 vccd1 vccd1 _19983_/D
+ sky130_fd_sc_hd__a211o_1
X_12059_ _12059_/A1 _12058_/X _12055_/X _12059_/C1 vssd1 vssd1 vccd1 vccd1 _12059_/X
+ sky130_fd_sc_hd__a211o_2
X_19724_ _19759_/CLK _19724_/D vssd1 vssd1 vccd1 vccd1 _19724_/Q sky130_fd_sc_hd__dfxtp_2
Xfanout1861 _19169_/Q vssd1 vssd1 vccd1 vccd1 _18765_/B sky130_fd_sc_hd__buf_12
XFILLER_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1872 _12504_/B vssd1 vssd1 vccd1 vccd1 _09507_/A sky130_fd_sc_hd__buf_8
XFILLER_42_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1883 _14112_/A vssd1 vssd1 vccd1 vccd1 _09609_/A sky130_fd_sc_hd__buf_6
XFILLER_38_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1894 fanout1905/X vssd1 vssd1 vccd1 vccd1 _18752_/A sky130_fd_sc_hd__buf_6
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_281_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16867_ _16887_/A _16867_/B vssd1 vssd1 vccd1 vccd1 _16867_/Y sky130_fd_sc_hd__nor2_1
X_19655_ _20410_/CLK _19655_/D vssd1 vssd1 vccd1 vccd1 _19655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18606_ _18842_/A _18606_/B vssd1 vssd1 vccd1 vccd1 _20924_/D sky130_fd_sc_hd__nor2_1
X_15818_ _09784_/B _15984_/A2 _15984_/B1 _09782_/A _15890_/A vssd1 vssd1 vccd1 vccd1
+ _15818_/X sky130_fd_sc_hd__a221o_1
XFILLER_281_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19586_ _20665_/CLK _19586_/D vssd1 vssd1 vccd1 vccd1 _19586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16798_ _16718_/X _16797_/X _13468_/B vssd1 vssd1 vccd1 vccd1 _16798_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_213_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18537_ _18932_/A _18537_/B vssd1 vssd1 vccd1 vccd1 _20905_/D sky130_fd_sc_hd__nor2_1
XFILLER_240_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15749_ _20966_/Q _16045_/A2 _16016_/S _20838_/Q _15748_/X vssd1 vssd1 vccd1 vccd1
+ _15749_/X sky130_fd_sc_hd__a221o_1
XFILLER_178_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18468_ _18589_/B _12557_/Y _12592_/C _18474_/S _20884_/Q vssd1 vssd1 vccd1 vccd1
+ _18468_/X sky130_fd_sc_hd__a32o_1
XFILLER_178_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17419_ _17420_/A _20256_/Q _17432_/A _17418_/Y vssd1 vssd1 vccd1 vccd1 _20255_/D
+ sky130_fd_sc_hd__o211a_1
X_18399_ _20854_/Q _18180_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18400_/B sky130_fd_sc_hd__mux2_1
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20430_ _20561_/CLK _20430_/D vssd1 vssd1 vccd1 vccd1 _20430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20361_ _20685_/CLK _20361_/D vssd1 vssd1 vccd1 vccd1 _20361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20292_ _20296_/CLK _20292_/D vssd1 vssd1 vccd1 vccd1 _20292_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_195_wb_clk_i _20408_/CLK vssd1 vssd1 vccd1 vccd1 _20706_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20268_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09606_ _09606_/A _09606_/B vssd1 vssd1 vccd1 vccd1 _12975_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09537_ _19151_/Q _19150_/Q vssd1 vssd1 vccd1 vccd1 _12490_/B sky130_fd_sc_hd__nand2_4
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11430_ _20135_/Q _20103_/Q _12133_/S vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__mux2_1
X_20628_ _20660_/CLK _20628_/D vssd1 vssd1 vccd1 vccd1 _20628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11361_ _19275_/Q _20062_/Q _12300_/S vssd1 vssd1 vccd1 vccd1 _11361_/X sky130_fd_sc_hd__mux2_1
X_20559_ _20559_/CLK _20559_/D vssd1 vssd1 vccd1 vccd1 _20559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10312_ _20539_/Q _10324_/S vssd1 vssd1 vccd1 vccd1 _10312_/X sky130_fd_sc_hd__or2_1
X_13100_ _13100_/A _13100_/B vssd1 vssd1 vccd1 vccd1 _13100_/X sky130_fd_sc_hd__and2_1
X_14080_ _19199_/Q _14104_/A2 _14079_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1 _19199_/D
+ sky130_fd_sc_hd__o211a_1
X_11292_ _20397_/Q _20333_/Q _20625_/Q _20589_/Q _11292_/S0 _11026_/C vssd1 vssd1
+ vccd1 vccd1 _11292_/X sky130_fd_sc_hd__mux4_1
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13031_ _20962_/Q _20896_/Q vssd1 vssd1 vccd1 vccd1 _13031_/Y sky130_fd_sc_hd__nor2_1
X_10243_ _12403_/A1 _13698_/A _12403_/B1 vssd1 vssd1 vccd1 vccd1 _10243_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_267_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10174_ _19878_/Q _19779_/Q _10174_/S vssd1 vssd1 vccd1 vccd1 _10174_/X sky130_fd_sc_hd__mux2_1
Xfanout1102 _17878_/A1 vssd1 vssd1 vccd1 vccd1 _17178_/A1 sky130_fd_sc_hd__buf_4
Xfanout1113 _11807_/X vssd1 vssd1 vccd1 vccd1 _17944_/A1 sky130_fd_sc_hd__buf_2
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1124 _17902_/A1 vssd1 vssd1 vccd1 vccd1 _17202_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1135 _10681_/X vssd1 vssd1 vccd1 vccd1 _17893_/A1 sky130_fd_sc_hd__buf_8
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17770_ _20549_/Q _17910_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20549_/D sky130_fd_sc_hd__mux2_1
Xfanout1146 _17908_/A1 vssd1 vssd1 vccd1 vccd1 _17942_/A1 sky130_fd_sc_hd__buf_2
X_14982_ _15022_/A _15022_/B _15022_/C vssd1 vssd1 vccd1 vccd1 _14987_/B sky130_fd_sc_hd__or3_4
Xfanout1157 _09631_/X vssd1 vssd1 vccd1 vccd1 _12153_/A1 sky130_fd_sc_hd__buf_8
Xfanout1168 _14898_/Y vssd1 vssd1 vccd1 vccd1 _16050_/A1 sky130_fd_sc_hd__buf_4
XFILLER_248_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1179 _12516_/Y vssd1 vssd1 vccd1 vccd1 _13350_/B sky130_fd_sc_hd__buf_4
XFILLER_219_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16721_ _20397_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16721_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13933_ _19137_/Q _13941_/B _13946_/B1 _13388_/C vssd1 vssd1 vccd1 vccd1 _19137_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19440_ _21047_/A _19440_/D vssd1 vssd1 vccd1 vccd1 _19440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16652_ _19909_/Q _17096_/A1 _16666_/S vssd1 vssd1 vccd1 vccd1 _19909_/D sky130_fd_sc_hd__mux2_1
X_13864_ _19084_/Q _13953_/A2 _13881_/B1 _19150_/Q _16197_/A vssd1 vssd1 vccd1 vccd1
+ _19084_/D sky130_fd_sc_hd__o221a_1
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15603_ _20801_/Q _15016_/A _15601_/X _15602_/X vssd1 vssd1 vccd1 vccd1 _15603_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_223_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19371_ _20662_/CLK _19371_/D vssd1 vssd1 vccd1 vccd1 _19371_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ _12906_/A _12815_/B vssd1 vssd1 vccd1 vccd1 _13362_/A sky130_fd_sc_hd__xnor2_4
XFILLER_90_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16583_ _16591_/A _16583_/B vssd1 vssd1 vccd1 vccd1 _19857_/D sky130_fd_sc_hd__or2_1
XFILLER_222_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13795_ _13798_/A1 _13802_/A1 _13685_/B _13805_/B1 input241/X vssd1 vssd1 vccd1 vccd1
+ _13795_/X sky130_fd_sc_hd__a32o_1
XFILLER_43_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18322_ _18322_/A _18323_/B _18322_/C _18138_/B vssd1 vssd1 vccd1 vccd1 _18563_/C
+ sky130_fd_sc_hd__or4b_2
XFILLER_16_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _20927_/Q _15567_/A2 _15533_/X vssd1 vssd1 vccd1 vccd1 _15534_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12746_ _12747_/A _12747_/B _12747_/C vssd1 vssd1 vccd1 vccd1 _12749_/C sky130_fd_sc_hd__a21oi_4
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18253_ _19546_/Q _18313_/B vssd1 vssd1 vccd1 vccd1 _18253_/Y sky130_fd_sc_hd__nand2b_2
X_15465_ _15465_/A _15465_/B vssd1 vssd1 vccd1 vccd1 _15465_/Y sky130_fd_sc_hd__nand2_1
X_12677_ _12675_/B _12675_/C _13501_/A _12676_/A vssd1 vssd1 vccd1 vccd1 _12678_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17204_ _20168_/Q _17695_/A1 _17212_/S vssd1 vssd1 vccd1 vccd1 _20168_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14416_ _14416_/A _14424_/B vssd1 vssd1 vccd1 vccd1 _14416_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18184_ _18213_/B _14171_/B _18183_/Y vssd1 vssd1 vccd1 vccd1 _18480_/B sky130_fd_sc_hd__o21ai_4
X_11628_ _12191_/C1 _11933_/S _11627_/X _10409_/A vssd1 vssd1 vccd1 vccd1 _11628_/X
+ sky130_fd_sc_hd__a31o_1
X_15396_ _15396_/A1 _15381_/X _15395_/X vssd1 vssd1 vccd1 vccd1 _16804_/B sky130_fd_sc_hd__a21oi_4
XFILLER_200_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17135_ _20103_/Q _17869_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20103_/D sky130_fd_sc_hd__mux2_1
X_14347_ _13205_/A _14346_/X _13399_/Y vssd1 vssd1 vccd1 vccd1 _14348_/C sky130_fd_sc_hd__o21a_1
XFILLER_171_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ _09986_/C _11558_/X _12006_/S vssd1 vssd1 vccd1 vccd1 _11559_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17066_ _20038_/Q _17693_/A1 _17078_/S vssd1 vssd1 vccd1 vccd1 _20038_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ _14278_/A _14278_/B vssd1 vssd1 vccd1 vccd1 _14283_/A sky130_fd_sc_hd__nor2_2
XFILLER_143_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16017_ _20976_/Q _16045_/A2 _16016_/X _16017_/C1 vssd1 vssd1 vccd1 vccd1 _16017_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13229_ _13373_/A _13229_/B _13229_/C vssd1 vssd1 vccd1 vccd1 _13229_/X sky130_fd_sc_hd__and3_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_6__f_wb_clk_i clkbuf_3_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_6__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17968_ _20727_/Q _17971_/C _18064_/A vssd1 vssd1 vccd1 vccd1 _17968_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_257_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19707_ _20757_/CLK _19707_/D vssd1 vssd1 vccd1 vccd1 _19707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1680 _12007_/A1 vssd1 vssd1 vccd1 vccd1 _12003_/A sky130_fd_sc_hd__buf_4
XFILLER_214_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16919_ _16916_/Y _16918_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16919_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_272_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1691 _10937_/A vssd1 vssd1 vccd1 vccd1 _11026_/A sky130_fd_sc_hd__buf_2
X_17899_ _20670_/Q _17899_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20670_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19638_ _20660_/CLK _19638_/D vssd1 vssd1 vccd1 vccd1 _19638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19569_ _19577_/CLK _19569_/D vssd1 vssd1 vccd1 vccd1 _19569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20413_ _20421_/CLK _20413_/D vssd1 vssd1 vccd1 vccd1 _20413_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_88_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20344_ _20668_/CLK _20344_/D vssd1 vssd1 vccd1 vccd1 _20344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20275_ _21018_/CLK _20275_/D vssd1 vssd1 vccd1 vccd1 _20275_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput205 localMemory_wb_adr_i[23] vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__buf_6
XFILLER_130_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput216 localMemory_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_hd__buf_12
XFILLER_89_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput227 localMemory_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_hd__buf_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput238 localMemory_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_hd__buf_12
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput249 localMemory_wb_sel_i[2] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_hd__clkbuf_2
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10930_ _19161_/Q _12569_/A vssd1 vssd1 vccd1 vccd1 _10930_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_92_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20426_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_245_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10861_ _10859_/X _10860_/X _12414_/S vssd1 vssd1 vccd1 vccd1 _10861_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_wb_clk_i _20408_/CLK vssd1 vssd1 vccd1 vccd1 _20675_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_231_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _19502_/Q _19501_/Q _12639_/A vssd1 vssd1 vccd1 vccd1 _12781_/B sky130_fd_sc_hd__and3_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13573_/Y _13576_/X _13552_/A vssd1 vssd1 vccd1 vccd1 _13580_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10792_ _12357_/A1 _10790_/X _10791_/X vssd1 vssd1 vccd1 vccd1 _10792_/X sky130_fd_sc_hd__o21a_1
XFILLER_231_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _19118_/Q _19117_/Q vssd1 vssd1 vccd1 vccd1 _12531_/Y sky130_fd_sc_hd__nor2_4
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _19531_/Q _15402_/A _15249_/Y _16165_/C1 vssd1 vssd1 vccd1 vccd1 _19531_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ _14895_/A _14898_/A vssd1 vssd1 vccd1 vccd1 _12462_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14201_ _14201_/A _14201_/B vssd1 vssd1 vccd1 vccd1 _14201_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_8_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11413_ _13424_/A _11754_/A _11411_/X vssd1 vssd1 vccd1 vccd1 _11413_/Y sky130_fd_sc_hd__a21oi_2
X_15181_ _14841_/S _15180_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _15181_/X sky130_fd_sc_hd__o21a_1
X_12393_ _19653_/Q _19959_/Q _12397_/S vssd1 vssd1 vccd1 vccd1 _12393_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14132_ _14130_/B _14131_/Y _14202_/S vssd1 vssd1 vccd1 vccd1 _14132_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11344_ _09503_/A _11339_/X _11340_/X vssd1 vssd1 vccd1 vccd1 _11344_/X sky130_fd_sc_hd__o21a_1
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14063_ _14081_/A _14069_/B _14063_/C vssd1 vssd1 vccd1 vccd1 _14063_/X sky130_fd_sc_hd__or3_1
XFILLER_180_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18940_ _19110_/Q _18954_/A2 _18967_/B1 _15898_/A vssd1 vssd1 vccd1 vccd1 _18941_/B
+ sky130_fd_sc_hd__a22o_1
X_11275_ _11275_/A _11275_/B _11275_/C vssd1 vssd1 vccd1 vccd1 _11275_/X sky130_fd_sc_hd__or3_1
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ _20972_/Q _20906_/Q vssd1 vssd1 vccd1 vccd1 _13086_/B sky130_fd_sc_hd__nor2_1
X_10226_ _11008_/A1 _20508_/Q _10235_/S _10225_/X vssd1 vssd1 vccd1 vccd1 _10226_/X
+ sky130_fd_sc_hd__o211a_1
X_18871_ _19100_/Q _18974_/A2 _18974_/B1 _13427_/C vssd1 vssd1 vccd1 vccd1 _18872_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17822_ _20597_/Q _17894_/A1 _17844_/S vssd1 vssd1 vccd1 vccd1 _20597_/D sky130_fd_sc_hd__mux2_1
X_10157_ _12230_/A1 _19910_/Q _11359_/S _10145_/X vssd1 vssd1 vccd1 vccd1 _10157_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_255_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17753_ _20532_/Q _17893_/A1 _17776_/S vssd1 vssd1 vccd1 vccd1 _20532_/D sky130_fd_sc_hd__mux2_1
X_14965_ _15019_/B _15019_/C _15308_/C vssd1 vssd1 vccd1 vccd1 _14965_/X sky130_fd_sc_hd__and3_1
X_10088_ _10356_/A _19346_/Q _20701_/Q _10518_/S _11304_/S vssd1 vssd1 vccd1 vccd1
+ _10088_/X sky130_fd_sc_hd__a221o_1
XFILLER_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16704_ _19959_/Q _17114_/A1 _16704_/S vssd1 vssd1 vccd1 vccd1 _19959_/D sky130_fd_sc_hd__mux2_1
X_13916_ _19123_/Q _13919_/S _13915_/Y _18710_/A vssd1 vssd1 vccd1 vccd1 _19123_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17684_ _20468_/Q _17684_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20468_/D sky130_fd_sc_hd__mux2_1
X_14896_ _11305_/B _11312_/X _15528_/B vssd1 vssd1 vccd1 vccd1 _14896_/X sky130_fd_sc_hd__mux2_1
XFILLER_262_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16635_ _19894_/Q _17706_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19894_/D sky130_fd_sc_hd__mux2_1
X_19423_ _20714_/CLK _19423_/D vssd1 vssd1 vccd1 vccd1 _19423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _20217_/Q _13844_/B _13844_/X vssd1 vssd1 vccd1 vccd1 _13847_/X sky130_fd_sc_hd__a21bo_1
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16566_ _19849_/Q _16566_/A2 _16566_/B1 input19/X vssd1 vssd1 vccd1 vccd1 _16567_/B
+ sky130_fd_sc_hd__o22a_1
X_19354_ _20713_/CLK _19354_/D vssd1 vssd1 vccd1 vccd1 _19354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13778_ _13698_/X _13741_/B _13741_/Y _13699_/Y _13777_/X vssd1 vssd1 vccd1 vccd1
+ _13779_/B sky130_fd_sc_hd__o221a_4
XFILLER_210_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15517_ _16049_/A1 _15506_/X _15516_/X vssd1 vssd1 vccd1 vccd1 _16842_/B sky130_fd_sc_hd__a21oi_4
X_18305_ _18553_/B vssd1 vssd1 vccd1 vccd1 _18305_/Y sky130_fd_sc_hd__clkinv_4
X_19285_ _20081_/CLK _19285_/D vssd1 vssd1 vccd1 vccd1 _19285_/Q sky130_fd_sc_hd__dfxtp_1
X_12729_ _12740_/B _12729_/B vssd1 vssd1 vccd1 vccd1 _12729_/X sky130_fd_sc_hd__or2_1
X_16497_ _19804_/Q _17649_/A1 _16521_/S vssd1 vssd1 vccd1 vccd1 _19804_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18236_ _20801_/Q _18235_/Y _18236_/S vssd1 vssd1 vccd1 vccd1 _18237_/B sky130_fd_sc_hd__mux2_1
X_15448_ _20924_/Q _15567_/A2 _15447_/X vssd1 vssd1 vccd1 vccd1 _15448_/X sky130_fd_sc_hd__o21a_1
X_18167_ _18414_/A _18167_/B vssd1 vssd1 vccd1 vccd1 _20787_/D sky130_fd_sc_hd__and2_1
XFILLER_157_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15379_ _12578_/B _12773_/X _11398_/S vssd1 vssd1 vccd1 vccd1 _15379_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17118_ _20086_/Q _17780_/A1 _17132_/S vssd1 vssd1 vccd1 vccd1 _20086_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18098_ _20774_/Q _18101_/C _18104_/A vssd1 vssd1 vccd1 vccd1 _18098_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_172_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17049_ _17851_/A _17851_/B _17049_/C vssd1 vssd1 vccd1 vccd1 _17049_/X sky130_fd_sc_hd__and3_4
X_09940_ _09941_/B vssd1 vssd1 vccd1 vccd1 _09940_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20060_ _20467_/CLK _20060_/D vssd1 vssd1 vccd1 vccd1 _20060_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout906 _15018_/X vssd1 vssd1 vccd1 vccd1 _15322_/C sky130_fd_sc_hd__buf_6
Xfanout917 _14946_/Y vssd1 vssd1 vccd1 vccd1 _15934_/B1 sky130_fd_sc_hd__buf_12
X_09871_ _20354_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _09871_/X sky130_fd_sc_hd__or2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 _14933_/Y vssd1 vssd1 vccd1 vccd1 _15989_/A2 sky130_fd_sc_hd__clkbuf_4
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 _15292_/S vssd1 vssd1 vccd1 vccd1 _15357_/S sky130_fd_sc_hd__buf_4
XFILLER_258_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ _20962_/CLK _20962_/D vssd1 vssd1 vccd1 vccd1 _20962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20893_ _20959_/CLK _20893_/D vssd1 vssd1 vccd1 vccd1 _20893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20327_ _20579_/CLK _20327_/D vssd1 vssd1 vccd1 vccd1 _20327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11060_ _11239_/A1 _13960_/A2 _11059_/X _11239_/B1 _19833_/Q vssd1 vssd1 vccd1 vccd1
+ _16073_/A sky130_fd_sc_hd__o32ai_4
XFILLER_89_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20258_ _20261_/CLK _20258_/D vssd1 vssd1 vccd1 vccd1 _20258_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_277_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ _12020_/C1 _10010_/X _11872_/A vssd1 vssd1 vccd1 vccd1 _10011_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20189_ _20428_/CLK _20189_/D vssd1 vssd1 vccd1 vccd1 _20189_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _19122_/Q _14764_/A2 _14749_/X _14758_/C1 vssd1 vssd1 vccd1 vccd1 _19499_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11962_ _19554_/Q _12155_/A2 _12155_/B1 _19618_/Q vssd1 vssd1 vccd1 vccd1 _11962_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13701_ _13702_/B vssd1 vssd1 vccd1 vccd1 _13701_/Y sky130_fd_sc_hd__inv_2
X_10913_ _09618_/A _12371_/A1 _19338_/Q _12302_/S vssd1 vssd1 vccd1 vccd1 _10913_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_205_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _19440_/Q _17930_/A1 _14685_/S vssd1 vssd1 vccd1 vccd1 _19440_/D sky130_fd_sc_hd__mux2_1
XFILLER_244_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _11903_/A1 _12120_/A1 _19359_/Q _12129_/S vssd1 vssd1 vccd1 vccd1 _11893_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_233_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16420_ _19753_/Q _16420_/B vssd1 vssd1 vccd1 vccd1 _16426_/C sky130_fd_sc_hd__and2_2
X_13632_ _15954_/A _13189_/B _16233_/B _13478_/B vssd1 vssd1 vccd1 vccd1 _13632_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_72_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10844_ _10842_/X _10843_/X _12324_/S vssd1 vssd1 vccd1 vccd1 _10844_/X sky130_fd_sc_hd__mux2_1
XFILLER_260_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16351_ _19727_/Q _16354_/C _18835_/A vssd1 vssd1 vccd1 vccd1 _16351_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_213_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13563_ _13563_/A _13564_/B _13562_/X vssd1 vssd1 vccd1 vccd1 _13563_/X sky130_fd_sc_hd__or3b_2
XFILLER_12_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10775_ _20403_/Q _20339_/Q _20631_/Q _20595_/Q _12339_/S0 _12337_/C vssd1 vssd1
+ vccd1 vccd1 _10775_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15302_ _11787_/A _15494_/B _15301_/X vssd1 vssd1 vccd1 vccd1 _15326_/C sky130_fd_sc_hd__a21oi_1
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ _12519_/C _13192_/A _12514_/C _12588_/C vssd1 vssd1 vccd1 vccd1 _12515_/C
+ sky130_fd_sc_hd__or4_1
X_19070_ _20415_/Q vssd1 vssd1 vccd1 vccd1 _20415_/D sky130_fd_sc_hd__clkbuf_2
X_16282_ _20623_/Q _17015_/B _19701_/D vssd1 vssd1 vccd1 vccd1 _19698_/D sky130_fd_sc_hd__and3_1
XFILLER_9_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13494_ _13612_/A _13663_/B _15127_/A _13493_/Y _19661_/D vssd1 vssd1 vccd1 vccd1
+ _13494_/X sky130_fd_sc_hd__a32o_4
X_18021_ _20746_/Q _18024_/C vssd1 vssd1 vccd1 vccd1 _18022_/B sky130_fd_sc_hd__and2_1
X_15233_ _21016_/Q _20984_/Q _15309_/S vssd1 vssd1 vccd1 vccd1 _15233_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12445_ _12447_/B _12445_/B vssd1 vssd1 vccd1 vccd1 _12446_/A sky130_fd_sc_hd__nand2b_1
XFILLER_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15164_ _15157_/Y _15163_/A _15611_/S vssd1 vssd1 vccd1 vccd1 _15164_/X sky130_fd_sc_hd__mux2_2
X_12376_ _12374_/X _12375_/X _12376_/S vssd1 vssd1 vccd1 vccd1 _12376_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14115_ _16133_/A _13860_/X _14524_/A1 vssd1 vssd1 vccd1 vccd1 _14115_/Y sky130_fd_sc_hd__a21oi_4
X_11327_ _10465_/A _11243_/X _10032_/Y vssd1 vssd1 vccd1 vccd1 _11327_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19972_ _20751_/CLK _19972_/D vssd1 vssd1 vccd1 vccd1 _19972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15095_ _15220_/A _15095_/B _15096_/B vssd1 vssd1 vccd1 vccd1 _15095_/X sky130_fd_sc_hd__and3_1
XFILLER_125_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14046_ _19182_/Q _14082_/A2 _14045_/X _16087_/B1 vssd1 vssd1 vccd1 vccd1 _19182_/D
+ sky130_fd_sc_hd__o211a_1
X_18923_ _21003_/Q _18971_/B vssd1 vssd1 vccd1 vccd1 _18923_/Y sky130_fd_sc_hd__nand2_1
X_11258_ _11258_/A1 _19462_/Q _19430_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _11258_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10209_ _20380_/Q _20444_/Q _10217_/S vssd1 vssd1 vccd1 vccd1 _10209_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18854_ _20993_/Q _18861_/B vssd1 vssd1 vccd1 vccd1 _18854_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11189_ _19495_/Q _11189_/B vssd1 vssd1 vccd1 vccd1 _11189_/Y sky130_fd_sc_hd__nor2_2
XFILLER_268_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17805_ _20582_/Q _17805_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20582_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18785_ _19087_/Q _18785_/A2 _12592_/C _13496_/Y _18949_/A2 vssd1 vssd1 vccd1 vccd1
+ _18785_/X sky130_fd_sc_hd__a221o_1
X_15997_ _16046_/A1 _15996_/X _15992_/X vssd1 vssd1 vccd1 vccd1 _15997_/X sky130_fd_sc_hd__o21a_4
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14948_ _14948_/A _14983_/A vssd1 vssd1 vccd1 vccd1 _14948_/Y sky130_fd_sc_hd__nor2_8
X_17736_ _20517_/Q _17910_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20517_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14879_ _09556_/X _09562_/X _14897_/A _12575_/Y vssd1 vssd1 vccd1 vccd1 _14881_/B
+ sky130_fd_sc_hd__o31a_1
X_17667_ _20453_/Q _17804_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20453_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19406_ _20565_/CLK _19406_/D vssd1 vssd1 vccd1 vccd1 _19406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16618_ _19877_/Q _17689_/A1 _16632_/S vssd1 vssd1 vccd1 vccd1 _19877_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17598_ _20356_/Q _17909_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20356_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19337_ _20565_/CLK _19337_/D vssd1 vssd1 vccd1 vccd1 _19337_/Q sky130_fd_sc_hd__dfxtp_1
X_16549_ _16567_/A _16549_/B vssd1 vssd1 vccd1 vccd1 _19840_/D sky130_fd_sc_hd__or2_1
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19268_ _20694_/CLK _19268_/D vssd1 vssd1 vccd1 vccd1 _19268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _18223_/B _14239_/B _18218_/Y vssd1 vssd1 vccd1 vccd1 _18502_/B sky130_fd_sc_hd__o21ai_4
X_19199_ _20426_/CLK _19199_/D vssd1 vssd1 vccd1 vccd1 _19199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20112_ _20579_/CLK _20112_/D vssd1 vssd1 vccd1 vccd1 _20112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09923_ _20482_/Q _11616_/B _12015_/A1 vssd1 vssd1 vccd1 vccd1 _09923_/X sky130_fd_sc_hd__a21o_1
Xfanout703 _16576_/A2 vssd1 vssd1 vccd1 vccd1 _16592_/A2 sky130_fd_sc_hd__buf_4
Xfanout714 _16576_/B1 vssd1 vssd1 vccd1 vccd1 _16592_/B1 sky130_fd_sc_hd__buf_4
XFILLER_113_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout725 _13244_/X vssd1 vssd1 vccd1 vccd1 _16240_/A1 sky130_fd_sc_hd__buf_6
XFILLER_259_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20043_ _20645_/CLK _20043_/D vssd1 vssd1 vccd1 vccd1 _20043_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout736 _18982_/X vssd1 vssd1 vccd1 vccd1 _19046_/C1 sky130_fd_sc_hd__buf_6
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout747 _18985_/B vssd1 vssd1 vccd1 vccd1 _19046_/A2 sky130_fd_sc_hd__buf_4
XFILLER_113_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09854_ _09851_/X _09852_/X _09853_/X _12103_/A1 _18765_/B vssd1 vssd1 vccd1 vccd1
+ _09854_/X sky130_fd_sc_hd__a221o_1
XFILLER_213_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout758 _18840_/B vssd1 vssd1 vccd1 vccd1 _18861_/B sky130_fd_sc_hd__buf_4
XFILLER_86_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout769 _18683_/B vssd1 vssd1 vccd1 vccd1 _18651_/B sky130_fd_sc_hd__buf_4
XFILLER_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09785_ _19549_/Q _09613_/A _09613_/B _19613_/Q vssd1 vssd1 vccd1 vccd1 _09785_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_107 _16242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_118 _16237_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _13660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20945_ _21009_/CLK _20945_/D vssd1 vssd1 vccd1 vccd1 _20945_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _21041_/CLK _20876_/D vssd1 vssd1 vccd1 vccd1 _20876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10560_ _10035_/Y _10554_/X _10559_/X _10549_/A _10024_/X vssd1 vssd1 vccd1 vccd1
+ _10561_/B sky130_fd_sc_hd__a32o_2
XFILLER_195_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10491_ _20343_/Q _11270_/A2 _10897_/A3 _11170_/B1 vssd1 vssd1 vccd1 vccd1 _10491_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_108_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12230_ _12230_/A1 _20522_/Q _12317_/S _12212_/X vssd1 vssd1 vccd1 vccd1 _12230_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12161_ _20653_/Q _20617_/Q _12182_/S vssd1 vssd1 vccd1 vccd1 _12161_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11112_ _20399_/Q _20335_/Q _20627_/Q _20591_/Q _12339_/S0 _12254_/C vssd1 vssd1
+ vccd1 vccd1 _11112_/X sky130_fd_sc_hd__mux4_1
XFILLER_162_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12092_ _19424_/Q _20583_/Q _12097_/S vssd1 vssd1 vccd1 vccd1 _12092_/X sky130_fd_sc_hd__mux2_1
XFILLER_268_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ _20153_/Q _11379_/B _11378_/S vssd1 vssd1 vccd1 vccd1 _11043_/X sky130_fd_sc_hd__o21a_1
X_15920_ _15890_/B _15903_/Y _15919_/X _15976_/B2 vssd1 vssd1 vccd1 vccd1 _15920_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15851_ _19726_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15851_/X sky130_fd_sc_hd__or2_1
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _19148_/Q _14802_/A2 _14801_/X _14802_/C1 vssd1 vssd1 vccd1 vccd1 _19525_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18570_ _19495_/Q _18570_/B vssd1 vssd1 vccd1 vccd1 _18570_/Y sky130_fd_sc_hd__nand2_2
X_15782_ _16051_/A1 _15768_/X _16051_/B1 vssd1 vssd1 vccd1 vccd1 _15782_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_224_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12994_ _19237_/Q _13390_/B vssd1 vssd1 vccd1 vccd1 _13255_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ _19490_/Q _17112_/A1 _14733_/S vssd1 vssd1 vccd1 vccd1 _19490_/D sky130_fd_sc_hd__mux2_1
X_17521_ _17525_/A1 _17520_/Y _17430_/A vssd1 vssd1 vccd1 vccd1 _20295_/D sky130_fd_sc_hd__a21oi_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ _11943_/X _11944_/X _11945_/S vssd1 vssd1 vccd1 vccd1 _11945_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_630 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_641 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_652 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17452_ _17452_/A _17456_/B vssd1 vssd1 vccd1 vccd1 _17454_/C sky130_fd_sc_hd__nor2_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14664_ _19426_/Q _17112_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19426_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11876_ _11877_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11878_/A sky130_fd_sc_hd__nor2_2
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _18086_/A _16403_/B _16404_/B vssd1 vssd1 vccd1 vccd1 _19746_/D sky130_fd_sc_hd__nor3_1
XFILLER_221_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ _13626_/A1 _13361_/B _15494_/A _13626_/B2 vssd1 vssd1 vccd1 vccd1 _13615_/X
+ sky130_fd_sc_hd__a22o_2
X_10827_ _10825_/X _10826_/X _11359_/S vssd1 vssd1 vccd1 vccd1 _10827_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17383_ _20240_/Q _17401_/A2 _17382_/X _18752_/A vssd1 vssd1 vccd1 vccd1 _20240_/D
+ sky130_fd_sc_hd__o211a_1
X_14595_ _19361_/Q _17947_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19361_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19122_ _19698_/CLK _19122_/D vssd1 vssd1 vccd1 vccd1 _19122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ _16338_/C _16334_/B vssd1 vssd1 vccd1 vccd1 _19720_/D sky130_fd_sc_hd__nor2_1
X_13546_ _20920_/Q _13598_/A2 _18589_/B vssd1 vssd1 vccd1 vccd1 _13546_/X sky130_fd_sc_hd__a21o_1
X_10758_ _19273_/Q _20060_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10758_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19053_ _20398_/Q vssd1 vssd1 vccd1 vccd1 _20398_/D sky130_fd_sc_hd__clkbuf_2
X_16265_ _19681_/Q _17696_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19681_/D sky130_fd_sc_hd__mux2_1
X_13477_ _19830_/Q _16594_/B vssd1 vssd1 vccd1 vccd1 _13477_/X sky130_fd_sc_hd__and2_1
XFILLER_127_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10689_ _19630_/Q _19936_/Q _19274_/Q _20061_/Q _11116_/S _12406_/C vssd1 vssd1 vccd1
+ vccd1 _10689_/X sky130_fd_sc_hd__mux4_1
XFILLER_200_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18004_ _18094_/A _18004_/B _18005_/B vssd1 vssd1 vccd1 vccd1 _20739_/D sky130_fd_sc_hd__nor3_1
X_15216_ _14841_/S _15215_/X _15214_/X _15612_/S vssd1 vssd1 vccd1 vccd1 _15216_/X
+ sky130_fd_sc_hd__o211a_1
X_12428_ _19428_/Q _20587_/Q _12428_/S vssd1 vssd1 vccd1 vccd1 _12428_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16196_ _19622_/Q _16049_/X _16196_/S vssd1 vssd1 vccd1 vccd1 _16197_/B sky130_fd_sc_hd__mux2_1
XFILLER_154_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput306 _13613_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[10] sky130_fd_sc_hd__buf_4
XFILLER_160_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput317 _13623_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[20] sky130_fd_sc_hd__buf_4
X_15147_ _15396_/A1 _15130_/X _15146_/X vssd1 vssd1 vccd1 vccd1 _16743_/B sky130_fd_sc_hd__a21oi_4
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput328 _13540_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[5] sky130_fd_sc_hd__buf_4
XFILLER_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ _11201_/A _12350_/X _12358_/X _12342_/Y vssd1 vssd1 vccd1 vccd1 _12359_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_114_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput339 _13697_/Y vssd1 vssd1 vccd1 vccd1 core_wb_data_o[14] sky130_fd_sc_hd__buf_4
XFILLER_236_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15078_ _11033_/S _11219_/X _15528_/B vssd1 vssd1 vccd1 vccd1 _15078_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19955_ _20647_/CLK _19955_/D vssd1 vssd1 vccd1 vccd1 _19955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14029_ _14029_/A1 _14038_/A2 _10379_/X _14035_/B1 _19858_/Q vssd1 vssd1 vccd1 vccd1
+ _14099_/C sky130_fd_sc_hd__o32a_1
X_18906_ _19105_/Q _18954_/A2 _18974_/B1 _15762_/A vssd1 vssd1 vccd1 vccd1 _18907_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_256_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19886_ _20710_/CLK _19886_/D vssd1 vssd1 vccd1 vccd1 _19886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18837_ _18968_/A _18837_/B vssd1 vssd1 vccd1 vccd1 _18837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_256_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09570_ _12569_/A _12578_/A vssd1 vssd1 vccd1 vccd1 _13661_/A sky130_fd_sc_hd__nand2_4
XFILLER_282_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18768_ _19494_/Q _18901_/S _18766_/Y _19117_/Q vssd1 vssd1 vccd1 vccd1 _18768_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_67_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17719_ _20500_/Q _17893_/A1 _17742_/S vssd1 vssd1 vccd1 vccd1 _20500_/D sky130_fd_sc_hd__mux2_1
XFILLER_222_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18699_ _20950_/Q _18180_/Y _18707_/S vssd1 vssd1 vccd1 vccd1 _18700_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_149_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19506_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_282_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20730_ _20763_/CLK _20730_/D vssd1 vssd1 vccd1 vccd1 _20730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20661_ _20667_/CLK _20661_/D vssd1 vssd1 vccd1 vccd1 _20661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20592_ _20660_/CLK _20592_/D vssd1 vssd1 vccd1 vccd1 _20592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout500 _17813_/X vssd1 vssd1 vccd1 vccd1 _17842_/S sky130_fd_sc_hd__buf_12
Xfanout511 _17745_/X vssd1 vssd1 vccd1 vccd1 _17776_/S sky130_fd_sc_hd__buf_6
Xfanout1509 _11979_/S vssd1 vssd1 vccd1 vccd1 _11889_/S sky130_fd_sc_hd__buf_6
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout522 _17657_/S vssd1 vssd1 vccd1 vccd1 _17674_/S sky130_fd_sc_hd__buf_12
X_09906_ _11922_/A1 _13726_/A _12158_/B1 vssd1 vssd1 vccd1 vccd1 _09906_/X sky130_fd_sc_hd__o21a_1
XFILLER_160_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout533 _17540_/X vssd1 vssd1 vccd1 vccd1 _17567_/S sky130_fd_sc_hd__buf_4
XFILLER_76_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout544 _17144_/S vssd1 vssd1 vccd1 vccd1 _17146_/S sky130_fd_sc_hd__buf_12
Xfanout555 _17049_/X vssd1 vssd1 vccd1 vccd1 _17080_/S sky130_fd_sc_hd__buf_6
XFILLER_258_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout566 _16620_/S vssd1 vssd1 vccd1 vccd1 _16637_/S sky130_fd_sc_hd__buf_12
X_20026_ _20690_/CLK _20026_/D vssd1 vssd1 vccd1 vccd1 _20026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout577 _16275_/S vssd1 vssd1 vccd1 vccd1 _16277_/S sky130_fd_sc_hd__buf_12
X_09837_ _09835_/X _09836_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _09837_/X sky130_fd_sc_hd__mux2_1
XFILLER_274_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout588 _14738_/Y vssd1 vssd1 vccd1 vccd1 _14798_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout599 _14635_/X vssd1 vssd1 vccd1 vccd1 _14664_/S sky130_fd_sc_hd__buf_12
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09768_ _09765_/X _09767_/X _09776_/S vssd1 vssd1 vccd1 vccd1 _09768_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_206_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09699_ _20388_/Q _20452_/Q _11889_/S vssd1 vssd1 vccd1 vccd1 _09699_/X sky130_fd_sc_hd__mux2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11730_/A _11730_/B vssd1 vssd1 vccd1 vccd1 _13419_/A sky130_fd_sc_hd__nor2_8
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ _21025_/CLK _20928_/D vssd1 vssd1 vccd1 vccd1 _20928_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _20383_/Q _20447_/Q _11665_/S vssd1 vssd1 vccd1 vccd1 _11661_/X sky130_fd_sc_hd__mux2_1
X_20859_ _20861_/CLK _20859_/D vssd1 vssd1 vccd1 vccd1 _20859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13400_ _13205_/A _19237_/Q _16191_/A _13399_/Y vssd1 vssd1 vccd1 vccd1 _13411_/A
+ sky130_fd_sc_hd__o211a_4
X_10612_ _20406_/Q _10603_/B _10611_/X _10630_/C1 vssd1 vssd1 vccd1 vccd1 _10612_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14380_ _19240_/Q _14438_/A2 _14379_/X _14794_/C1 vssd1 vssd1 vccd1 vccd1 _19240_/D
+ sky130_fd_sc_hd__o211a_1
X_11592_ _11977_/A1 _11578_/X _11579_/X vssd1 vssd1 vccd1 vccd1 _11592_/X sky130_fd_sc_hd__o21a_1
X_13331_ _14306_/A1 _19233_/Q _14776_/C1 _13330_/X vssd1 vssd1 vccd1 vccd1 _13361_/C
+ sky130_fd_sc_hd__o211a_1
X_10543_ _19536_/Q _09596_/A _09613_/B _19600_/Q _11246_/A1 vssd1 vssd1 vccd1 vccd1
+ _10543_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16050_ _16050_/A1 _16049_/X _16037_/Y vssd1 vssd1 vccd1 vccd1 _16050_/X sky130_fd_sc_hd__a21o_1
X_13262_ _13257_/X _13261_/X _13205_/A vssd1 vssd1 vccd1 vccd1 _13262_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10474_ _19537_/Q _09596_/B _10473_/Y vssd1 vssd1 vccd1 vccd1 _10474_/X sky130_fd_sc_hd__a21o_4
XFILLER_170_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15001_ _14983_/A _14959_/B _14997_/X vssd1 vssd1 vccd1 vccd1 _15001_/Y sky130_fd_sc_hd__o21bai_1
X_12213_ _19958_/Q _12213_/B vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__or2_1
XFILLER_182_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ _18765_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13193_/Y sky130_fd_sc_hd__nor2_2
XFILLER_151_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12144_ _12144_/A1 _12143_/X _12140_/X _12144_/C1 vssd1 vssd1 vccd1 vccd1 _12144_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19740_ _20757_/CLK _19740_/D vssd1 vssd1 vccd1 vccd1 _19740_/Q sky130_fd_sc_hd__dfxtp_1
X_16952_ _16950_/Y _16951_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16952_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12075_ _13670_/A1 _17878_/A1 _12074_/X _12075_/C1 vssd1 vssd1 vccd1 vccd1 _12075_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_256_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11026_ _11026_/A _20660_/Q _11026_/C vssd1 vssd1 vccd1 vccd1 _11026_/X sky130_fd_sc_hd__or3_1
X_15903_ _15903_/A _15903_/B vssd1 vssd1 vccd1 vccd1 _15903_/Y sky130_fd_sc_hd__nor2_1
X_19671_ _20679_/CLK _19671_/D vssd1 vssd1 vccd1 vccd1 _19671_/Q sky130_fd_sc_hd__dfxtp_1
X_16883_ _19701_/Q _19698_/Q vssd1 vssd1 vccd1 vccd1 _16885_/A sky130_fd_sc_hd__nand2_8
XFILLER_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18622_ _18856_/A _18622_/B vssd1 vssd1 vccd1 vccd1 _20928_/D sky130_fd_sc_hd__nor2_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _15882_/A1 _15823_/X _15824_/X _15833_/X vssd1 vssd1 vccd1 vccd1 _15834_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_264_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ _18560_/A _18553_/B vssd1 vssd1 vccd1 vccd1 _18553_/X sky130_fd_sc_hd__or2_1
X_12977_ _19087_/Q _19086_/Q _09588_/C _12976_/Y _14112_/C vssd1 vssd1 vccd1 vccd1
+ _12978_/B sky130_fd_sc_hd__a41o_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15765_ _13415_/A _12565_/B _15983_/A _15437_/B _15764_/X vssd1 vssd1 vccd1 vccd1
+ _15765_/X sky130_fd_sc_hd__a221o_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _20287_/Q _17524_/B vssd1 vssd1 vccd1 vccd1 _17504_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14716_ _19473_/Q _17163_/A1 _14719_/S vssd1 vssd1 vccd1 vccd1 _19473_/D sky130_fd_sc_hd__mux2_1
X_11928_ _11926_/X _11927_/X _12006_/S vssd1 vssd1 vccd1 vccd1 _11928_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18484_ _20888_/Q fanout753/X _18483_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18485_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15696_ _20804_/Q _15941_/A2 _15689_/X _15882_/A1 _15695_/X vssd1 vssd1 vccd1 vccd1
+ _15696_/X sky130_fd_sc_hd__a221o_1
XFILLER_221_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_460 _19245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_471 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_482 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17435_ _17442_/A _17451_/B _17337_/B vssd1 vssd1 vccd1 vccd1 _17454_/A sky130_fd_sc_hd__o21ai_1
X_14647_ _19409_/Q _17931_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19409_/D sky130_fd_sc_hd__mux2_1
XANTENNA_493 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11859_ _19422_/Q _20581_/Q _11947_/S vssd1 vssd1 vccd1 vccd1 _11859_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_18 _15535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ _19344_/Q _17930_/A1 _14599_/S vssd1 vssd1 vccd1 vccd1 _19344_/D sky130_fd_sc_hd__mux2_1
X_17366_ _20231_/Q _17378_/A2 _17370_/B1 _20280_/Q _17370_/C1 vssd1 vssd1 vccd1 vccd1
+ _17366_/X sky130_fd_sc_hd__a221o_1
XANTENNA_29 _15820_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19105_ _19228_/CLK _19105_/D vssd1 vssd1 vccd1 vccd1 _19105_/Q sky130_fd_sc_hd__dfxtp_4
X_16317_ _19714_/Q _16316_/B _18414_/A vssd1 vssd1 vccd1 vccd1 _16318_/B sky130_fd_sc_hd__o21ai_1
XFILLER_201_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13529_ _13545_/B _13529_/B vssd1 vssd1 vccd1 vccd1 _13529_/X sky130_fd_sc_hd__and2b_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17297_ _20204_/Q _17327_/A2 _17330_/C1 vssd1 vssd1 vccd1 vccd1 _17297_/X sky130_fd_sc_hd__a21o_1
XFILLER_186_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16248_ _19664_/Q _17922_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19664_/D sky130_fd_sc_hd__mux2_1
X_19036_ _18285_/Y _19046_/A2 _19048_/B1 _12550_/C _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19036_/X sky130_fd_sc_hd__a221o_1
XFILLER_146_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16179_ _16179_/A _16179_/B vssd1 vssd1 vccd1 vccd1 _19613_/D sky130_fd_sc_hd__and2_1
XFILLER_142_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19938_ _20438_/CLK _19938_/D vssd1 vssd1 vccd1 vccd1 _19938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19869_ _20465_/CLK _19869_/D vssd1 vssd1 vccd1 vccd1 _19869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09622_ _11101_/A _10979_/C vssd1 vssd1 vccd1 vccd1 _09622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09553_ _12464_/A _12464_/C _09552_/B _12574_/A vssd1 vssd1 vccd1 vccd1 _09567_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_243_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09484_ _17402_/A vssd1 vssd1 vccd1 vccd1 _17443_/A sky130_fd_sc_hd__clkinv_4
XFILLER_52_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20713_ _20713_/CLK _20713_/D vssd1 vssd1 vccd1 vccd1 _20713_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20644_ _20676_/CLK _20644_/D vssd1 vssd1 vccd1 vccd1 _20644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20575_ _20716_/CLK _20575_/D vssd1 vssd1 vccd1 vccd1 _20575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20718_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10190_ _20410_/Q _20346_/Q _20638_/Q _20602_/Q _11211_/S _11191_/C vssd1 vssd1 vccd1
+ vccd1 _10190_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1306 _12962_/S vssd1 vssd1 vccd1 vccd1 _12964_/A2 sky130_fd_sc_hd__buf_6
Xfanout1317 _14878_/B vssd1 vssd1 vccd1 vccd1 _15984_/B1 sky130_fd_sc_hd__buf_6
XFILLER_238_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1328 _16030_/D1 vssd1 vssd1 vccd1 vccd1 _15890_/A sky130_fd_sc_hd__buf_6
XFILLER_278_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1339 _09688_/Y vssd1 vssd1 vccd1 vccd1 _09689_/D sky130_fd_sc_hd__buf_6
XFILLER_87_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12900_ _13221_/B _12900_/B vssd1 vssd1 vccd1 vccd1 _13116_/B sky130_fd_sc_hd__nor2_1
X_20009_ _20751_/CLK _20009_/D vssd1 vssd1 vccd1 vccd1 _20009_/Q sky130_fd_sc_hd__dfxtp_2
X_13880_ _19098_/Q _14527_/A2 _13900_/A2 _19164_/Q _16195_/A vssd1 vssd1 vccd1 vccd1
+ _19098_/D sky130_fd_sc_hd__o221a_1
XFILLER_272_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12831_ _12866_/A _12864_/B vssd1 vssd1 vccd1 vccd1 _13300_/A sky130_fd_sc_hd__nand2b_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _14878_/B _15549_/X _10198_/A vssd1 vssd1 vccd1 vccd1 _15550_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _19504_/Q _12782_/A vssd1 vssd1 vccd1 vccd1 _12762_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_203_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _19279_/Q _17096_/A1 _14516_/S vssd1 vssd1 vccd1 vccd1 _19279_/D sky130_fd_sc_hd__mux2_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11713_ _12102_/A1 _19352_/Q _20707_/Q _12025_/S vssd1 vssd1 vccd1 vccd1 _11713_/X
+ sky130_fd_sc_hd__a22o_1
X_15481_ _20861_/Q _15480_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15481_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _12693_/Y sky130_fd_sc_hd__nor2_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17220_ _20182_/Q _17224_/B vssd1 vssd1 vccd1 vccd1 _17220_/X sky130_fd_sc_hd__or2_1
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14432_ _14432_/A _14432_/B vssd1 vssd1 vccd1 vccd1 _14433_/B sky130_fd_sc_hd__nor2_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11872_/A _12023_/S _11641_/X _11643_/X vssd1 vssd1 vccd1 vccd1 _11644_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_174_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17151_ _17745_/A _17676_/B _17151_/C vssd1 vssd1 vccd1 vccd1 _17151_/X sky130_fd_sc_hd__and3_4
XFILLER_167_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14363_ _19518_/Q _14364_/B vssd1 vssd1 vccd1 vccd1 _14363_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11575_ _11575_/A _11575_/B vssd1 vssd1 vccd1 vccd1 _13421_/A sky130_fd_sc_hd__nor2_4
Xinput16 core_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_4
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 core_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_4
X_16102_ _11242_/X _16126_/A2 _16101_/X vssd1 vssd1 vccd1 vccd1 _19575_/D sky130_fd_sc_hd__o21a_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput38 core_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_4
X_13314_ split6/X _13310_/X _13313_/X vssd1 vssd1 vccd1 vccd1 _13314_/Y sky130_fd_sc_hd__a21oi_1
X_17082_ _17082_/A _17812_/A vssd1 vssd1 vccd1 vccd1 _17083_/C sky130_fd_sc_hd__nor2_1
X_10526_ _11290_/A _19907_/Q _11292_/S0 _20032_/Q vssd1 vssd1 vccd1 vccd1 _10526_/X
+ sky130_fd_sc_hd__o22a_1
Xinput49 dout0[15] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14294_ _14417_/S _14294_/B vssd1 vssd1 vccd1 vccd1 _14294_/X sky130_fd_sc_hd__or2_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16033_ _16005_/A1 _12617_/Y _16032_/X _12708_/B vssd1 vssd1 vccd1 vccd1 _16033_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ _13245_/A _13245_/B vssd1 vssd1 vccd1 vccd1 _16241_/B sky130_fd_sc_hd__nand2_1
X_10457_ _19537_/Q _09596_/A _09613_/B _19601_/Q _11246_/A1 vssd1 vssd1 vccd1 vccd1
+ _10457_/Y sky130_fd_sc_hd__a221oi_4
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _12199_/B _13183_/B _12197_/Y vssd1 vssd1 vccd1 vccd1 _13182_/B sky130_fd_sc_hd__a21oi_4
XFILLER_112_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10388_ _19777_/Q _11305_/B _11304_/S vssd1 vssd1 vccd1 vccd1 _10388_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12127_ _20146_/Q _20114_/Q _12133_/S vssd1 vssd1 vccd1 vccd1 _12127_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_5__f_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17984_ _17984_/A _17984_/B vssd1 vssd1 vccd1 vccd1 _20732_/D sky130_fd_sc_hd__nor2_1
XFILLER_257_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19723_ _21026_/CLK _19723_/D vssd1 vssd1 vccd1 vccd1 _19723_/Q sky130_fd_sc_hd__dfxtp_1
X_16935_ _16932_/Y _16934_/Y _16822_/A vssd1 vssd1 vccd1 vccd1 _16935_/Y sky130_fd_sc_hd__a21oi_4
Xfanout1840 _12125_/A1 vssd1 vssd1 vccd1 vccd1 _11514_/A1 sky130_fd_sc_hd__buf_8
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12058_ _12056_/X _12057_/X _12058_/S vssd1 vssd1 vccd1 vccd1 _12058_/X sky130_fd_sc_hd__mux2_1
Xfanout1851 _11281_/A vssd1 vssd1 vccd1 vccd1 _13192_/A sky130_fd_sc_hd__buf_12
XFILLER_238_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1862 _12850_/A1 vssd1 vssd1 vccd1 vccd1 _12020_/C1 sky130_fd_sc_hd__buf_6
XFILLER_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1873 _19166_/Q vssd1 vssd1 vccd1 vccd1 _12504_/B sky130_fd_sc_hd__buf_6
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1884 _19116_/Q vssd1 vssd1 vccd1 vccd1 _14112_/A sky130_fd_sc_hd__buf_4
X_11009_ _19801_/Q _11009_/A2 _11007_/X _11009_/B2 _11008_/X vssd1 vssd1 vccd1 vccd1
+ _11009_/X sky130_fd_sc_hd__o221a_1
X_19654_ _20664_/CLK _19654_/D vssd1 vssd1 vccd1 vccd1 _19654_/Q sky130_fd_sc_hd__dfxtp_1
X_16866_ _16982_/B1 _16863_/X _16865_/X _16866_/B2 vssd1 vssd1 vccd1 vccd1 _16867_/B
+ sky130_fd_sc_hd__o2bb2a_4
Xfanout1895 _18734_/A vssd1 vssd1 vccd1 vccd1 _18740_/A sky130_fd_sc_hd__buf_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18605_ _18496_/X _18621_/A2 _18603_/Y _18604_/Y vssd1 vssd1 vccd1 vccd1 _18606_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_225_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15817_ _11748_/Y _15925_/B _15219_/Y _15816_/Y vssd1 vssd1 vccd1 vccd1 _15817_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_280_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19585_ _20665_/CLK _19585_/D vssd1 vssd1 vccd1 vccd1 _19585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16797_ _19222_/Q _16862_/A2 _16713_/X _16794_/Y _16796_/X vssd1 vssd1 vccd1 vccd1
+ _16797_/X sky130_fd_sc_hd__o2111a_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18536_ _20905_/Q fanout750/X _18535_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18537_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _20934_/Q _16044_/A2 _15747_/X vssd1 vssd1 vccd1 vccd1 _15748_/X sky130_fd_sc_hd__o21a_1
XFILLER_252_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18467_ _18474_/S _18467_/B vssd1 vssd1 vccd1 vccd1 _18467_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_290 input221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15679_ _19544_/Q _16007_/A _15677_/X _15678_/X _16189_/A vssd1 vssd1 vccd1 vccd1
+ _19544_/D sky130_fd_sc_hd__o221a_1
XFILLER_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17418_ _17443_/A _17420_/A _20256_/Q vssd1 vssd1 vccd1 vccd1 _17418_/Y sky130_fd_sc_hd__o21ai_1
X_18398_ _18418_/A _18398_/B vssd1 vssd1 vccd1 vccd1 _20853_/D sky130_fd_sc_hd__and2_1
X_17349_ _20223_/Q _17363_/A2 _17348_/X _18692_/A vssd1 vssd1 vccd1 vccd1 _20223_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20360_ _20706_/CLK _20360_/D vssd1 vssd1 vccd1 vccd1 _20360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19019_ _21028_/Q _19015_/B _19018_/X _18724_/A vssd1 vssd1 vccd1 vccd1 _21028_/D
+ sky130_fd_sc_hd__o211a_1
X_20291_ _20291_/CLK _20291_/D vssd1 vssd1 vccd1 vccd1 _20291_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_88_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_164_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21011_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09605_ _09610_/A _19090_/Q _19089_/Q _19088_/Q vssd1 vssd1 vccd1 vccd1 _09606_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_84_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_260_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09536_ _19156_/Q _19155_/Q _13869_/A vssd1 vssd1 vccd1 vccd1 _12480_/A sky130_fd_sc_hd__and3_2
XFILLER_243_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20627_ _20686_/CLK _20627_/D vssd1 vssd1 vccd1 vccd1 _20627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ _12230_/A1 _19905_/Q _11359_/S _11348_/X vssd1 vssd1 vccd1 vccd1 _11360_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20558_ _20690_/CLK _20558_/D vssd1 vssd1 vccd1 vccd1 _20558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10311_ _20036_/Q _10485_/S vssd1 vssd1 vccd1 vccd1 _10311_/X sky130_fd_sc_hd__or2_1
XFILLER_285_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11291_ _19366_/Q _11291_/A2 _11289_/X _11291_/B2 _11290_/X vssd1 vssd1 vccd1 vccd1
+ _11291_/X sky130_fd_sc_hd__o221a_1
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20489_ _20641_/CLK _20489_/D vssd1 vssd1 vccd1 vccd1 _20489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030_ _20964_/Q _20898_/Q vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__nand2_2
X_10242_ _12245_/A1 _17901_/A1 _10241_/X vssd1 vssd1 vccd1 vccd1 _13698_/A sky130_fd_sc_hd__o21ai_4
XFILLER_180_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10173_ _10262_/A _19475_/Q _19443_/Q _10174_/S vssd1 vssd1 vccd1 vccd1 _10173_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1103 _12040_/X vssd1 vssd1 vccd1 vccd1 _17878_/A1 sky130_fd_sc_hd__buf_6
XFILLER_79_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1114 _17876_/A1 vssd1 vssd1 vccd1 vccd1 _17910_/A1 sky130_fd_sc_hd__buf_4
Xfanout1125 _17902_/A1 vssd1 vssd1 vccd1 vccd1 _17693_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1136 _09947_/X vssd1 vssd1 vccd1 vccd1 _17800_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_94_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1147 _17908_/A1 vssd1 vssd1 vccd1 vccd1 _17874_/A1 sky130_fd_sc_hd__clkbuf_4
X_14981_ _14981_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _15022_/C sky130_fd_sc_hd__or2_2
Xfanout1158 _09631_/X vssd1 vssd1 vccd1 vccd1 _12074_/B1 sky130_fd_sc_hd__buf_4
XFILLER_282_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1169 _14897_/Y vssd1 vssd1 vccd1 vccd1 _15644_/A1 sky130_fd_sc_hd__buf_6
X_16720_ _16720_/A _16720_/B _16720_/C _16720_/D vssd1 vssd1 vccd1 vccd1 _16720_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_75_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13932_ _19136_/Q _13941_/B _13932_/B1 _13361_/A vssd1 vssd1 vccd1 vccd1 _19136_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_262_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13863_ _13863_/A _13863_/B vssd1 vssd1 vccd1 vccd1 _13863_/Y sky130_fd_sc_hd__nand2_1
X_16651_ _19908_/Q _17095_/A1 _16666_/S vssd1 vssd1 vccd1 vccd1 _19908_/D sky130_fd_sc_hd__mux2_1
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15602_ input270/X _15013_/Y _15596_/X _15606_/A1 vssd1 vssd1 vccd1 vccd1 _15602_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_216_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12814_ _12906_/A _12815_/B vssd1 vssd1 vccd1 vccd1 _13264_/B sky130_fd_sc_hd__nand2_1
XFILLER_234_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19370_ _20667_/CLK _19370_/D vssd1 vssd1 vccd1 vccd1 _19370_/Q sky130_fd_sc_hd__dfxtp_1
X_16582_ _19857_/Q _16592_/A2 _16592_/B1 input28/X vssd1 vssd1 vccd1 vccd1 _16583_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13794_ _13798_/A1 _13826_/A1 _13718_/B _13826_/B1 input240/X vssd1 vssd1 vccd1 vccd1
+ _13794_/X sky130_fd_sc_hd__a32o_1
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18321_ _18981_/C _18323_/B _18139_/B vssd1 vssd1 vccd1 vccd1 _18755_/A sky130_fd_sc_hd__or3b_1
XFILLER_231_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15533_ _20895_/Q _15937_/A2 _15566_/B1 _15532_/X _15937_/C1 vssd1 vssd1 vccd1 vccd1
+ _15533_/X sky130_fd_sc_hd__a221o_1
X_12745_ _12464_/A _09541_/Y split6/A _12710_/B vssd1 vssd1 vccd1 vccd1 _12747_/C
+ sky130_fd_sc_hd__o211a_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _18724_/A _18252_/B vssd1 vssd1 vccd1 vccd1 _20804_/D sky130_fd_sc_hd__and2_1
X_15464_ _13459_/Y _15494_/B _15219_/Y vssd1 vssd1 vccd1 vccd1 _15465_/B sky130_fd_sc_hd__o21a_1
XFILLER_230_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12676_ _12676_/A _12676_/B vssd1 vssd1 vccd1 vccd1 _13501_/C sky130_fd_sc_hd__nor2_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _14400_/Y _14405_/B _14402_/B vssd1 vssd1 vccd1 vccd1 _14424_/B sky130_fd_sc_hd__o21ai_2
X_17203_ _20167_/Q _17869_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20167_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11627_ _20416_/Q _20352_/Q _20644_/Q _20608_/Q _11932_/S0 _12008_/C vssd1 vssd1
+ vccd1 vccd1 _11627_/X sky130_fd_sc_hd__mux4_1
X_15395_ _19710_/Q _15394_/X _15395_/S vssd1 vssd1 vccd1 vccd1 _15395_/X sky130_fd_sc_hd__mux2_2
X_18183_ _19532_/Q _18213_/B vssd1 vssd1 vccd1 vccd1 _18183_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14346_ _14427_/A _14342_/B _14345_/X vssd1 vssd1 vccd1 vccd1 _14346_/X sky130_fd_sc_hd__a21bo_1
X_17134_ _20102_/Q _17202_/A1 _17146_/S vssd1 vssd1 vccd1 vccd1 _20102_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11558_ _11946_/A1 _19350_/Q _20705_/Q _11860_/B2 vssd1 vssd1 vccd1 vccd1 _11558_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17065_ _20037_/Q _17099_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20037_/D sky130_fd_sc_hd__mux2_1
X_10509_ _19504_/Q _15589_/S vssd1 vssd1 vccd1 vccd1 _10509_/Y sky130_fd_sc_hd__nor2_2
XFILLER_171_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14277_ _19230_/Q _14398_/A2 _14276_/X _14772_/C1 vssd1 vssd1 vccd1 vccd1 _19230_/D
+ sky130_fd_sc_hd__o211a_1
X_11489_ _11487_/X _11488_/X _12189_/A vssd1 vssd1 vccd1 vccd1 _11489_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16016_ _16015_/X _20848_/Q _16016_/S vssd1 vssd1 vccd1 vccd1 _16016_/X sky130_fd_sc_hd__mux2_1
X_13228_ _20972_/Q _13397_/B _13226_/Y _13227_/Y _18767_/A vssd1 vssd1 vccd1 vccd1
+ _13229_/C sky130_fd_sc_hd__a221o_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _10367_/Y _13423_/B _15580_/S vssd1 vssd1 vccd1 vccd1 _13422_/B sky130_fd_sc_hd__a21bo_4
XFILLER_98_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _20726_/Q _17965_/B _17966_/Y vssd1 vssd1 vccd1 vccd1 _20726_/D sky130_fd_sc_hd__o21a_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19706_ _20759_/CLK _19706_/D vssd1 vssd1 vccd1 vccd1 _19706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_254_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1670 _14029_/A1 vssd1 vssd1 vccd1 vccd1 _14041_/A1 sky130_fd_sc_hd__buf_4
X_16918_ _16885_/A _16917_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16918_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_239_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1681 _12008_/A vssd1 vssd1 vccd1 vccd1 _12007_/A1 sky130_fd_sc_hd__buf_4
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1692 _11021_/A vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__clkbuf_8
X_17898_ _20669_/Q _17898_/A1 _17912_/S vssd1 vssd1 vccd1 vccd1 _20669_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19637_ _20539_/CLK _19637_/D vssd1 vssd1 vccd1 vccd1 _19637_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 ANTENNA_548/DIODE sky130_fd_sc_hd__clkbuf_16
XFILLER_81_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16849_ _16849_/A _16849_/B vssd1 vssd1 vccd1 vccd1 _16849_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19568_ _19577_/CLK _19568_/D vssd1 vssd1 vccd1 vccd1 _19568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_281_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18519_ _18891_/A _18519_/B vssd1 vssd1 vccd1 vccd1 _20899_/D sky130_fd_sc_hd__nor2_1
XFILLER_22_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19499_ _19505_/CLK _19499_/D vssd1 vssd1 vccd1 vccd1 _19499_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20412_ _20465_/CLK _20412_/D vssd1 vssd1 vccd1 vccd1 _20412_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_175_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20343_ _20635_/CLK _20343_/D vssd1 vssd1 vccd1 vccd1 _20343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20274_ _20818_/CLK _20274_/D vssd1 vssd1 vccd1 vccd1 _20274_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_249_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput206 localMemory_wb_adr_i[2] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput217 localMemory_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_hd__buf_12
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput228 localMemory_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_hd__buf_12
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput239 localMemory_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_hd__buf_12
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10860_ _20402_/Q _20338_/Q _20630_/Q _20594_/Q _12352_/S _12337_/C vssd1 vssd1 vccd1
+ vccd1 _10860_/X sky130_fd_sc_hd__mux4_1
XFILLER_232_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09519_ input54/X vssd1 vssd1 vccd1 vccd1 _09519_/Y sky130_fd_sc_hd__inv_2
XFILLER_213_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10791_ _12427_/A1 _19340_/Q _20695_/Q _11126_/B _12419_/C1 vssd1 vssd1 vccd1 vccd1
+ _10791_/X sky130_fd_sc_hd__a221o_1
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12530_ _13552_/A _19215_/Q _12529_/X vssd1 vssd1 vccd1 vccd1 _13478_/A sky130_fd_sc_hd__o21a_4
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20687_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12461_ _14894_/A _14897_/A vssd1 vssd1 vccd1 vccd1 _15468_/A sky130_fd_sc_hd__nor2_8
XFILLER_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14200_ _14189_/A _14191_/B _14189_/B vssd1 vssd1 vccd1 vccd1 _14201_/B sky130_fd_sc_hd__a21boi_4
XFILLER_138_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11412_ _10112_/A _11412_/B vssd1 vssd1 vccd1 vccd1 _11754_/A sky130_fd_sc_hd__and2b_1
X_15180_ _14885_/B _14839_/X _15215_/S vssd1 vssd1 vccd1 vccd1 _15180_/X sky130_fd_sc_hd__mux2_1
X_12392_ _12399_/A1 _12391_/X _12388_/X _12392_/C1 vssd1 vssd1 vccd1 vccd1 _12392_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _14131_/A _14131_/B vssd1 vssd1 vccd1 vccd1 _14131_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_153_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11343_ _11341_/X _11342_/X _12376_/S vssd1 vssd1 vccd1 vccd1 _11343_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14062_ _19190_/Q _14082_/A2 _14061_/X _16143_/A vssd1 vssd1 vccd1 vccd1 _19190_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11274_ _19798_/Q _09689_/D _11272_/X _11274_/B2 _11273_/X vssd1 vssd1 vccd1 vccd1
+ _11275_/C sky130_fd_sc_hd__o221a_1
XFILLER_106_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13013_ _20972_/Q _20906_/Q vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__and2_2
X_10225_ _20540_/Q _10986_/B vssd1 vssd1 vccd1 vccd1 _10225_/X sky130_fd_sc_hd__or2_1
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18870_ _18877_/A _18870_/B vssd1 vssd1 vccd1 vccd1 _20995_/D sky130_fd_sc_hd__nor2_1
XFILLER_95_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17821_ _20596_/Q _17893_/A1 _17844_/S vssd1 vssd1 vccd1 vccd1 _20596_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10156_ _10154_/X _10155_/X _11359_/S vssd1 vssd1 vccd1 vccd1 _10156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17752_ _20531_/Q _17892_/A1 _17776_/S vssd1 vssd1 vccd1 vccd1 _20531_/D sky130_fd_sc_hd__mux2_1
X_14964_ _14983_/A _15020_/A vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__or2_2
X_10087_ _10082_/X _10086_/X _15678_/A1 vssd1 vssd1 vccd1 vccd1 _10087_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16703_ _19958_/Q _17915_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19958_/D sky130_fd_sc_hd__mux2_1
XFILLER_247_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13915_ _13915_/A _13919_/S vssd1 vssd1 vccd1 vccd1 _13915_/Y sky130_fd_sc_hd__nand2_1
X_17683_ _20467_/Q _17683_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20467_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14895_ _14895_/A _15096_/A vssd1 vssd1 vccd1 vccd1 _14895_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19422_ _20713_/CLK _19422_/D vssd1 vssd1 vccd1 vccd1 _19422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16634_ _19893_/Q _17112_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19893_/D sky130_fd_sc_hd__mux2_1
XFILLER_235_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13846_ _20261_/Q _20258_/Q _13846_/C vssd1 vssd1 vccd1 vccd1 _17335_/B sky130_fd_sc_hd__nor3_4
XFILLER_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19353_ _20708_/CLK _19353_/D vssd1 vssd1 vccd1 vccd1 _19353_/Q sky130_fd_sc_hd__dfxtp_1
X_16565_ _16593_/A _16565_/B vssd1 vssd1 vccd1 vccd1 _19848_/D sky130_fd_sc_hd__or2_1
XFILLER_204_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13777_ _13777_/A _13777_/B vssd1 vssd1 vccd1 vccd1 _13777_/X sky130_fd_sc_hd__or2_1
X_10989_ _11336_/A _20692_/Q _10986_/B _10987_/X _10988_/X vssd1 vssd1 vccd1 vccd1
+ _10989_/X sky130_fd_sc_hd__a311o_1
XFILLER_16_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18304_ _18313_/B _14413_/B _18303_/Y vssd1 vssd1 vccd1 vccd1 _18553_/B sky130_fd_sc_hd__o21ai_4
X_15516_ _19714_/Q _15395_/S _15515_/X vssd1 vssd1 vccd1 vccd1 _15516_/X sky130_fd_sc_hd__o21a_1
XFILLER_231_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19284_ _20446_/CLK _19284_/D vssd1 vssd1 vccd1 vccd1 _19284_/Q sky130_fd_sc_hd__dfxtp_1
X_12728_ _19506_/Q _12754_/A vssd1 vssd1 vccd1 vccd1 _12729_/B sky130_fd_sc_hd__nor2_1
X_16496_ _19803_/Q _17751_/A1 _16521_/S vssd1 vssd1 vccd1 vccd1 _19803_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18235_ _18511_/B vssd1 vssd1 vccd1 vccd1 _18235_/Y sky130_fd_sc_hd__inv_4
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12659_ _12657_/X _12658_/Y _12752_/B vssd1 vssd1 vccd1 vccd1 _12662_/B sky130_fd_sc_hd__a21o_1
X_15447_ _20892_/Q _14971_/A _15566_/B1 _15446_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15447_/X sky130_fd_sc_hd__a221o_1
XFILLER_276_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18166_ _20787_/Q _18165_/Y _18236_/S vssd1 vssd1 vccd1 vccd1 _18167_/B sky130_fd_sc_hd__mux2_1
XFILLER_157_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15378_ _15378_/A _15378_/B _15377_/X vssd1 vssd1 vccd1 vccd1 _15378_/X sky130_fd_sc_hd__or3b_1
XFILLER_209_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17117_ _17745_/A _17676_/B _17117_/C vssd1 vssd1 vccd1 vccd1 _17117_/X sky130_fd_sc_hd__and3_4
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ _19235_/Q _14438_/A2 _14328_/X _14780_/C1 vssd1 vssd1 vccd1 vccd1 _19235_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18097_ _20773_/Q _18095_/B _18096_/Y vssd1 vssd1 vccd1 vccd1 _20773_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17048_ _17082_/A _17744_/A vssd1 vssd1 vccd1 vccd1 _17049_/C sky130_fd_sc_hd__nor2_1
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _12156_/A1 _09869_/X _09865_/X vssd1 vssd1 vccd1 vccd1 _09870_/X sky130_fd_sc_hd__a21o_1
Xfanout907 _16042_/A2 vssd1 vssd1 vccd1 vccd1 _16018_/A2 sky130_fd_sc_hd__buf_6
XFILLER_258_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout918 _16041_/A2 vssd1 vssd1 vccd1 vccd1 _15445_/A2 sky130_fd_sc_hd__buf_4
XFILLER_135_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout929 _15595_/A2 vssd1 vssd1 vccd1 vccd1 _15475_/A2 sky130_fd_sc_hd__buf_6
XFILLER_140_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ _21019_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _18999_/X sky130_fd_sc_hd__or2_1
XFILLER_86_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20961_ _20962_/CLK _20961_/D vssd1 vssd1 vccd1 vccd1 _20961_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_227_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20892_ _20990_/CLK _20892_/D vssd1 vssd1 vccd1 vccd1 _20892_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_198_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20326_ _20714_/CLK _20326_/D vssd1 vssd1 vccd1 vccd1 _20326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20257_ _20261_/CLK _20257_/D vssd1 vssd1 vccd1 vccd1 _20257_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_103_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ _10006_/X _10009_/X _11949_/S vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20188_ _20688_/CLK _20188_/D vssd1 vssd1 vccd1 vccd1 _20188_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ _11946_/A1 _20385_/Q _20449_/Q _11944_/S _11946_/C1 vssd1 vssd1 vccd1 vccd1
+ _09999_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11961_ _13434_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__or2_1
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10912_ _20561_/Q _12295_/B _10911_/X _11338_/A1 vssd1 vssd1 vccd1 vccd1 _10912_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _13735_/A _13698_/X _13699_/Y _13659_/A vssd1 vssd1 vccd1 vccd1 _13702_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_245_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _19439_/Q _17929_/A1 _14699_/S vssd1 vssd1 vccd1 vccd1 _19439_/D sky130_fd_sc_hd__mux2_1
X_11892_ _20582_/Q _11897_/B _11891_/X _11892_/C1 vssd1 vssd1 vccd1 vccd1 _11892_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13631_ _13714_/S _13631_/B vssd1 vssd1 vccd1 vccd1 _16233_/B sky130_fd_sc_hd__nor2_8
X_10843_ _19272_/Q _20059_/Q _12323_/S vssd1 vssd1 vccd1 vccd1 _10843_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13562_ _13049_/Y _13050_/X _13051_/X _13064_/X vssd1 vssd1 vccd1 vccd1 _13562_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16350_ _16354_/C _16350_/B vssd1 vssd1 vccd1 vccd1 _19726_/D sky130_fd_sc_hd__nor2_1
X_10774_ _19372_/Q _12255_/A2 _10772_/X _09738_/A _10773_/X vssd1 vssd1 vccd1 vccd1
+ _10774_/X sky130_fd_sc_hd__o221a_1
XFILLER_201_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12513_ _12513_/A _12513_/B _12513_/C _12513_/D vssd1 vssd1 vccd1 vccd1 _12588_/C
+ sky130_fd_sc_hd__or4_1
X_15301_ _15303_/B _15127_/B _15220_/A vssd1 vssd1 vccd1 vccd1 _15301_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16281_ _20622_/Q _17015_/B _19701_/D vssd1 vssd1 vccd1 vccd1 _19697_/D sky130_fd_sc_hd__and3_1
XFILLER_12_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13493_ _16241_/A _13907_/A vssd1 vssd1 vccd1 vccd1 _13493_/Y sky130_fd_sc_hd__nor2_2
XFILLER_185_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18020_ _18104_/A _18020_/B _18024_/C vssd1 vssd1 vccd1 vccd1 _20745_/D sky130_fd_sc_hd__nor3_1
X_15232_ input5/X _15334_/B vssd1 vssd1 vccd1 vccd1 _15232_/X sky130_fd_sc_hd__or2_1
X_12444_ _12450_/B _12444_/B vssd1 vssd1 vccd1 vccd1 _12445_/B sky130_fd_sc_hd__and2_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15163_ _15163_/A vssd1 vssd1 vccd1 vccd1 _15163_/Y sky130_fd_sc_hd__inv_2
X_12375_ _20148_/Q _20116_/Q _12375_/S vssd1 vssd1 vccd1 vccd1 _12375_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14114_ _12584_/A _14111_/Y _14113_/X vssd1 vssd1 vccd1 vccd1 _14114_/X sky130_fd_sc_hd__o21a_1
XFILLER_158_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11326_ _11326_/A _11326_/B _11326_/C vssd1 vssd1 vccd1 vccd1 _11326_/X sky130_fd_sc_hd__and3_1
X_19971_ _20268_/CLK _19971_/D vssd1 vssd1 vccd1 vccd1 _19971_/Q sky130_fd_sc_hd__dfxtp_1
X_15094_ _15644_/A1 _16732_/B _15078_/X vssd1 vssd1 vccd1 vccd1 _15094_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_180_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14045_ _14081_/A _16133_/B _14045_/C vssd1 vssd1 vccd1 vccd1 _14045_/X sky130_fd_sc_hd__or3_1
X_18922_ _18655_/Y _18970_/A2 _18920_/Y _18921_/Y vssd1 vssd1 vccd1 vccd1 _18922_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11257_ _19865_/Q _19766_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _11257_/X sky130_fd_sc_hd__mux2_1
X_10208_ _20476_/Q _20316_/Q _10217_/S vssd1 vssd1 vccd1 vccd1 _10208_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18853_ _18616_/Y _18867_/A2 _18851_/Y _18852_/Y vssd1 vssd1 vccd1 vccd1 _18853_/X
+ sky130_fd_sc_hd__a22o_1
X_11188_ _15155_/S vssd1 vssd1 vccd1 vccd1 _15067_/S sky130_fd_sc_hd__inv_2
XFILLER_122_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17804_ _20581_/Q _17804_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20581_/D sky130_fd_sc_hd__mux2_1
X_10139_ _11338_/A1 _10136_/X _10138_/X vssd1 vssd1 vccd1 vccd1 _10139_/X sky130_fd_sc_hd__a21o_1
X_18784_ _19120_/Q _18968_/A vssd1 vssd1 vccd1 vccd1 _18784_/X sky130_fd_sc_hd__or2_1
XFILLER_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15996_ _20975_/Q _16045_/A2 _15996_/B1 _20847_/Q _15995_/X vssd1 vssd1 vccd1 vccd1
+ _15996_/X sky130_fd_sc_hd__a221o_1
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17735_ _20516_/Q _17909_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20516_/D sky130_fd_sc_hd__mux2_1
X_14947_ _20722_/Q _15445_/A2 _15445_/B1 _20754_/Q vssd1 vssd1 vccd1 vccd1 _14947_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17666_ _20452_/Q _17666_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20452_/D sky130_fd_sc_hd__mux2_1
X_14878_ _14878_/A _14878_/B vssd1 vssd1 vccd1 vccd1 _14878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19405_ _20586_/CLK _19405_/D vssd1 vssd1 vccd1 vccd1 _19405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16617_ _19876_/Q _17163_/A1 _16620_/S vssd1 vssd1 vccd1 vccd1 _19876_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13829_ _19999_/Q split1/A _13783_/X split2/X vssd1 vssd1 vccd1 vccd1 _13829_/X sky130_fd_sc_hd__a22o_4
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17597_ _20355_/Q _09790_/X _17601_/S vssd1 vssd1 vccd1 vccd1 _20355_/D sky130_fd_sc_hd__mux2_1
XFILLER_245_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_250_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19336_ _20720_/CLK _19336_/D vssd1 vssd1 vccd1 vccd1 _19336_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16548_ _19840_/Q _16566_/A2 _16566_/B1 input41/X vssd1 vssd1 vccd1 vccd1 _16549_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_206_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19267_ _20315_/CLK _19267_/D vssd1 vssd1 vccd1 vccd1 _19267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16479_ _19788_/Q _17802_/A1 _16483_/S vssd1 vssd1 vccd1 vccd1 _19788_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18218_ _19539_/Q _18248_/B vssd1 vssd1 vccd1 vccd1 _18218_/Y sky130_fd_sc_hd__nand2b_2
X_19198_ _20659_/CLK _19198_/D vssd1 vssd1 vccd1 vccd1 _19198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18149_ _12945_/A _19115_/Q _18149_/S vssd1 vssd1 vccd1 vccd1 _18318_/B sky130_fd_sc_hd__mux2_1
XFILLER_116_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20111_ _20482_/CLK _20111_/D vssd1 vssd1 vccd1 vccd1 _20111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09922_ _09986_/A _20386_/Q _20450_/Q _09928_/S _11946_/C1 vssd1 vssd1 vccd1 vccd1
+ _09922_/X sky130_fd_sc_hd__a221o_1
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout704 _16578_/A2 vssd1 vssd1 vccd1 vccd1 _16576_/A2 sky130_fd_sc_hd__buf_4
Xfanout715 _16578_/B1 vssd1 vssd1 vccd1 vccd1 _16576_/B1 sky130_fd_sc_hd__buf_4
Xfanout726 _13481_/A vssd1 vssd1 vccd1 vccd1 _13626_/A1 sky130_fd_sc_hd__buf_4
X_20042_ _20677_/CLK _20042_/D vssd1 vssd1 vccd1 vccd1 _20042_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout737 _18982_/X vssd1 vssd1 vccd1 vccd1 _19048_/C1 sky130_fd_sc_hd__clkbuf_4
X_09853_ _09829_/A _20387_/Q _20451_/Q _10397_/S vssd1 vssd1 vccd1 vccd1 _09853_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout748 _18985_/B vssd1 vssd1 vccd1 vccd1 _19048_/A2 sky130_fd_sc_hd__buf_4
XFILLER_259_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout759 _18840_/B vssd1 vssd1 vccd1 vccd1 _18819_/B sky130_fd_sc_hd__buf_6
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09784_ _09784_/A _09784_/B vssd1 vssd1 vccd1 vccd1 _13413_/A sky130_fd_sc_hd__nor2_8
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_108 _13474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_269_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20944_ _21000_/CLK _20944_/D vssd1 vssd1 vccd1 vccd1 _20944_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_119 _16239_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20875_ _21040_/CLK _20875_/D vssd1 vssd1 vccd1 vccd1 _20875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _20635_/Q _10897_/A3 _11274_/B2 vssd1 vssd1 vccd1 vccd1 _10490_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _19165_/Q _19925_/Q _12464_/C vssd1 vssd1 vccd1 vccd1 _12160_/X sky130_fd_sc_hd__and3_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _19368_/Q _12255_/A2 _11109_/X _12412_/B2 _11110_/X vssd1 vssd1 vccd1 vccd1
+ _11111_/X sky130_fd_sc_hd__o221a_1
X_20309_ _20718_/CLK _20309_/D vssd1 vssd1 vccd1 vccd1 _20309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12091_ _12089_/X _12090_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _12091_/X sky130_fd_sc_hd__mux2_1
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _19665_/Q _11042_/B vssd1 vssd1 vccd1 vccd1 _11042_/X sky130_fd_sc_hd__or2_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15850_ _19726_/Q _15961_/A2 _15961_/B1 _19758_/Q vssd1 vssd1 vccd1 vccd1 _15850_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _19525_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14801_/X sky130_fd_sc_hd__or2_1
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15781_ _15973_/A1 _15780_/X _15768_/X vssd1 vssd1 vccd1 vccd1 _15781_/X sky130_fd_sc_hd__a21o_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _19236_/Q _19235_/Q _19234_/Q _13296_/B vssd1 vssd1 vccd1 vccd1 _13390_/B
+ sky130_fd_sc_hd__and4_4
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _20295_/Q _17522_/B vssd1 vssd1 vccd1 vccd1 _17520_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _19489_/Q _17947_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19489_/D sky130_fd_sc_hd__mux2_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ _20143_/Q _20111_/Q _11944_/S vssd1 vssd1 vccd1 vccd1 _11944_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_620 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_631 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_642 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17451_ _17451_/A _17451_/B vssd1 vssd1 vccd1 vccd1 _17456_/B sky130_fd_sc_hd__or2_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_653 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11875_ _19518_/Q _15849_/A _15895_/S vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__mux2_8
X_14663_ _19425_/Q _17947_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19425_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _19745_/Q _19746_/Q _16402_/C vssd1 vssd1 vccd1 vccd1 _16404_/B sky130_fd_sc_hd__and3_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ _20123_/Q _20091_/Q _12300_/S vssd1 vssd1 vccd1 vccd1 _10826_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13614_ _19661_/D _13458_/Y _13459_/Y _13663_/B vssd1 vssd1 vccd1 vccd1 _13614_/X
+ sky130_fd_sc_hd__a22o_4
X_17382_ _20239_/Q _17390_/A2 _17382_/B1 _20288_/Q _17400_/C1 vssd1 vssd1 vccd1 vccd1
+ _17382_/X sky130_fd_sc_hd__a221o_1
X_14594_ _19360_/Q _17806_/A1 _14594_/S vssd1 vssd1 vccd1 vccd1 _19360_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19121_ _19505_/CLK _19121_/D vssd1 vssd1 vccd1 vccd1 _19121_/Q sky130_fd_sc_hd__dfxtp_1
X_16333_ _19720_/Q _16332_/B _18720_/A vssd1 vssd1 vccd1 vccd1 _16334_/B sky130_fd_sc_hd__o21ai_1
X_10757_ _12396_/A1 _19903_/Q _12395_/S _10740_/X vssd1 vssd1 vccd1 vccd1 _10757_/X
+ sky130_fd_sc_hd__o211a_1
X_13545_ _19221_/Q _13545_/B vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__or2_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19052_ _20397_/Q vssd1 vssd1 vccd1 vccd1 _20397_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13476_ _13469_/Y _13472_/A _13474_/X vssd1 vssd1 vccd1 vccd1 _13476_/X sky130_fd_sc_hd__a21o_1
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16264_ _19680_/Q _17695_/A1 _16272_/S vssd1 vssd1 vccd1 vccd1 _19680_/D sky130_fd_sc_hd__mux2_1
X_10688_ _19805_/Q _12412_/A2 _10686_/X _12412_/B2 _10687_/X vssd1 vssd1 vccd1 vccd1
+ _10688_/X sky130_fd_sc_hd__o221a_1
XFILLER_173_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18003_ _20739_/Q _20738_/Q _18003_/C vssd1 vssd1 vccd1 vccd1 _18005_/B sky130_fd_sc_hd__and3_1
XFILLER_127_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12427_ _12427_/A1 _19364_/Q _20719_/Q _12428_/S _11378_/S vssd1 vssd1 vccd1 vccd1
+ _12427_/X sky130_fd_sc_hd__a221o_1
X_15215_ _14848_/X _14865_/X _15215_/S vssd1 vssd1 vccd1 vccd1 _15215_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16195_ _16195_/A _16195_/B vssd1 vssd1 vccd1 vccd1 _19621_/D sky130_fd_sc_hd__and2_1
XFILLER_127_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput307 _13614_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[11] sky130_fd_sc_hd__buf_4
X_12358_ _11118_/A _12353_/Y _12355_/Y _12357_/Y _12431_/A1 vssd1 vssd1 vccd1 vccd1
+ _12358_/X sky130_fd_sc_hd__a221o_1
X_15146_ _19704_/Q _15145_/X _15454_/S vssd1 vssd1 vccd1 vccd1 _15146_/X sky130_fd_sc_hd__mux2_2
Xoutput318 _13624_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[21] sky130_fd_sc_hd__buf_4
Xoutput329 _13555_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[6] sky130_fd_sc_hd__buf_4
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11309_ _11309_/A1 _11304_/X _11308_/X _10260_/S vssd1 vssd1 vccd1 vccd1 _11309_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15077_ _15075_/A _15075_/B _15185_/B _15075_/Y vssd1 vssd1 vccd1 vccd1 _15077_/X
+ sky130_fd_sc_hd__o211a_1
X_19954_ _20047_/CLK _19954_/D vssd1 vssd1 vccd1 vccd1 _19954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12289_ _15982_/A _15982_/B _11748_/Y _11883_/X _12207_/Y vssd1 vssd1 vccd1 vccd1
+ _12454_/A sky130_fd_sc_hd__o2111ai_4
XFILLER_114_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14028_ _19176_/Q _14043_/A2 _14040_/B1 _14027_/X _16127_/B1 vssd1 vssd1 vccd1 vccd1
+ _19176_/D sky130_fd_sc_hd__o221a_1
X_18905_ _18905_/A _18905_/B vssd1 vssd1 vccd1 vccd1 _21000_/D sky130_fd_sc_hd__nor2_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19885_ _20708_/CLK _19885_/D vssd1 vssd1 vccd1 vccd1 _19885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_206_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18836_ _19095_/Q _12589_/B _12590_/Y _13459_/Y vssd1 vssd1 vccd1 vccd1 _18837_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_256_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18767_ _18767_/A _18767_/B vssd1 vssd1 vccd1 vccd1 _18767_/X sky130_fd_sc_hd__or2_1
XFILLER_83_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15979_ _15979_/A _15979_/B _15814_/A vssd1 vssd1 vccd1 vccd1 _15979_/X sky130_fd_sc_hd__or3b_2
XFILLER_243_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17718_ _20499_/Q _17892_/A1 _17742_/S vssd1 vssd1 vccd1 vccd1 _20499_/D sky130_fd_sc_hd__mux2_1
XFILLER_209_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18698_ _18698_/A _18698_/B vssd1 vssd1 vccd1 vccd1 _20949_/D sky130_fd_sc_hd__and2_1
XFILLER_35_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17649_ _20435_/Q _17649_/A1 _17657_/S vssd1 vssd1 vccd1 vccd1 _20435_/D sky130_fd_sc_hd__mux2_1
XFILLER_243_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20660_ _20660_/CLK _20660_/D vssd1 vssd1 vccd1 vccd1 _20660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_189_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19523_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19319_ _20646_/CLK _19319_/D vssd1 vssd1 vccd1 vccd1 _19319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20591_ _20686_/CLK _20591_/D vssd1 vssd1 vccd1 vccd1 _20591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_118_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20949_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout501 _17813_/X vssd1 vssd1 vccd1 vccd1 _17840_/S sky130_fd_sc_hd__buf_4
X_09905_ _12157_/A1 _09936_/A2 _09904_/X _12153_/B1 vssd1 vssd1 vccd1 vccd1 _13726_/A
+ sky130_fd_sc_hd__o211ai_4
Xfanout512 _17711_/X vssd1 vssd1 vccd1 vccd1 _17740_/S sky130_fd_sc_hd__buf_12
Xfanout523 _17642_/X vssd1 vssd1 vccd1 vccd1 _17657_/S sky130_fd_sc_hd__buf_12
XFILLER_116_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout534 _17570_/S vssd1 vssd1 vccd1 vccd1 _17572_/S sky130_fd_sc_hd__buf_12
XFILLER_86_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout545 _17132_/S vssd1 vssd1 vccd1 vccd1 _17149_/S sky130_fd_sc_hd__buf_12
XFILLER_116_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout556 _16673_/X vssd1 vssd1 vccd1 vccd1 _16702_/S sky130_fd_sc_hd__buf_12
X_20025_ _20660_/CLK _20025_/D vssd1 vssd1 vccd1 vccd1 _20025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_274_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout567 _16605_/X vssd1 vssd1 vccd1 vccd1 _16620_/S sky130_fd_sc_hd__buf_12
XFILLER_100_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09836_ _20419_/Q _20355_/Q _20647_/Q _20611_/Q _10092_/S _12084_/C vssd1 vssd1 vccd1
+ vccd1 _09836_/X sky130_fd_sc_hd__mux4_1
XFILLER_247_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout578 _16272_/S vssd1 vssd1 vccd1 vccd1 _16275_/S sky130_fd_sc_hd__buf_12
XFILLER_258_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout589 _14774_/A2 vssd1 vssd1 vccd1 vccd1 _14764_/A2 sky130_fd_sc_hd__buf_4
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09767_ _20324_/Q _11936_/S _09766_/X vssd1 vssd1 vccd1 vccd1 _09767_/X sky130_fd_sc_hd__a21o_1
XFILLER_273_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09698_ _20484_/Q _20324_/Q _11889_/S vssd1 vssd1 vccd1 vccd1 _09698_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20927_ _21025_/CLK _20927_/D vssd1 vssd1 vccd1 vccd1 _20927_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _20479_/Q _20319_/Q _12053_/S vssd1 vssd1 vccd1 vccd1 _11660_/X sky130_fd_sc_hd__mux2_1
X_20858_ _21018_/CLK _20858_/D vssd1 vssd1 vccd1 vccd1 _20858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10611_ _20342_/Q _10611_/B _11693_/B vssd1 vssd1 vccd1 vccd1 _10611_/X sky130_fd_sc_hd__or3_1
XFILLER_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ _11576_/X _11577_/X _11980_/S vssd1 vssd1 vccd1 vccd1 _11591_/X sky130_fd_sc_hd__mux2_1
X_20789_ _20856_/CLK _20789_/D vssd1 vssd1 vccd1 vccd1 _20789_/Q sky130_fd_sc_hd__dfxtp_1
X_13330_ _13325_/X _13329_/X _14295_/C1 vssd1 vssd1 vccd1 vccd1 _13330_/X sky130_fd_sc_hd__a21o_1
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10542_ _10641_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _13611_/A sky130_fd_sc_hd__xnor2_4
XFILLER_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13261_ _13397_/B _13258_/X _13259_/Y _13260_/Y _18651_/B vssd1 vssd1 vccd1 vccd1
+ _13261_/X sky130_fd_sc_hd__o311a_2
X_10473_ _10561_/A _10472_/X _10457_/Y vssd1 vssd1 vccd1 vccd1 _10473_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ _20554_/Q _12316_/S vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__or2_1
X_15000_ _15308_/B _14997_/C _14972_/B _14991_/X vssd1 vssd1 vccd1 vccd1 _15000_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_136_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13192_ _13192_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13192_/Y sky130_fd_sc_hd__nor2_8
XFILLER_194_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12143_ _12141_/X _12142_/X _12143_/S vssd1 vssd1 vccd1 vccd1 _12143_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_4__f_wb_clk_i clkbuf_3_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_4__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_269_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16951_ input59/X input94/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16951_/X sky130_fd_sc_hd__mux2_8
XFILLER_1_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12074_ _12059_/X _12073_/X _12074_/B1 vssd1 vssd1 vccd1 vccd1 _12074_/X sky130_fd_sc_hd__a21o_2
XFILLER_278_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11025_ _11026_/A _20496_/Q _10345_/S _20528_/Q vssd1 vssd1 vccd1 vccd1 _11025_/X
+ sky130_fd_sc_hd__o22a_1
X_15902_ _13432_/A _16054_/B _15900_/X _15901_/X vssd1 vssd1 vccd1 vccd1 _15903_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19670_ _20559_/CLK _19670_/D vssd1 vssd1 vccd1 vccd1 _19670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16882_ _16878_/Y _16879_/X _16881_/X _16932_/A1 vssd1 vssd1 vccd1 vccd1 _16882_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18621_ _18508_/X _18621_/A2 _18619_/Y _18620_/Y vssd1 vssd1 vccd1 vccd1 _18622_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15833_ _19757_/Q _15999_/A2 _15832_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15833_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _18960_/A _18552_/B vssd1 vssd1 vccd1 vccd1 _20910_/D sky130_fd_sc_hd__nor2_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _09940_/Y _15984_/A2 _15984_/B1 _09941_/A _15890_/A vssd1 vssd1 vccd1 vccd1
+ _15764_/X sky130_fd_sc_hd__a221o_2
X_12976_ _12976_/A _12976_/B vssd1 vssd1 vccd1 vccd1 _12976_/Y sky130_fd_sc_hd__nor2_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17505_/A1 _17502_/Y _18980_/A vssd1 vssd1 vccd1 vccd1 _20286_/D sky130_fd_sc_hd__a21oi_1
X_14715_ _19472_/Q _17930_/A1 _14719_/S vssd1 vssd1 vccd1 vccd1 _19472_/D sky130_fd_sc_hd__mux2_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18483_ _18570_/B _18483_/B vssd1 vssd1 vccd1 vccd1 _18483_/X sky130_fd_sc_hd__or2_2
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _19648_/Q _19954_/Q _19292_/Q _20079_/Q _09931_/S _09986_/C vssd1 vssd1 vccd1
+ vccd1 _11927_/X sky130_fd_sc_hd__mux4_1
X_15695_ _16046_/A1 _15694_/X _15690_/X vssd1 vssd1 vccd1 vccd1 _15695_/X sky130_fd_sc_hd__o21a_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_450 _13775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_461 _19245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_472 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17434_ _17434_/A _17434_/B vssd1 vssd1 vccd1 vccd1 _20261_/D sky130_fd_sc_hd__and2_1
XFILLER_260_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_483 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14646_ _19408_/Q _17930_/A1 _14650_/S vssd1 vssd1 vccd1 vccd1 _19408_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_494 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11858_ _11856_/X _11857_/X _12006_/S vssd1 vssd1 vccd1 vccd1 _11858_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_19 _15535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ input162/X input137/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__mux2_8
XFILLER_202_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17365_ _20231_/Q _17371_/A2 _17364_/X _18702_/A vssd1 vssd1 vccd1 vccd1 _20231_/D
+ sky130_fd_sc_hd__o211a_1
X_14577_ _19343_/Q _17929_/A1 _14594_/S vssd1 vssd1 vccd1 vccd1 _19343_/D sky130_fd_sc_hd__mux2_1
X_11789_ _15433_/A _15433_/B _11768_/X _11773_/X _11788_/X vssd1 vssd1 vccd1 vccd1
+ _11789_/X sky130_fd_sc_hd__a2111o_1
Xclkbuf_leaf_211_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20682_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_19104_ _19511_/CLK _19104_/D vssd1 vssd1 vccd1 vccd1 _19104_/Q sky130_fd_sc_hd__dfxtp_4
X_16316_ _19714_/Q _16316_/B vssd1 vssd1 vccd1 vccd1 _16322_/C sky130_fd_sc_hd__and2_2
XFILLER_203_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13528_ _19219_/Q _19218_/Q _13498_/B _19220_/Q vssd1 vssd1 vccd1 vccd1 _13529_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17296_ _17296_/A _17329_/S _17305_/C vssd1 vssd1 vccd1 vccd1 _17296_/X sky130_fd_sc_hd__and3_1
XFILLER_201_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19035_ _21036_/Q _19049_/A2 _19034_/X _18734_/A vssd1 vssd1 vccd1 vccd1 _21036_/D
+ sky130_fd_sc_hd__o211a_1
X_16247_ _19663_/Q _17921_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19663_/D sky130_fd_sc_hd__mux2_1
XFILLER_173_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13459_ _13459_/A _13459_/B vssd1 vssd1 vccd1 vccd1 _13459_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_284_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16178_ _19613_/Q _15807_/X _16178_/S vssd1 vssd1 vccd1 vccd1 _16179_/B sky130_fd_sc_hd__mux2_1
XFILLER_217_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15129_ _15129_/A0 _12668_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _15129_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19937_ _20633_/CLK _19937_/D vssd1 vssd1 vccd1 vccd1 _19937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19868_ _20565_/CLK _19868_/D vssd1 vssd1 vccd1 vccd1 _19868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09621_ _09621_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09621_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18819_ _20988_/Q _18819_/B vssd1 vssd1 vccd1 vccd1 _18819_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19799_ _20670_/CLK _19799_/D vssd1 vssd1 vccd1 vccd1 _19799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09552_ _12468_/C _09552_/B vssd1 vssd1 vccd1 vccd1 _13635_/A sky130_fd_sc_hd__nor2_2
XFILLER_271_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09483_ _20298_/Q vssd1 vssd1 vccd1 vccd1 _17526_/C sky130_fd_sc_hd__inv_2
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20712_ _20712_/CLK _20712_/D vssd1 vssd1 vccd1 vccd1 _20712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20643_ _20675_/CLK _20643_/D vssd1 vssd1 vccd1 vccd1 _20643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20574_ _20574_/CLK _20574_/D vssd1 vssd1 vccd1 vccd1 _20574_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20273_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1307 _12962_/S vssd1 vssd1 vccd1 vccd1 _12950_/B2 sky130_fd_sc_hd__buf_4
XFILLER_132_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20472_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1318 _14878_/B vssd1 vssd1 vccd1 vccd1 _16057_/A2 sky130_fd_sc_hd__buf_2
Xfanout1329 _16030_/D1 vssd1 vssd1 vccd1 vccd1 _12579_/D sky130_fd_sc_hd__buf_6
XFILLER_132_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20008_ _20751_/CLK _20008_/D vssd1 vssd1 vccd1 vccd1 _20008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09819_ _20044_/Q _19919_/Q _10426_/S vssd1 vssd1 vccd1 vccd1 _09819_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_274_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12830_ _12829_/B _12829_/C _12829_/D _12839_/A vssd1 vssd1 vccd1 vccd1 _12864_/B
+ sky130_fd_sc_hd__o22ai_4
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_227_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12759_/X _12771_/B vssd1 vssd1 vccd1 vccd1 _13448_/A sky130_fd_sc_hd__and2b_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _19278_/Q _17095_/A1 _14516_/S vssd1 vssd1 vccd1 vccd1 _19278_/D sky130_fd_sc_hd__mux2_1
XFILLER_230_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _12102_/A1 _19480_/Q _19448_/Q _12025_/S vssd1 vssd1 vccd1 vccd1 _11712_/X
+ sky130_fd_sc_hd__a22o_1
X_12692_ _12693_/A _13526_/A _12692_/C _12692_/D vssd1 vssd1 vccd1 vccd1 _12699_/B
+ sky130_fd_sc_hd__or4_1
X_15480_ _20957_/Q _15568_/A2 _15568_/B1 _20829_/Q _15479_/X vssd1 vssd1 vccd1 vccd1
+ _15480_/X sky130_fd_sc_hd__a221o_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14431_ _20297_/Q _14431_/A2 _14431_/B1 input239/X vssd1 vssd1 vccd1 vccd1 _14435_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11872_/A _12006_/S _11642_/X _12012_/S vssd1 vssd1 vccd1 vccd1 _11643_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17150_ _17744_/A _17184_/A vssd1 vssd1 vccd1 vccd1 _17151_/C sky130_fd_sc_hd__nor2_1
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14362_ _20290_/Q _14431_/A2 _14431_/B1 input231/X vssd1 vssd1 vccd1 vccd1 _14364_/B
+ sky130_fd_sc_hd__a22o_2
X_11574_ _11574_/A _11735_/B vssd1 vssd1 vccd1 vccd1 _11575_/B sky130_fd_sc_hd__and2_2
XFILLER_155_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 core_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_4
X_16101_ _19575_/Q _16127_/A2 _16107_/B1 vssd1 vssd1 vccd1 vccd1 _16101_/X sky130_fd_sc_hd__o21a_1
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 core_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10525_ _10516_/X _10524_/X _10525_/S vssd1 vssd1 vccd1 vccd1 _10525_/X sky130_fd_sc_hd__mux2_2
Xinput39 core_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_4
X_13313_ _20926_/Q _13602_/A1 _13311_/X _13312_/Y _18612_/B vssd1 vssd1 vccd1 vccd1
+ _13313_/X sky130_fd_sc_hd__a221o_1
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17081_ _20053_/Q _17674_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20053_/D sky130_fd_sc_hd__mux2_1
X_14293_ _14293_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14293_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_182_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16032_ _15544_/A _16024_/X _16031_/X vssd1 vssd1 vccd1 vccd1 _16032_/X sky130_fd_sc_hd__o21a_1
X_13244_ _13245_/A _13245_/B vssd1 vssd1 vccd1 vccd1 _13244_/X sky130_fd_sc_hd__and2_4
XFILLER_171_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ _10456_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10456_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13175_ _12034_/Y _13431_/B _12036_/B vssd1 vssd1 vccd1 vccd1 _13183_/B sky130_fd_sc_hd__o21a_4
XFILLER_272_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10387_ _19876_/Q _10400_/S vssd1 vssd1 vccd1 vccd1 _10387_/X sky130_fd_sc_hd__or2_1
XFILLER_272_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _19690_/Q _20178_/Q _12133_/S vssd1 vssd1 vccd1 vccd1 _12126_/X sky130_fd_sc_hd__mux2_1
X_17983_ _20732_/Q _17985_/C _18416_/A vssd1 vssd1 vccd1 vccd1 _17984_/B sky130_fd_sc_hd__o21ai_1
XFILLER_96_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19722_ _21026_/CLK _19722_/D vssd1 vssd1 vccd1 vccd1 _19722_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1830 _19174_/Q vssd1 vssd1 vccd1 vccd1 _11670_/S sky130_fd_sc_hd__buf_12
X_16934_ _16885_/A _16933_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16934_/Y sky130_fd_sc_hd__o21bai_4
X_12057_ _10430_/S _12050_/X _12051_/X vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__o21a_1
Xfanout1841 _10057_/S vssd1 vssd1 vccd1 vccd1 _10430_/S sky130_fd_sc_hd__buf_6
Xfanout1852 _19170_/Q vssd1 vssd1 vccd1 vccd1 _11281_/A sky130_fd_sc_hd__buf_12
X_11008_ _11008_/A1 _19305_/Q _11008_/A3 _10235_/S vssd1 vssd1 vccd1 vccd1 _11008_/X
+ sky130_fd_sc_hd__o31a_1
Xfanout1863 _15678_/A1 vssd1 vssd1 vccd1 vccd1 _12850_/A1 sky130_fd_sc_hd__buf_12
X_19653_ _20463_/CLK _19653_/D vssd1 vssd1 vccd1 vccd1 _19653_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1874 _09731_/A vssd1 vssd1 vccd1 vccd1 _12429_/A1 sky130_fd_sc_hd__buf_6
XFILLER_78_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1885 _19097_/Q vssd1 vssd1 vccd1 vccd1 _12967_/B sky130_fd_sc_hd__buf_8
X_16865_ _16884_/S _09527_/Y _16809_/X _16864_/Y vssd1 vssd1 vccd1 vccd1 _16865_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_65_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1896 _18736_/A vssd1 vssd1 vccd1 vccd1 _18734_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_253_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18604_ _19504_/Q _18604_/B vssd1 vssd1 vccd1 vccd1 _18604_/Y sky130_fd_sc_hd__nand2_1
XFILLER_219_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15816_ _15816_/A _15925_/B vssd1 vssd1 vccd1 vccd1 _15816_/Y sky130_fd_sc_hd__nand2_1
XFILLER_281_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19584_ _20665_/CLK _19584_/D vssd1 vssd1 vccd1 vccd1 _19584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16796_ _19091_/Q _16996_/B1 _16795_/X vssd1 vssd1 vccd1 vccd1 _16796_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18535_ _18651_/B _18535_/B vssd1 vssd1 vccd1 vccd1 _18535_/X sky130_fd_sc_hd__or2_2
XFILLER_206_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _20902_/Q _16043_/A2 _16043_/B1 _15746_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _15747_/X sky130_fd_sc_hd__a221o_1
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12959_ _16719_/B _12959_/B vssd1 vssd1 vccd1 vccd1 _16710_/A sky130_fd_sc_hd__or2_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18466_ _18570_/B _18466_/B vssd1 vssd1 vccd1 vccd1 _18467_/B sky130_fd_sc_hd__or2_1
XFILLER_233_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15678_ _15678_/A1 _12581_/B _16007_/A vssd1 vssd1 vccd1 vccd1 _15678_/X sky130_fd_sc_hd__a21bo_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 _20623_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_291 input222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17417_ _17402_/Y _17416_/X _17415_/X _17434_/A vssd1 vssd1 vccd1 vccd1 _20254_/D
+ sky130_fd_sc_hd__o211a_1
X_14629_ _19393_/Q _17913_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19393_/D sky130_fd_sc_hd__mux2_1
X_18397_ _20853_/Q _18175_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18398_/B sky130_fd_sc_hd__mux2_1
XFILLER_159_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ _20222_/Q _17356_/A2 _17362_/B1 _20271_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17348_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17279_ _20198_/Q _17330_/A2 _17290_/C _17278_/Y _17279_/C1 vssd1 vssd1 vccd1 vccd1
+ _17279_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19018_ _18240_/Y _19048_/A2 _19017_/X _12551_/C _19048_/C1 vssd1 vssd1 vccd1 vccd1
+ _19018_/X sky130_fd_sc_hd__a221o_1
X_20290_ _20296_/CLK _20290_/D vssd1 vssd1 vccd1 vccd1 _20290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_0_0_wb_clk_i ANTENNA_548/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_114_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09604_ _09604_/A _17850_/A _17884_/A vssd1 vssd1 vccd1 vccd1 _09607_/B sky130_fd_sc_hd__or3_2
XFILLER_249_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09535_ _19155_/Q _13869_/A vssd1 vssd1 vccd1 vccd1 _09555_/C sky130_fd_sc_hd__nand2_2
XFILLER_83_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_133_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _20980_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20626_ _20659_/CLK _20626_/D vssd1 vssd1 vccd1 vccd1 _20626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20557_ _20557_/CLK _20557_/D vssd1 vssd1 vccd1 vccd1 _20557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ _11101_/A _10308_/X _10309_/X _12311_/C1 vssd1 vssd1 vccd1 vccd1 _10310_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_138_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11290_ _11290_/A _20657_/Q _11290_/C vssd1 vssd1 vccd1 vccd1 _11290_/X sky130_fd_sc_hd__or3_1
XFILLER_164_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20488_ _20716_/CLK _20488_/D vssd1 vssd1 vccd1 vccd1 _20488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10241_ _11012_/A _10240_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _10241_/X sky130_fd_sc_hd__o21a_1
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10172_ _10168_/X _10171_/X _11375_/S vssd1 vssd1 vccd1 vccd1 _10172_/X sky130_fd_sc_hd__mux2_1
Xfanout1104 _17111_/A1 vssd1 vssd1 vccd1 vccd1 _17947_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1115 _11807_/X vssd1 vssd1 vccd1 vccd1 _17876_/A1 sky130_fd_sc_hd__buf_4
Xfanout1126 _17936_/A1 vssd1 vssd1 vccd1 vccd1 _17902_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_266_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14980_ _15314_/B _14980_/B _14980_/C vssd1 vssd1 vccd1 vccd1 _14980_/X sky130_fd_sc_hd__or3_1
Xfanout1137 _09947_/X vssd1 vssd1 vccd1 vccd1 _17940_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_266_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1148 _09790_/X vssd1 vssd1 vccd1 vccd1 _17908_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1159 _09631_/X vssd1 vssd1 vccd1 vccd1 _11012_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13931_ _19135_/Q _13943_/S _13932_/B1 _13361_/C vssd1 vssd1 vccd1 vccd1 _19135_/D
+ sky130_fd_sc_hd__o22a_1
Xwire1254 _13468_/Y vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__buf_12
XFILLER_86_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ _19907_/Q _17060_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19907_/D sky130_fd_sc_hd__mux2_1
X_13862_ _16133_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _13862_/X sky130_fd_sc_hd__and2_4
XFILLER_75_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15601_ _20865_/Q _15600_/X _15601_/S vssd1 vssd1 vccd1 vccd1 _15601_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12813_ _19514_/Q _12916_/A2 _12812_/X _12916_/B2 vssd1 vssd1 vccd1 vccd1 _12815_/B
+ sky130_fd_sc_hd__o22a_4
X_16581_ _16591_/A _16581_/B vssd1 vssd1 vccd1 vccd1 _19856_/D sky130_fd_sc_hd__or2_1
XFILLER_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13793_ _13798_/A1 _13826_/A1 _13676_/B _13826_/B1 input237/X vssd1 vssd1 vccd1 vccd1
+ _13793_/X sky130_fd_sc_hd__a32o_1
XFILLER_262_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18320_ _18320_/A _18457_/B vssd1 vssd1 vccd1 vccd1 _18981_/C sky130_fd_sc_hd__or2_4
XFILLER_27_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ _21025_/Q _20993_/Q _15993_/S vssd1 vssd1 vccd1 vccd1 _15532_/X sky130_fd_sc_hd__mux2_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _19507_/Q _12744_/B vssd1 vssd1 vccd1 vccd1 _12747_/B sky130_fd_sc_hd__or2_4
XFILLER_215_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _20804_/Q _18250_/Y _18316_/S vssd1 vssd1 vccd1 vccd1 _18252_/B sky130_fd_sc_hd__mux2_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15463_ _11764_/Y _11765_/X _15127_/B vssd1 vssd1 vccd1 vccd1 _15465_/A sky130_fd_sc_hd__a21o_1
X_12675_ _12675_/A _12675_/B _12675_/C vssd1 vssd1 vccd1 vccd1 _12676_/B sky130_fd_sc_hd__and3_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17202_ _20166_/Q _17202_/A1 _17214_/S vssd1 vssd1 vccd1 vccd1 _20166_/D sky130_fd_sc_hd__mux2_1
X_14414_ _14426_/A _14424_/A vssd1 vssd1 vccd1 vccd1 _14416_/A sky130_fd_sc_hd__or2_1
X_18182_ _18708_/A _18182_/B vssd1 vssd1 vccd1 vccd1 _20790_/D sky130_fd_sc_hd__and2_1
X_11626_ _11624_/X _11625_/X _11641_/S vssd1 vssd1 vccd1 vccd1 _11626_/X sky130_fd_sc_hd__mux2_1
X_15394_ _19742_/Q _15453_/A2 _15382_/X _15021_/A _15393_/X vssd1 vssd1 vccd1 vccd1
+ _15394_/X sky130_fd_sc_hd__a221o_1
X_17133_ _20101_/Q _17692_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20101_/D sky130_fd_sc_hd__mux2_1
X_14345_ _14427_/A _14345_/B _14354_/B vssd1 vssd1 vccd1 vccd1 _14345_/X sky130_fd_sc_hd__or3b_1
X_11557_ _12008_/A _19478_/Q _19446_/Q _09931_/S vssd1 vssd1 vccd1 vccd1 _11557_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17064_ _20036_/Q _17934_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20036_/D sky130_fd_sc_hd__mux2_1
X_10508_ _10540_/A _10540_/B vssd1 vssd1 vccd1 vccd1 _10641_/A sky130_fd_sc_hd__nand2_4
XFILLER_170_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11488_ _20135_/Q _20103_/Q _12174_/S vssd1 vssd1 vccd1 vccd1 _11488_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14276_ _14397_/A _14397_/B _14276_/C vssd1 vssd1 vccd1 vccd1 _14276_/X sky130_fd_sc_hd__or3_1
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16015_ _20944_/Q _16044_/A2 _16014_/X vssd1 vssd1 vccd1 vccd1 _16015_/X sky130_fd_sc_hd__o21a_1
X_13227_ _13227_/A _13272_/B vssd1 vssd1 vccd1 vccd1 _13227_/Y sky130_fd_sc_hd__nor2_1
X_10439_ _11281_/A _20065_/Q _11268_/C vssd1 vssd1 vccd1 vccd1 _10439_/X sky130_fd_sc_hd__and3_1
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _10198_/A _13424_/B _15549_/S vssd1 vssd1 vccd1 vccd1 _13423_/B sky130_fd_sc_hd__a21bo_4
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12110_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12109_/Y sky130_fd_sc_hd__nor2_2
X_17966_ _18056_/A _17971_/C vssd1 vssd1 vccd1 vccd1 _17966_/Y sky130_fd_sc_hd__nor2_1
XFILLER_239_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13089_ _13009_/Y _13121_/A _13120_/B vssd1 vssd1 vccd1 vccd1 _13135_/A sky130_fd_sc_hd__o21a_1
XFILLER_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_273_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19705_ _20759_/CLK _19705_/D vssd1 vssd1 vccd1 vccd1 _19705_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1660 _09646_/Y vssd1 vssd1 vccd1 vccd1 _14038_/A2 sky130_fd_sc_hd__buf_4
X_16917_ input55/X input90/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16917_/X sky130_fd_sc_hd__mux2_8
XFILLER_66_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1671 _14002_/A1 vssd1 vssd1 vccd1 vccd1 _14029_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_111_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17897_ _20668_/Q split4/X _17912_/S vssd1 vssd1 vccd1 vccd1 _20668_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1682 _12008_/A vssd1 vssd1 vccd1 vccd1 _11851_/A sky130_fd_sc_hd__buf_6
XFILLER_226_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1693 _10937_/A vssd1 vssd1 vccd1 vccd1 _11021_/A sky130_fd_sc_hd__buf_6
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19636_ _20633_/CLK _19636_/D vssd1 vssd1 vccd1 vccd1 _19636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16848_ _16932_/B1 _16845_/X _16847_/X _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16849_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_265_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19567_ _19577_/CLK _19567_/D vssd1 vssd1 vccd1 vccd1 _19567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16779_ input98/X input73/X _16799_/S vssd1 vssd1 vccd1 vccd1 _16780_/A sky130_fd_sc_hd__mux2_2
XFILLER_241_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18518_ _20899_/Q _18559_/B _18517_/X _18458_/B vssd1 vssd1 vccd1 vccd1 _18519_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_222_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19498_ _21023_/CLK _19498_/D vssd1 vssd1 vccd1 vccd1 _19498_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18449_ _20879_/Q _18305_/Y _18449_/S vssd1 vssd1 vccd1 vccd1 _18450_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20411_ _20635_/CLK _20411_/D vssd1 vssd1 vccd1 vccd1 _20411_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_175_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20342_ _20666_/CLK _20342_/D vssd1 vssd1 vccd1 vccd1 _20342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20273_ _20273_/CLK _20273_/D vssd1 vssd1 vccd1 vccd1 _20273_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_89_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_276_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput207 localMemory_wb_adr_i[3] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__clkbuf_2
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput218 localMemory_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_hd__buf_12
Xinput229 localMemory_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__buf_12
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ input43/X vssd1 vssd1 vccd1 vccd1 _09518_/Y sky130_fd_sc_hd__inv_2
X_10790_ _19404_/Q _20563_/Q _11126_/B vssd1 vssd1 vccd1 vccd1 _10790_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12460_ _12449_/A _12450_/A _12445_/B _12447_/B vssd1 vssd1 vccd1 vccd1 _12463_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _10197_/A _11411_/B vssd1 vssd1 vccd1 vccd1 _11411_/X sky130_fd_sc_hd__and2b_1
X_12391_ _12389_/X _12390_/X _12391_/S vssd1 vssd1 vccd1 vccd1 _12391_/X sky130_fd_sc_hd__mux2_1
X_20609_ _20681_/CLK _20609_/D vssd1 vssd1 vccd1 vccd1 _20609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11342_ _20126_/Q _20094_/Q _11342_/S vssd1 vssd1 vccd1 vccd1 _11342_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14130_ _19495_/Q _14130_/B vssd1 vssd1 vccd1 vccd1 _14131_/B sky130_fd_sc_hd__xor2_4
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20465_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14061_ _14081_/A _14069_/B _14061_/C vssd1 vssd1 vccd1 vccd1 _14061_/X sky130_fd_sc_hd__or3_1
X_11273_ _11273_/A1 _19302_/Q _09623_/B _10322_/S vssd1 vssd1 vccd1 vccd1 _11273_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_141_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10224_ _20037_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _10224_/X sky130_fd_sc_hd__or2_1
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13012_ _20973_/Q _20907_/Q vssd1 vssd1 vccd1 vccd1 _13012_/X sky130_fd_sc_hd__or2_1
XFILLER_279_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17820_ _20595_/Q _17892_/A1 _17844_/S vssd1 vssd1 vccd1 vccd1 _20595_/D sky130_fd_sc_hd__mux2_1
X_10155_ _19811_/Q _19315_/Q _12296_/S vssd1 vssd1 vccd1 vccd1 _10155_/X sky130_fd_sc_hd__mux2_1
X_17751_ _20530_/Q _17751_/A1 _17776_/S vssd1 vssd1 vccd1 vccd1 _20530_/D sky130_fd_sc_hd__mux2_1
XFILLER_254_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14963_ _14983_/A _15020_/A vssd1 vssd1 vccd1 vccd1 _14963_/Y sky130_fd_sc_hd__nor2_1
X_10086_ _10083_/X _10085_/X _12514_/C vssd1 vssd1 vccd1 vccd1 _10086_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16702_ _19957_/Q _17705_/A1 _16702_/S vssd1 vssd1 vccd1 vccd1 _19957_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13914_ _19122_/Q _13919_/S _13913_/Y _18710_/A vssd1 vssd1 vccd1 vccd1 _19122_/D
+ sky130_fd_sc_hd__o211a_1
X_17682_ _20466_/Q _17857_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20466_/D sky130_fd_sc_hd__mux2_1
XFILLER_247_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14894_ _14894_/A _14897_/B vssd1 vssd1 vccd1 vccd1 _16037_/B sky130_fd_sc_hd__nor2_4
XFILLER_235_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19421_ _20580_/CLK _19421_/D vssd1 vssd1 vccd1 vccd1 _19421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_236_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16633_ _19892_/Q _17947_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19892_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13845_ _20260_/Q _20259_/Q _20257_/Q vssd1 vssd1 vccd1 vccd1 _13846_/C sky130_fd_sc_hd__or3b_2
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19352_ _20715_/CLK _19352_/D vssd1 vssd1 vccd1 vccd1 _19352_/Q sky130_fd_sc_hd__dfxtp_1
X_16564_ _19848_/Q _16576_/A2 _16576_/B1 input18/X vssd1 vssd1 vccd1 vccd1 _16565_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_216_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13776_ _12328_/Y _13730_/B _13776_/B1 vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__o21a_2
X_10988_ _11336_/A _11008_/A1 _19337_/Q _12377_/S vssd1 vssd1 vccd1 vccd1 _10988_/X
+ sky130_fd_sc_hd__a31o_1
X_18303_ _19556_/Q _18313_/B vssd1 vssd1 vccd1 vccd1 _18303_/Y sky130_fd_sc_hd__nand2b_2
X_15515_ _19746_/Q _15604_/A2 _15514_/X _16048_/C1 vssd1 vssd1 vccd1 vccd1 _15515_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_200_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19283_ _20573_/CLK _19283_/D vssd1 vssd1 vccd1 vccd1 _19283_/Q sky130_fd_sc_hd__dfxtp_1
X_12727_ _12468_/B _12832_/B split6/A _12710_/B vssd1 vssd1 vccd1 vccd1 _12736_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_200_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16495_ _19802_/Q _17890_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19802_/D sky130_fd_sc_hd__mux2_1
XFILLER_70_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18234_ _18248_/B _14269_/B _18233_/Y vssd1 vssd1 vccd1 vccd1 _18511_/B sky130_fd_sc_hd__o21ai_4
X_15446_ _21022_/Q _20990_/Q _15508_/S vssd1 vssd1 vccd1 vccd1 _15446_/X sky130_fd_sc_hd__mux2_1
X_12658_ _12658_/A _12784_/B vssd1 vssd1 vccd1 vccd1 _12658_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18165_ _18463_/B vssd1 vssd1 vccd1 vccd1 _18165_/Y sky130_fd_sc_hd__inv_2
X_11609_ _11594_/X _11608_/X _12153_/A1 vssd1 vssd1 vccd1 vccd1 _11609_/X sky130_fd_sc_hd__a21o_1
X_15377_ _15258_/A _15373_/X _15376_/Y _14843_/S vssd1 vssd1 vccd1 vccd1 _15377_/X
+ sky130_fd_sc_hd__o22a_1
X_12589_ _12589_/A _12589_/B _12589_/C vssd1 vssd1 vccd1 vccd1 _12592_/B sky130_fd_sc_hd__or3_1
XFILLER_144_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17116_ _17918_/A _17184_/A vssd1 vssd1 vccd1 vccd1 _17117_/C sky130_fd_sc_hd__nor2_1
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14328_ _14397_/A _14437_/B _14328_/C vssd1 vssd1 vccd1 vccd1 _14328_/X sky130_fd_sc_hd__or3_1
XFILLER_209_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18096_ _18096_/A _18101_/C vssd1 vssd1 vccd1 vccd1 _18096_/Y sky130_fd_sc_hd__nor2_1
XFILLER_209_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17047_ _20020_/Q _16706_/X _17046_/X vssd1 vssd1 vccd1 vccd1 _20021_/D sky130_fd_sc_hd__a21oi_1
XFILLER_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14259_ _19508_/Q _14259_/B vssd1 vssd1 vccd1 vccd1 _14260_/C sky130_fd_sc_hd__xnor2_1
XFILLER_143_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 _14996_/X vssd1 vssd1 vccd1 vccd1 _16042_/A2 sky130_fd_sc_hd__buf_4
Xfanout919 _16011_/A2 vssd1 vssd1 vccd1 vccd1 _16041_/A2 sky130_fd_sc_hd__buf_8
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18998_ _18190_/Y _18983_/B _19002_/B1 _18997_/X vssd1 vssd1 vccd1 vccd1 _21018_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _20718_/Q _17949_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20718_/D sky130_fd_sc_hd__mux2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1490 _09728_/X vssd1 vssd1 vccd1 vccd1 _09839_/A sky130_fd_sc_hd__buf_12
XFILLER_66_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20960_ _21024_/CLK _20960_/D vssd1 vssd1 vccd1 vccd1 _20960_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_238_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_285_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19619_ _20263_/CLK _19619_/D vssd1 vssd1 vccd1 vccd1 _19619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20891_ _21023_/CLK _20891_/D vssd1 vssd1 vccd1 vccd1 _20891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20325_ _21046_/A _20325_/D vssd1 vssd1 vccd1 vccd1 _20325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20256_ _20261_/CLK _20256_/D vssd1 vssd1 vccd1 vccd1 _20256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_249_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20187_ _20688_/CLK _20187_/D vssd1 vssd1 vccd1 vccd1 _20187_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09998_ _12015_/A1 _09996_/X _09997_/X vssd1 vssd1 vccd1 vccd1 _09998_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_103_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11960_ _13433_/A _11960_/B vssd1 vssd1 vccd1 vccd1 _12290_/A sky130_fd_sc_hd__xnor2_2
XFILLER_229_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10911_ _19402_/Q _12296_/S vssd1 vssd1 vccd1 vccd1 _10911_/X sky130_fd_sc_hd__or2_1
XFILLER_218_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _19423_/Q _11891_/B vssd1 vssd1 vccd1 vccd1 _11891_/X sky130_fd_sc_hd__or2_1
XFILLER_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _13478_/B _13220_/Y _15949_/B _13765_/A vssd1 vssd1 vccd1 vccd1 _13630_/X
+ sky130_fd_sc_hd__a22o_4
X_10842_ _20027_/Q _19902_/Q _10842_/S vssd1 vssd1 vccd1 vccd1 _10842_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13561_ _12652_/B _13558_/Y _13560_/X vssd1 vssd1 vccd1 vccd1 _13561_/Y sky130_fd_sc_hd__a21oi_2
X_10773_ _12337_/A _20663_/Q _12254_/C vssd1 vssd1 vccd1 vccd1 _10773_/X sky130_fd_sc_hd__or3_1
XFILLER_197_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15300_ _13150_/A _14878_/B _15299_/X vssd1 vssd1 vccd1 vccd1 _15326_/B sky130_fd_sc_hd__a21oi_1
XFILLER_197_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ _13897_/A _12512_/B _12517_/C _12584_/B vssd1 vssd1 vccd1 vccd1 _12515_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_185_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16280_ _20621_/Q _17015_/B _19701_/D vssd1 vssd1 vccd1 vccd1 _19696_/D sky130_fd_sc_hd__and3_1
X_13492_ _12584_/A _19217_/Q _13491_/X vssd1 vssd1 vccd1 vccd1 _13907_/A sky130_fd_sc_hd__a21oi_4
XFILLER_200_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15231_ _20726_/Q _15445_/A2 _15445_/B1 _20758_/Q vssd1 vssd1 vccd1 vccd1 _15231_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ _12436_/A _12443_/B vssd1 vssd1 vccd1 vccd1 _12444_/B sky130_fd_sc_hd__nand2b_1
XFILLER_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15162_ _15161_/Y _15159_/Y _15357_/S vssd1 vssd1 vccd1 vccd1 _15163_/A sky130_fd_sc_hd__mux2_1
X_12374_ _19692_/Q _20180_/Q _12375_/S vssd1 vssd1 vccd1 vccd1 _12374_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14113_ _18152_/B _14119_/A _14121_/A _17952_/B vssd1 vssd1 vccd1 vccd1 _14113_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_181_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11325_ _19535_/Q _09596_/A _11225_/B _19599_/Q _09686_/Y vssd1 vssd1 vccd1 vccd1
+ _11325_/X sky130_fd_sc_hd__a221o_1
XFILLER_176_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15093_ _15019_/A _15079_/X _15092_/X vssd1 vssd1 vccd1 vccd1 _16732_/B sky130_fd_sc_hd__a21oi_4
X_19970_ _19970_/CLK _19970_/D vssd1 vssd1 vccd1 vccd1 _19970_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14044_ _14105_/A _14069_/B vssd1 vssd1 vccd1 vccd1 _14044_/Y sky130_fd_sc_hd__nor2_1
X_11256_ _11254_/X _11255_/X _11256_/S vssd1 vssd1 vccd1 vccd1 _11256_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18921_ _19140_/Q _18976_/A2 _18767_/B vssd1 vssd1 vccd1 vccd1 _18921_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10207_ _19542_/Q _09596_/B _10199_/X _10206_/Y vssd1 vssd1 vccd1 vccd1 _10207_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_122_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11187_ _11185_/X _11186_/Y _11313_/B vssd1 vssd1 vccd1 vccd1 _11187_/X sky130_fd_sc_hd__a21o_1
X_18852_ _19130_/Q _12533_/B _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18852_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_268_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10138_ _19475_/Q _09695_/Y _10137_/X _12377_/S vssd1 vssd1 vccd1 vccd1 _10138_/X
+ sky130_fd_sc_hd__a211o_1
X_17803_ _20580_/Q _17943_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20580_/D sky130_fd_sc_hd__mux2_1
XFILLER_283_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18783_ _18783_/A _18783_/B vssd1 vssd1 vccd1 vccd1 _20982_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ _20943_/Q _15995_/A2 _15994_/X vssd1 vssd1 vccd1 vccd1 _15995_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17734_ _20515_/Q _17908_/A1 _17738_/S vssd1 vssd1 vccd1 vccd1 _20515_/D sky130_fd_sc_hd__mux2_1
XFILLER_282_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14946_ _14948_/A _14980_/C vssd1 vssd1 vccd1 vccd1 _14946_/Y sky130_fd_sc_hd__nor2_2
X_10069_ _19635_/Q _10502_/A2 _10066_/X _10067_/X _10068_/X vssd1 vssd1 vccd1 vccd1
+ _10069_/X sky130_fd_sc_hd__o221a_1
XFILLER_76_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17665_ _20451_/Q _17802_/A1 _17669_/S vssd1 vssd1 vccd1 vccd1 _20451_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14877_ _15468_/A _14877_/B vssd1 vssd1 vccd1 vccd1 _14893_/B sky130_fd_sc_hd__and2_1
XFILLER_251_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19404_ _20563_/CLK _19404_/D vssd1 vssd1 vccd1 vccd1 _19404_/Q sky130_fd_sc_hd__dfxtp_1
X_16616_ _19875_/Q _17930_/A1 _16620_/S vssd1 vssd1 vccd1 vccd1 _19875_/D sky130_fd_sc_hd__mux2_1
X_13828_ _19998_/Q split1/A _13782_/X split2/A vssd1 vssd1 vccd1 vccd1 _13828_/X sky130_fd_sc_hd__a22o_4
XFILLER_223_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17596_ _20354_/Q _17835_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20354_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19335_ _20638_/CLK _19335_/D vssd1 vssd1 vccd1 vccd1 _19335_/Q sky130_fd_sc_hd__dfxtp_1
X_16547_ _16551_/A _16547_/B vssd1 vssd1 vccd1 vccd1 _19839_/D sky130_fd_sc_hd__or2_1
XFILLER_232_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ _13759_/A _13759_/B vssd1 vssd1 vccd1 vccd1 _13760_/B sky130_fd_sc_hd__nor2_8
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19266_ _20812_/CLK _19266_/D vssd1 vssd1 vccd1 vccd1 _19266_/Q sky130_fd_sc_hd__dfxtp_1
X_16478_ _19787_/Q _17801_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19787_/D sky130_fd_sc_hd__mux2_1
X_18217_ _18414_/A _18217_/B vssd1 vssd1 vccd1 vccd1 _20797_/D sky130_fd_sc_hd__and2_1
X_15429_ _15520_/B2 _15428_/X _15412_/X _15405_/Y vssd1 vssd1 vccd1 vccd1 _15429_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_19197_ _19704_/CLK _19197_/D vssd1 vssd1 vccd1 vccd1 _19197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18148_ _16711_/A _19108_/Q _18148_/S vssd1 vssd1 vccd1 vccd1 _18318_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18079_ _20767_/Q _18079_/B vssd1 vssd1 vccd1 vccd1 _18085_/C sky130_fd_sc_hd__and2_2
XFILLER_172_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20110_ _20481_/CLK _20110_/D vssd1 vssd1 vccd1 vccd1 _20110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09921_ _12015_/A1 _09920_/X _09919_/X vssd1 vssd1 vccd1 vccd1 _09921_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_252_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout705 _16566_/A2 vssd1 vssd1 vccd1 vccd1 _16578_/A2 sky130_fd_sc_hd__buf_6
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout716 _16566_/B1 vssd1 vssd1 vccd1 vccd1 _16578_/B1 sky130_fd_sc_hd__buf_6
X_20041_ _20480_/CLK _20041_/D vssd1 vssd1 vccd1 vccd1 _20041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout727 _13142_/X vssd1 vssd1 vccd1 vccd1 _13481_/A sky130_fd_sc_hd__buf_4
X_09852_ _20483_/Q _10397_/S _12100_/B1 vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__o21a_1
XFILLER_213_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout738 _14397_/A vssd1 vssd1 vccd1 vccd1 _14437_/A sky130_fd_sc_hd__buf_4
Xfanout749 _18472_/X vssd1 vssd1 vccd1 vccd1 _18985_/B sky130_fd_sc_hd__buf_6
XFILLER_258_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_252_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09783_/A _11799_/B vssd1 vssd1 vccd1 vccd1 _09784_/B sky130_fd_sc_hd__and2_4
XFILLER_274_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_109 _13474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20943_ _21009_/CLK _20943_/D vssd1 vssd1 vccd1 vccd1 _20943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _20969_/CLK _20874_/D vssd1 vssd1 vccd1 vccd1 _20874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11110_ _12332_/A _20659_/Q _12254_/C vssd1 vssd1 vccd1 vccd1 _11110_/X sky130_fd_sc_hd__or3_1
X_20308_ _20468_/CLK _20308_/D vssd1 vssd1 vccd1 vccd1 _20308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_3__f_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20408_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ _19688_/Q _20176_/Q _12097_/S vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11041_ _12429_/A1 _11039_/X _11040_/X vssd1 vssd1 vccd1 vccd1 _11041_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20239_ _21010_/CLK _20239_/D vssd1 vssd1 vccd1 vccd1 _20239_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_276_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_264_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _19147_/Q _14802_/A2 _14799_/X _17536_/D vssd1 vssd1 vccd1 vccd1 _19524_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _15882_/A1 _15769_/X _15770_/X _15779_/X vssd1 vssd1 vccd1 vccd1 _15780_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_218_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12992_ _19234_/Q _13296_/B vssd1 vssd1 vccd1 vccd1 _13365_/B sky130_fd_sc_hd__and2_2
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _19488_/Q _17806_/A1 _14733_/S vssd1 vssd1 vccd1 vccd1 _19488_/D sky130_fd_sc_hd__mux2_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11943_ _19687_/Q _20175_/Q _11944_/S vssd1 vssd1 vccd1 vccd1 _11943_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_610 input228/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_621 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_632 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _17457_/B _17443_/D _17446_/A _17452_/A vssd1 vssd1 vccd1 vccd1 _17454_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_643 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14662_ _19424_/Q _17806_/A1 _14662_/S vssd1 vssd1 vccd1 vccd1 _19424_/D sky130_fd_sc_hd__mux2_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _12194_/A1 _17910_/A1 _11873_/X _12194_/B2 vssd1 vssd1 vccd1 vccd1 _15849_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_73_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_654 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _19745_/Q _16402_/C _19746_/Q vssd1 vssd1 vccd1 vccd1 _16403_/B sky130_fd_sc_hd__a21oi_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13613_ _19661_/D _13610_/X _13612_/X _13663_/B vssd1 vssd1 vccd1 vccd1 _13613_/X
+ sky130_fd_sc_hd__a22o_4
X_10825_ _19667_/Q _20155_/Q _11358_/S vssd1 vssd1 vccd1 vccd1 _10825_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17381_ _20239_/Q _17381_/A2 _17380_/X _18740_/A vssd1 vssd1 vccd1 vccd1 _20239_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14593_ _19359_/Q _17945_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19359_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19120_ _19696_/CLK _19120_/D vssd1 vssd1 vccd1 vccd1 _19120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16332_ _19720_/Q _16332_/B vssd1 vssd1 vccd1 vccd1 _16338_/C sky130_fd_sc_hd__and2_2
X_13544_ _13544_/A _13544_/B vssd1 vssd1 vccd1 vccd1 _13544_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10756_ _10754_/X _10755_/X _12395_/S vssd1 vssd1 vccd1 vccd1 _10756_/X sky130_fd_sc_hd__mux2_1
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051_ _19051_/A _19051_/B vssd1 vssd1 vccd1 vccd1 _21044_/D sky130_fd_sc_hd__or2_1
XFILLER_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16263_ _19679_/Q _17869_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19679_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ _13469_/Y _13472_/A _13474_/X vssd1 vssd1 vccd1 vccd1 _13475_/X sky130_fd_sc_hd__a21bo_1
X_10687_ _10692_/A _19309_/Q _12406_/C vssd1 vssd1 vccd1 vccd1 _10687_/X sky130_fd_sc_hd__or3_1
X_18002_ _20738_/Q _18003_/C _20739_/Q vssd1 vssd1 vccd1 vccd1 _18004_/B sky130_fd_sc_hd__a21oi_1
XFILLER_200_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15214_ _15611_/S _15214_/B vssd1 vssd1 vccd1 vccd1 _15214_/X sky130_fd_sc_hd__or2_1
X_12426_ _12424_/X _12425_/X _12426_/S vssd1 vssd1 vccd1 vccd1 _12426_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16194_ _19621_/Q _16021_/X _16194_/S vssd1 vssd1 vccd1 vccd1 _16195_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15145_ _19736_/Q _15453_/A2 _15131_/X _15396_/A1 _15144_/X vssd1 vssd1 vccd1 vccd1
+ _15145_/X sky130_fd_sc_hd__a221o_1
XFILLER_142_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput308 _13615_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[12] sky130_fd_sc_hd__buf_4
XFILLER_126_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12357_ _12357_/A1 _12356_/X _11118_/A vssd1 vssd1 vccd1 vccd1 _12357_/Y sky130_fd_sc_hd__a21oi_1
Xoutput319 _13625_/Y vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[22] sky130_fd_sc_hd__buf_4
XFILLER_236_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11308_ _11305_/X _11306_/X _11307_/X _09507_/A _12514_/C vssd1 vssd1 vccd1 vccd1
+ _11308_/X sky130_fd_sc_hd__a221o_1
XFILLER_126_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15076_ _15076_/A _15494_/B vssd1 vssd1 vccd1 vccd1 _15076_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19953_ _20353_/CLK _19953_/D vssd1 vssd1 vccd1 vccd1 _19953_/Q sky130_fd_sc_hd__dfxtp_1
X_12288_ _12288_/A _12288_/B _12288_/C vssd1 vssd1 vccd1 vccd1 _12290_/D sky130_fd_sc_hd__and3_1
X_14027_ _19208_/Q _14097_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _14027_/X sky130_fd_sc_hd__mux2_1
X_18904_ _18526_/X _18964_/B _18902_/Y _18903_/Y vssd1 vssd1 vccd1 vccd1 _18905_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_206_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11239_ _11239_/A1 _13960_/A2 _11238_/X _11239_/B1 _19831_/Q vssd1 vssd1 vccd1 vccd1
+ _11239_/X sky130_fd_sc_hd__o32a_1
XFILLER_45_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19884_ _20081_/CLK _19884_/D vssd1 vssd1 vccd1 vccd1 _19884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18835_ _18835_/A _18835_/B vssd1 vssd1 vccd1 vccd1 _20990_/D sky130_fd_sc_hd__nor2_1
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18766_ _19118_/Q _18764_/X _18901_/S vssd1 vssd1 vccd1 vccd1 _18766_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15978_ _11367_/A _15978_/A2 _15954_/A _16063_/B2 vssd1 vssd1 vccd1 vccd1 _15979_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_283_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17717_ _20498_/Q _17751_/A1 _17742_/S vssd1 vssd1 vccd1 vccd1 _20498_/D sky130_fd_sc_hd__mux2_1
X_14929_ _14955_/B vssd1 vssd1 vccd1 vccd1 _15014_/B sky130_fd_sc_hd__inv_2
XFILLER_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_264_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18697_ _20949_/Q _18175_/Y _18719_/S vssd1 vssd1 vccd1 vccd1 _18698_/B sky130_fd_sc_hd__mux2_1
XFILLER_91_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17648_ _20434_/Q _17857_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20434_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17579_ _20337_/Q _17890_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20337_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19318_ _20673_/CLK _19318_/D vssd1 vssd1 vccd1 vccd1 _19318_/Q sky130_fd_sc_hd__dfxtp_1
X_20590_ _20659_/CLK _20590_/D vssd1 vssd1 vccd1 vccd1 _20590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19249_ _21016_/CLK _19249_/D vssd1 vssd1 vccd1 vccd1 _19249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_158_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20742_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_118_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout502 _17813_/X vssd1 vssd1 vccd1 vccd1 _17845_/S sky130_fd_sc_hd__buf_12
X_09904_ _09889_/X _09903_/X _12153_/A1 vssd1 vssd1 vccd1 vccd1 _09904_/X sky130_fd_sc_hd__a21o_2
XFILLER_104_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout513 _17711_/X vssd1 vssd1 vccd1 vccd1 _17738_/S sky130_fd_sc_hd__buf_4
XFILLER_263_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout524 _17608_/X vssd1 vssd1 vccd1 vccd1 _17637_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout535 _17540_/X vssd1 vssd1 vccd1 vccd1 _17570_/S sky130_fd_sc_hd__buf_12
XFILLER_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20024_ _20664_/CLK _20024_/D vssd1 vssd1 vccd1 vccd1 _20024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_258_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout546 _17144_/S vssd1 vssd1 vccd1 vccd1 _17132_/S sky130_fd_sc_hd__buf_12
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09835_ _19388_/Q _10603_/B _09833_/X _11718_/S _09834_/X vssd1 vssd1 vccd1 vccd1
+ _09835_/X sky130_fd_sc_hd__o221a_1
Xfanout557 _16673_/X vssd1 vssd1 vccd1 vccd1 _16701_/S sky130_fd_sc_hd__buf_4
Xfanout568 _16490_/X vssd1 vssd1 vccd1 vccd1 _16519_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_247_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout579 _16245_/X vssd1 vssd1 vccd1 vccd1 _16272_/S sky130_fd_sc_hd__buf_12
XFILLER_281_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09766_ _20484_/Q _11616_/B _12015_/A1 vssd1 vssd1 vccd1 vccd1 _09766_/X sky130_fd_sc_hd__a21o_1
XFILLER_58_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09697_ _11514_/A1 _20712_/Q _11599_/S _09696_/X vssd1 vssd1 vccd1 vccd1 _09697_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _21025_/CLK _20926_/D vssd1 vssd1 vccd1 vccd1 _20926_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ _21018_/CLK _20857_/D vssd1 vssd1 vccd1 vccd1 _20857_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _20598_/Q _10628_/S _10609_/X vssd1 vssd1 vccd1 vccd1 _10610_/X sky130_fd_sc_hd__a21o_1
XFILLER_211_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ _11581_/X _11583_/X _11589_/X _12135_/A _12137_/A1 vssd1 vssd1 vccd1 vccd1
+ _11590_/X sky130_fd_sc_hd__o221a_1
X_20788_ _20796_/CLK _20788_/D vssd1 vssd1 vccd1 vccd1 _20788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _10540_/A _10540_/B _10641_/B vssd1 vssd1 vccd1 vccd1 _13155_/A sky130_fd_sc_hd__a21o_2
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260_ _20969_/Q _13397_/B vssd1 vssd1 vccd1 vccd1 _13260_/Y sky130_fd_sc_hd__nand2_1
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10472_ _10035_/Y _10466_/X _10471_/X _10461_/X _10024_/X vssd1 vssd1 vccd1 vccd1
+ _10472_/X sky130_fd_sc_hd__a32o_2
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12211_ _20362_/Q _12295_/B vssd1 vssd1 vccd1 vccd1 _12211_/X sky130_fd_sc_hd__or2_1
XFILLER_157_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13191_ _16598_/A _16594_/B vssd1 vssd1 vccd1 vccd1 _13191_/X sky130_fd_sc_hd__and2_1
XFILLER_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12142_ _19394_/Q _20685_/Q _12148_/S vssd1 vssd1 vccd1 vccd1 _12142_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16950_ _19701_/Q _19699_/Q vssd1 vssd1 vccd1 vccd1 _16950_/Y sky130_fd_sc_hd__nand2_8
X_12073_ _12073_/A1 _12062_/X _12065_/X _12072_/X _12073_/C1 vssd1 vssd1 vccd1 vccd1
+ _12073_/X sky130_fd_sc_hd__a311o_1
XFILLER_123_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11024_ _11022_/X _11023_/X _11033_/S vssd1 vssd1 vccd1 vccd1 _11024_/X sky130_fd_sc_hd__mux2_1
X_15901_ _14837_/S _15258_/B _15262_/Y _15258_/A vssd1 vssd1 vccd1 vccd1 _15901_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16881_ _19231_/Q _17003_/B _16964_/B1 _19100_/Q _16880_/X vssd1 vssd1 vccd1 vccd1
+ _16881_/X sky130_fd_sc_hd__o221a_2
XFILLER_238_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832_ _20809_/Q _15941_/A2 _15825_/X _15941_/B2 _15831_/X vssd1 vssd1 vccd1 vccd1
+ _15832_/X sky130_fd_sc_hd__a221o_2
X_18620_ _19508_/Q _18628_/B vssd1 vssd1 vccd1 vccd1 _18620_/Y sky130_fd_sc_hd__nand2_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _20910_/Q fanout750/X _18550_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18552_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15763_ _15763_/A _15763_/B _15981_/B vssd1 vssd1 vccd1 vccd1 _15763_/Y sky130_fd_sc_hd__nand3_1
XFILLER_206_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _12975_/A _12975_/B _12975_/C _12975_/D vssd1 vssd1 vccd1 vccd1 _12975_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_45_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ _20286_/Q _17502_/B vssd1 vssd1 vccd1 vccd1 _17502_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14714_ _19471_/Q _17929_/A1 _14733_/S vssd1 vssd1 vccd1 vccd1 _19471_/D sky130_fd_sc_hd__mux2_1
X_18482_ _18598_/A _18482_/B vssd1 vssd1 vccd1 vccd1 _20887_/D sky130_fd_sc_hd__nor2_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _19823_/Q _12009_/A2 _11924_/X _11563_/S _11925_/X vssd1 vssd1 vccd1 vccd1
+ _11926_/X sky130_fd_sc_hd__o221a_1
X_15694_ _20964_/Q _15939_/A2 _15996_/B1 _20836_/Q _15693_/X vssd1 vssd1 vccd1 vccd1
+ _15694_/X sky130_fd_sc_hd__a221o_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_440 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_451 _13775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_462 _19245_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17433_ _20261_/Q _20254_/Q _17433_/S vssd1 vssd1 vccd1 vccd1 _17434_/B sky130_fd_sc_hd__mux2_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14645_ _19407_/Q _17929_/A1 _14662_/S vssd1 vssd1 vccd1 vccd1 _19407_/D sky130_fd_sc_hd__mux2_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_473 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11857_ _19686_/Q _20174_/Q _11944_/S vssd1 vssd1 vccd1 vccd1 _11857_/X sky130_fd_sc_hd__mux2_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_484 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_495 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10808_ _10553_/B _10124_/Y _10807_/X _10118_/X vssd1 vssd1 vccd1 vccd1 _10808_/Y
+ sky130_fd_sc_hd__o211ai_2
X_17364_ _20230_/Q _17364_/A2 _17370_/B1 _20279_/Q _17370_/C1 vssd1 vssd1 vccd1 vccd1
+ _17364_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14576_ _19342_/Q _17928_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19342_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11788_ _11788_/A _11788_/B _11788_/C vssd1 vssd1 vccd1 vccd1 _11788_/X sky130_fd_sc_hd__or3_4
X_16315_ _18086_/A _16315_/B _16316_/B vssd1 vssd1 vccd1 vccd1 _19713_/D sky130_fd_sc_hd__nor3_1
X_19103_ _19609_/CLK _19103_/D vssd1 vssd1 vccd1 vccd1 _19103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13527_ _13526_/A _13526_/B _13526_/C vssd1 vssd1 vccd1 vccd1 _13527_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17295_ _20204_/Q _17328_/A2 _17293_/X _17294_/X _17974_/B1 vssd1 vssd1 vccd1 vccd1
+ _20204_/D sky130_fd_sc_hd__o221a_1
X_10739_ _20531_/Q _12313_/S vssd1 vssd1 vccd1 vccd1 _10739_/X sky130_fd_sc_hd__or2_1
XFILLER_159_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19034_ _18280_/Y _19046_/A2 _19048_/B1 _12552_/A _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19034_/X sky130_fd_sc_hd__a221o_1
X_16246_ _19662_/Q _17780_/A1 _16275_/S vssd1 vssd1 vccd1 vccd1 _19662_/D sky130_fd_sc_hd__mux2_1
X_13458_ _14524_/A1 _09497_/Y _16241_/A _13457_/X vssd1 vssd1 vccd1 vccd1 _13458_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12409_ _12407_/X _12408_/X _12414_/S vssd1 vssd1 vccd1 vccd1 _12409_/X sky130_fd_sc_hd__mux2_1
X_16177_ _16191_/A _16177_/B vssd1 vssd1 vccd1 vccd1 _19612_/D sky130_fd_sc_hd__and2_1
X_13389_ _13389_/A _13389_/B _13389_/C vssd1 vssd1 vccd1 vccd1 _13389_/X sky130_fd_sc_hd__or3_2
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15128_ _11786_/C _15127_/B _15127_/Y _16030_/D1 vssd1 vssd1 vccd1 vccd1 _15128_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19936_ _20467_/CLK _19936_/D vssd1 vssd1 vccd1 vccd1 _19936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_269_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15059_ _14811_/X _14815_/X _15062_/S vssd1 vssd1 vccd1 vccd1 _15059_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19867_ _20720_/CLK _19867_/D vssd1 vssd1 vccd1 vccd1 _19867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09620_ _16454_/B _10152_/S _09619_/X _09616_/Y vssd1 vssd1 vccd1 vccd1 _09630_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_110_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18818_ _18596_/Y _18818_/A2 _18816_/Y _18817_/Y vssd1 vssd1 vccd1 vccd1 _18818_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_255_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19798_ _20379_/CLK _19798_/D vssd1 vssd1 vccd1 vccd1 _19798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09551_ _14895_/A _12510_/C vssd1 vssd1 vccd1 vccd1 _09552_/B sky130_fd_sc_hd__or2_2
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18749_ _20975_/Q _18305_/Y _18749_/S vssd1 vssd1 vccd1 vccd1 _18750_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09482_ _20794_/Q vssd1 vssd1 vccd1 vccd1 _09482_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20711_ _20711_/CLK _20711_/D vssd1 vssd1 vccd1 vccd1 _20711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20642_ _20685_/CLK _20642_/D vssd1 vssd1 vccd1 vccd1 _20642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20573_ _20573_/CLK _20573_/D vssd1 vssd1 vccd1 vccd1 _20573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1308 _14836_/S vssd1 vssd1 vccd1 vccd1 _14815_/S sky130_fd_sc_hd__buf_4
Xfanout1319 _12467_/Y vssd1 vssd1 vccd1 vccd1 _14878_/B sky130_fd_sc_hd__buf_6
XFILLER_87_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20007_ _20751_/CLK _20007_/D vssd1 vssd1 vccd1 vccd1 _20007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09818_ _09806_/S _09817_/X _09816_/X _12068_/C1 vssd1 vssd1 vccd1 vccd1 _09818_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_275_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_55_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20463_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_235_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09749_ _09748_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09749_/X sky130_fd_sc_hd__and2b_1
XFILLER_262_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_261_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12751_/X _12752_/Y _12757_/Y _12758_/X vssd1 vssd1 vccd1 vccd1 _12771_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _19883_/Q _11718_/S _11708_/B _11709_/X _11710_/X vssd1 vssd1 vccd1 vccd1
+ _11711_/X sky130_fd_sc_hd__a311o_1
XFILLER_203_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ _21011_/CLK _20909_/D vssd1 vssd1 vccd1 vccd1 _20909_/Q sky130_fd_sc_hd__dfxtp_1
X_12691_ _12693_/A _12692_/D vssd1 vssd1 vccd1 vccd1 _13526_/C sky130_fd_sc_hd__nor2_1
XFILLER_242_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _19245_/Q _14438_/A2 _14429_/X _14802_/C1 vssd1 vssd1 vccd1 vccd1 _19245_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _19642_/Q _19948_/Q _19286_/Q _20073_/Q _11642_/S0 _12003_/C vssd1 vssd1
+ vccd1 vccd1 _11642_/X sky130_fd_sc_hd__mux4_1
XFILLER_42_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14361_ _14361_/A _14361_/B vssd1 vssd1 vccd1 vccd1 _14366_/A sky130_fd_sc_hd__nor2_1
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ _11575_/A vssd1 vssd1 vccd1 vccd1 _13162_/A sky130_fd_sc_hd__inv_2
XFILLER_211_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16100_ _19574_/Q _16079_/B _16099_/X _16107_/B1 vssd1 vssd1 vccd1 vccd1 _19574_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput18 core_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_4
XFILLER_167_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13312_ _19227_/Q _13450_/A _14110_/B vssd1 vssd1 vccd1 vccd1 _13312_/Y sky130_fd_sc_hd__a21oi_1
X_17080_ _20052_/Q _17114_/A1 _17080_/S vssd1 vssd1 vccd1 vccd1 _20052_/D sky130_fd_sc_hd__mux2_1
X_10524_ _10516_/S _10519_/X _10523_/X vssd1 vssd1 vccd1 vccd1 _10524_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput29 core_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14292_ _14283_/A _14280_/Y _14282_/B vssd1 vssd1 vccd1 vccd1 _14302_/B sky130_fd_sc_hd__o21ai_2
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16031_ _16029_/X _16030_/X _15890_/B vssd1 vssd1 vccd1 vccd1 _16031_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13243_ _14780_/C1 _13220_/Y _13242_/X _13141_/X vssd1 vssd1 vccd1 vccd1 _13245_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_108_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10455_ _10640_/B _10455_/B vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__xor2_4
XFILLER_164_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13174_ _12109_/Y _13432_/B _12111_/B vssd1 vssd1 vccd1 vccd1 _13431_/B sky130_fd_sc_hd__o21a_4
X_10386_ _19538_/Q _09596_/B _10369_/X _10385_/Y vssd1 vssd1 vccd1 vccd1 _10386_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_163_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12125_ _12125_/A1 _12124_/X _12123_/X vssd1 vssd1 vccd1 vccd1 _12125_/X sky130_fd_sc_hd__o21a_1
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17982_ _20732_/Q _20731_/Q _17982_/C vssd1 vssd1 vccd1 vccd1 _17984_/A sky130_fd_sc_hd__and3_1
XFILLER_111_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1820 _19177_/Q vssd1 vssd1 vccd1 vccd1 _12519_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19721_ _21026_/CLK _19721_/D vssd1 vssd1 vccd1 vccd1 _19721_/Q sky130_fd_sc_hd__dfxtp_2
X_16933_ input57/X input92/X _16975_/S vssd1 vssd1 vccd1 vccd1 _16933_/X sky130_fd_sc_hd__mux2_8
X_12056_ _12048_/X _12049_/X _12056_/S vssd1 vssd1 vccd1 vccd1 _12056_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1831 _19173_/Q vssd1 vssd1 vccd1 vccd1 _12513_/D sky130_fd_sc_hd__buf_12
XFILLER_238_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1842 _12125_/A1 vssd1 vssd1 vccd1 vccd1 _10057_/S sky130_fd_sc_hd__buf_6
XFILLER_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1853 _09776_/S vssd1 vssd1 vccd1 vccd1 _11949_/S sky130_fd_sc_hd__buf_6
Xfanout1864 _11384_/S vssd1 vssd1 vccd1 vccd1 _12431_/A1 sky130_fd_sc_hd__buf_6
XFILLER_238_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11007_ _11008_/A1 _19900_/Q _10986_/B _20025_/Q vssd1 vssd1 vccd1 vccd1 _11007_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19652_ _20662_/CLK _19652_/D vssd1 vssd1 vccd1 vccd1 _19652_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1875 _12357_/A1 vssd1 vssd1 vccd1 vccd1 _12420_/B1 sky130_fd_sc_hd__buf_6
XFILLER_238_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16864_ _16884_/S input83/X vssd1 vssd1 vccd1 vccd1 _16864_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1886 _14802_/C1 vssd1 vssd1 vccd1 vccd1 _17434_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_237_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1897 _18736_/A vssd1 vssd1 vccd1 vccd1 _18748_/A sky130_fd_sc_hd__clkbuf_4
X_18603_ _20924_/Q _18619_/B vssd1 vssd1 vccd1 vccd1 _18603_/Y sky130_fd_sc_hd__nand2_1
X_15815_ _19549_/Q _15980_/A2 _15814_/Y _16191_/A vssd1 vssd1 vccd1 vccd1 _19549_/D
+ sky130_fd_sc_hd__o211a_1
X_19583_ _19590_/CLK _19583_/D vssd1 vssd1 vccd1 vccd1 _19583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16795_ _20404_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16795_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15746_ _21032_/Q _21000_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _15746_/X sky130_fd_sc_hd__mux2_1
X_18534_ _18932_/A _18534_/B vssd1 vssd1 vccd1 vccd1 _20904_/D sky130_fd_sc_hd__nor2_1
XFILLER_280_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12958_ _19251_/Q _12964_/A2 _16716_/A _19999_/Q vssd1 vssd1 vccd1 vccd1 _12959_/B
+ sky130_fd_sc_hd__a22o_2
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11909_ _20422_/Q _11915_/S _11895_/X _11917_/S vssd1 vssd1 vccd1 vccd1 _11909_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_261_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18465_ _18462_/X _18464_/X _18783_/A vssd1 vssd1 vccd1 vccd1 _20883_/D sky130_fd_sc_hd__a21oi_1
X_15677_ _13427_/B _15676_/X _16034_/S vssd1 vssd1 vccd1 vccd1 _15677_/X sky130_fd_sc_hd__mux2_1
XANTENNA_270 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12889_ _12889_/A _12889_/B vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__or2_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_281 _20623_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17416_ _20261_/Q _20253_/Q _17442_/A vssd1 vssd1 vccd1 vccd1 _17416_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_292 input222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14628_ _19392_/Q _17878_/A1 _14628_/S vssd1 vssd1 vccd1 vccd1 _19392_/D sky130_fd_sc_hd__mux2_1
X_18396_ _18396_/A _18396_/B vssd1 vssd1 vccd1 vccd1 _20852_/D sky130_fd_sc_hd__and2_1
XFILLER_159_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17347_ _20222_/Q _17363_/A2 _17346_/X _18694_/A vssd1 vssd1 vccd1 vccd1 _20222_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14559_ _19329_/Q _17111_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19329_/D sky130_fd_sc_hd__mux2_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ input272/X _17290_/B vssd1 vssd1 vccd1 vccd1 _17278_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16229_ _19652_/Q _17915_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19652_/D sky130_fd_sc_hd__mux2_1
X_19017_ _12555_/A _12555_/B _18760_/X vssd1 vssd1 vccd1 vccd1 _19017_/X sky130_fd_sc_hd__o21a_4
XFILLER_228_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19919_ _20479_/CLK _19919_/D vssd1 vssd1 vccd1 vccd1 _19919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_269_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_260_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_249_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09603_ _14668_/B _17538_/C _17709_/C vssd1 vssd1 vccd1 vccd1 _17884_/A sky130_fd_sc_hd__nand3_4
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ _19154_/Q _09734_/B vssd1 vssd1 vccd1 vccd1 _13869_/A sky130_fd_sc_hd__nor2_2
XFILLER_243_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_173_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21010_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_196_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20625_ _20657_/CLK _20625_/D vssd1 vssd1 vccd1 vccd1 _20625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_102_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20794_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_177_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20556_ _20688_/CLK _20556_/D vssd1 vssd1 vccd1 vccd1 _20556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20487_ _20583_/CLK _20487_/D vssd1 vssd1 vccd1 vccd1 _20487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10240_ _09689_/A _10232_/X _10239_/X _10223_/X vssd1 vssd1 vccd1 vccd1 _10240_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ _10169_/X _10170_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _10171_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput480 _19502_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[8] sky130_fd_sc_hd__buf_4
XFILLER_267_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1105 _17111_/A1 vssd1 vssd1 vccd1 vccd1 _17704_/A1 sky130_fd_sc_hd__clkbuf_2
Xfanout1116 _17870_/A1 vssd1 vssd1 vccd1 vccd1 _17695_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1127 _11534_/X vssd1 vssd1 vccd1 vccd1 _17936_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout1138 _09947_/X vssd1 vssd1 vccd1 vccd1 _17872_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout1149 _17943_/A1 vssd1 vssd1 vccd1 vccd1 _17666_/A1 sky130_fd_sc_hd__clkbuf_4
X_13930_ _19134_/Q _13932_/B1 _13906_/X _13345_/X vssd1 vssd1 vccd1 vccd1 _19134_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21039_ _21043_/CLK _21039_/D vssd1 vssd1 vccd1 vccd1 _21039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ _16066_/B _13860_/B _13860_/C _14244_/A1 vssd1 vssd1 vccd1 vccd1 _14073_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15600_ _20961_/Q _15939_/A2 _15996_/B1 _20833_/Q _15599_/X vssd1 vssd1 vccd1 vccd1
+ _15600_/X sky130_fd_sc_hd__a221o_4
XFILLER_216_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12812_ _12483_/Y _12811_/X _15741_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12812_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16580_ _19856_/Q _16592_/A2 _16592_/B1 input27/X vssd1 vssd1 vccd1 vccd1 _16581_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13792_ _13798_/A1 _13826_/A1 _13708_/B _13826_/B1 input226/X vssd1 vssd1 vccd1 vccd1
+ _13792_/X sky130_fd_sc_hd__a32o_2
XFILLER_222_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15531_ _20735_/Q _16041_/A2 _16041_/B1 _20767_/Q vssd1 vssd1 vccd1 vccd1 _15531_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12739_/Y _12742_/X _12716_/B vssd1 vssd1 vccd1 vccd1 _12747_/A sky130_fd_sc_hd__a21o_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _18520_/B vssd1 vssd1 vccd1 vccd1 _18250_/Y sky130_fd_sc_hd__clkinv_2
X_15462_ _19537_/Q _15402_/A _15461_/Y _16159_/C1 vssd1 vssd1 vccd1 vccd1 _19537_/D
+ sky130_fd_sc_hd__o211a_1
X_12674_ _12674_/A _12674_/B _12674_/C vssd1 vssd1 vccd1 vccd1 _12675_/C sky130_fd_sc_hd__nand3_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _20165_/Q _17692_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20165_/D sky130_fd_sc_hd__mux2_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14413_ _19523_/Q _14413_/B vssd1 vssd1 vccd1 vccd1 _14424_/A sky130_fd_sc_hd__and2_1
XFILLER_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18181_ _20790_/Q _18180_/Y _18311_/S vssd1 vssd1 vccd1 vccd1 _18182_/B sky130_fd_sc_hd__mux2_1
X_11625_ _12003_/A _19385_/Q _20676_/Q _11642_/S0 vssd1 vssd1 vccd1 vccd1 _11625_/X
+ sky130_fd_sc_hd__a22o_1
X_15393_ _17263_/A _15392_/X _15452_/S vssd1 vssd1 vccd1 vccd1 _15393_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17132_ _20100_/Q _17657_/A1 _17132_/S vssd1 vssd1 vccd1 vccd1 _20100_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14344_ _14343_/A _14343_/B _14343_/C vssd1 vssd1 vccd1 vccd1 _14354_/B sky130_fd_sc_hd__a21o_1
X_11556_ _19881_/Q _11563_/S _11616_/B _11554_/X _11555_/X vssd1 vssd1 vccd1 vccd1
+ _11556_/X sky130_fd_sc_hd__a311o_1
X_17063_ _20035_/Q _17097_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20035_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ _12517_/B _11367_/B _11398_/S vssd1 vssd1 vccd1 vccd1 _10540_/B sky130_fd_sc_hd__o21a_2
X_14275_ _14275_/A1 _14274_/X _13409_/X vssd1 vssd1 vccd1 vccd1 _14276_/C sky130_fd_sc_hd__o21a_1
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ _19679_/Q _20167_/Q _12174_/S vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16014_ _20912_/Q _16043_/A2 _16043_/B1 _16013_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _16014_/X sky130_fd_sc_hd__a221o_1
X_13226_ _13086_/A _13086_/B _13086_/C vssd1 vssd1 vccd1 vccd1 _13226_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_143_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _19377_/Q _10502_/A2 _10436_/X _12072_/A1 _10437_/X vssd1 vssd1 vccd1 vccd1
+ _10438_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13157_ _10113_/A _13425_/B _15500_/S vssd1 vssd1 vccd1 vccd1 _13424_/B sky130_fd_sc_hd__a21bo_4
X_10369_ _19538_/Q _09596_/A _09613_/B _19602_/Q _11246_/A1 vssd1 vssd1 vccd1 vccd1
+ _10369_/X sky130_fd_sc_hd__a221o_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12108_ _19520_/Q _15904_/A _15895_/S vssd1 vssd1 vccd1 vccd1 _12114_/B sky130_fd_sc_hd__mux2_8
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _20726_/Q _17965_/B vssd1 vssd1 vccd1 vccd1 _17971_/C sky130_fd_sc_hd__and2_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _20973_/Q _20907_/Q _13216_/A vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__a21oi_2
XFILLER_285_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19704_ _19704_/CLK _19704_/D vssd1 vssd1 vccd1 vccd1 _19704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12039_ _12039_/A1 _10470_/B split7/X vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__a21o_4
X_16916_ _16932_/A1 _16915_/X _16932_/B1 vssd1 vssd1 vccd1 vccd1 _16916_/Y sky130_fd_sc_hd__o21ai_2
Xfanout1650 _12531_/Y vssd1 vssd1 vccd1 vccd1 _18830_/A sky130_fd_sc_hd__clkbuf_4
Xfanout1661 _09646_/Y vssd1 vssd1 vccd1 vccd1 _14041_/A2 sky130_fd_sc_hd__buf_4
XFILLER_239_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1672 _13853_/B vssd1 vssd1 vccd1 vccd1 _14002_/A1 sky130_fd_sc_hd__clkbuf_8
X_17896_ _20667_/Q _17896_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20667_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1683 _11191_/A vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_66_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1694 _11191_/A vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__clkbuf_16
X_19635_ _20472_/CLK _19635_/D vssd1 vssd1 vccd1 vccd1 _19635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16847_ _16846_/A _09525_/Y _16809_/X _16846_/Y vssd1 vssd1 vccd1 vccd1 _16847_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_92_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19566_ _19590_/CLK _19566_/D vssd1 vssd1 vccd1 vccd1 _19566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_280_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16778_ _17008_/A1 _16777_/X _17008_/B1 vssd1 vssd1 vccd1 vccd1 _16778_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_34_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18517_ _18628_/B _18517_/B vssd1 vssd1 vccd1 vccd1 _18517_/X sky130_fd_sc_hd__or2_1
X_15729_ _15890_/B _15712_/Y _15728_/X _15976_/B2 vssd1 vssd1 vccd1 vccd1 _15729_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_206_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19497_ _19696_/CLK _19497_/D vssd1 vssd1 vccd1 vccd1 _19497_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20713_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18448_ _18736_/A _18448_/B vssd1 vssd1 vccd1 vccd1 _20878_/D sky130_fd_sc_hd__and2_1
XFILLER_61_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_279_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18379_ _18547_/B _18387_/B vssd1 vssd1 vccd1 vccd1 _18379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_239_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20410_ _20410_/CLK _20410_/D vssd1 vssd1 vccd1 vccd1 _20410_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_175_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20341_ _20341_/CLK _20341_/D vssd1 vssd1 vccd1 vccd1 _20341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20272_ _20273_/CLK _20272_/D vssd1 vssd1 vccd1 vccd1 _20272_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_249_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput208 localMemory_wb_adr_i[4] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__clkbuf_2
Xinput219 localMemory_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_hd__buf_12
XFILLER_102_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09517_ _19659_/Q vssd1 vssd1 vccd1 vccd1 _13853_/B sky130_fd_sc_hd__inv_6
XFILLER_253_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11410_ _11409_/A _10645_/A _11772_/A _11409_/X vssd1 vssd1 vccd1 vccd1 _11791_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_184_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20608_ _20676_/CLK _20608_/D vssd1 vssd1 vccd1 vccd1 _20608_/Q sky130_fd_sc_hd__dfxtp_1
X_12390_ _19396_/Q _20687_/Q _12397_/S vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11341_ _19670_/Q _20158_/Q _11342_/S vssd1 vssd1 vccd1 vccd1 _11341_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20539_ _20539_/CLK _20539_/D vssd1 vssd1 vccd1 vccd1 _20539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ _19189_/Q _14108_/A2 _14059_/X _16107_/B1 vssd1 vssd1 vccd1 vccd1 _19189_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11272_ _11273_/A1 _19897_/Q _10324_/S _20022_/Q vssd1 vssd1 vccd1 vccd1 _11272_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_153_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ _20973_/Q _20907_/Q vssd1 vssd1 vccd1 vccd1 _13011_/Y sky130_fd_sc_hd__nand2_1
X_10223_ _11101_/A _10221_/X _10222_/X _12311_/C1 vssd1 vssd1 vccd1 vccd1 _10223_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_180_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20665_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_239_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10154_ _19636_/Q _19942_/Q _11358_/S vssd1 vssd1 vccd1 vccd1 _10154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_267_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14962_ _14957_/B _15021_/B _15308_/C vssd1 vssd1 vccd1 vccd1 _14972_/A sky130_fd_sc_hd__o21a_1
X_17750_ _20529_/Q _17750_/A1 _17777_/S vssd1 vssd1 vccd1 vccd1 _20529_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10085_ _20313_/Q _10518_/S _10084_/X vssd1 vssd1 vccd1 vccd1 _10085_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16701_ _19956_/Q _17111_/A1 _16701_/S vssd1 vssd1 vccd1 vccd1 _19956_/D sky130_fd_sc_hd__mux2_1
X_13913_ _13913_/A _13919_/S vssd1 vssd1 vccd1 vccd1 _13913_/Y sky130_fd_sc_hd__nand2_1
X_17681_ _20465_/Q _17750_/A1 _17706_/S vssd1 vssd1 vccd1 vccd1 _20465_/D sky130_fd_sc_hd__mux2_1
X_14893_ _14893_/A _14893_/B _14891_/X vssd1 vssd1 vccd1 vccd1 _14893_/X sky130_fd_sc_hd__or3b_4
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19420_ _20579_/CLK _19420_/D vssd1 vssd1 vccd1 vccd1 _19420_/Q sky130_fd_sc_hd__dfxtp_1
X_13844_ _17226_/B _13844_/B _20216_/Q vssd1 vssd1 vccd1 vccd1 _13844_/X sky130_fd_sc_hd__or3b_1
XFILLER_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16632_ _19891_/Q _17806_/A1 _16632_/S vssd1 vssd1 vccd1 vccd1 _19891_/D sky130_fd_sc_hd__mux2_1
XFILLER_262_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19351_ _20574_/CLK _19351_/D vssd1 vssd1 vccd1 vccd1 _19351_/Q sky130_fd_sc_hd__dfxtp_1
X_16563_ _16591_/A _16563_/B vssd1 vssd1 vccd1 vccd1 _19847_/D sky130_fd_sc_hd__or2_1
XFILLER_222_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13775_ _13775_/A _13775_/B vssd1 vssd1 vccd1 vccd1 _13775_/X sky130_fd_sc_hd__and2_1
X_10987_ _20560_/Q _11169_/B _10986_/X _12304_/C1 vssd1 vssd1 vccd1 vccd1 _10987_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18302_ _18720_/A _18302_/B vssd1 vssd1 vccd1 vccd1 _20814_/D sky130_fd_sc_hd__and2_1
X_15514_ _20798_/Q _16047_/A2 _15512_/X _15513_/X vssd1 vssd1 vccd1 vccd1 _15514_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_231_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _12726_/A _12726_/B _12726_/C _12726_/D vssd1 vssd1 vccd1 vccd1 _12791_/A
+ sky130_fd_sc_hd__or4_4
X_16494_ _19801_/Q _17855_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19801_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19282_ _20692_/CLK _19282_/D vssd1 vssd1 vccd1 vccd1 _19282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15445_ _20732_/Q _15445_/A2 _15445_/B1 _20764_/Q vssd1 vssd1 vccd1 vccd1 _15445_/X
+ sky130_fd_sc_hd__a22o_1
X_18233_ _19542_/Q _18248_/B vssd1 vssd1 vccd1 vccd1 _18233_/Y sky130_fd_sc_hd__nand2b_4
X_12657_ _14803_/A1 _12657_/A2 _12682_/B _12656_/X vssd1 vssd1 vccd1 vccd1 _12657_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11608_ _12144_/C1 _11597_/X _11600_/X _11607_/X _12152_/A1 vssd1 vssd1 vccd1 vccd1
+ _11608_/X sky130_fd_sc_hd__a311o_1
XFILLER_128_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18164_ _18163_/A _14130_/B _18163_/Y vssd1 vssd1 vccd1 vccd1 _18463_/B sky130_fd_sc_hd__o21ai_2
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15376_ _15610_/A1 _15354_/A _15610_/B1 vssd1 vssd1 vccd1 vccd1 _15376_/Y sky130_fd_sc_hd__o21ai_2
X_12588_ _12588_/A _12588_/B _12588_/C _12588_/D vssd1 vssd1 vccd1 vccd1 _18765_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_8_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17115_ _20085_/Q _17917_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20085_/D sky130_fd_sc_hd__mux2_1
X_14327_ _13373_/A _14326_/X _13373_/Y vssd1 vssd1 vccd1 vccd1 _14328_/C sky130_fd_sc_hd__o21a_1
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11539_ _19678_/Q _09928_/S _11538_/X _09986_/C vssd1 vssd1 vccd1 vccd1 _11539_/X
+ sky130_fd_sc_hd__o211a_1
X_18095_ _20773_/Q _18095_/B vssd1 vssd1 vccd1 vccd1 _18101_/C sky130_fd_sc_hd__and2_2
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17046_ _20021_/Q _20020_/Q _18821_/A _17045_/X vssd1 vssd1 vccd1 vccd1 _17046_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14258_ _19508_/Q _14259_/B vssd1 vssd1 vccd1 vccd1 _14271_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ _13209_/A _13209_/B _13209_/C vssd1 vssd1 vccd1 vccd1 _13209_/Y sky130_fd_sc_hd__nand3_1
X_14189_ _14189_/A _14189_/B vssd1 vssd1 vccd1 vccd1 _14191_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout909 _15601_/S vssd1 vssd1 vccd1 vccd1 _15569_/S sky130_fd_sc_hd__buf_6
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _21018_/Q _18997_/B vssd1 vssd1 vccd1 vccd1 _18997_/X sky130_fd_sc_hd__or2_1
XFILLER_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _20717_/Q _17948_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20717_/D sky130_fd_sc_hd__mux2_1
XFILLER_273_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1480 _12426_/S vssd1 vssd1 vccd1 vccd1 _11945_/S sky130_fd_sc_hd__clkbuf_16
Xfanout1491 _12342_/A vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_238_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17879_ _20652_/Q _17913_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20652_/D sky130_fd_sc_hd__mux2_1
XFILLER_253_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19618_ _19618_/CLK _19618_/D vssd1 vssd1 vccd1 vccd1 _19618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20890_ _21019_/CLK _20890_/D vssd1 vssd1 vccd1 vccd1 _20890_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19549_ _20425_/CLK _19549_/D vssd1 vssd1 vccd1 vccd1 _19549_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20324_ _20580_/CLK _20324_/D vssd1 vssd1 vccd1 vccd1 _20324_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_2__f_wb_clk_i clkbuf_3_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_266_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20255_ _20261_/CLK _20255_/D vssd1 vssd1 vccd1 vccd1 _20255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_282_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20186_ _20428_/CLK _20186_/D vssd1 vssd1 vccd1 vccd1 _20186_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ _09752_/A _19482_/Q _19450_/Q _11936_/S _11946_/C1 vssd1 vssd1 vccd1 vccd1
+ _09997_/X sky130_fd_sc_hd__a221o_1
XFILLER_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10910_ _09689_/C _10898_/X _10901_/X _10909_/X vssd1 vssd1 vccd1 vccd1 _10928_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _11983_/A1 _19487_/Q _19455_/Q _11889_/S _11892_/C1 vssd1 vssd1 vccd1 vccd1
+ _11890_/X sky130_fd_sc_hd__a221o_1
XFILLER_260_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ _12309_/S _10840_/X _10839_/X _12318_/A1 vssd1 vssd1 vccd1 vccd1 _10841_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13560_ _20921_/Q _13598_/A2 _13575_/C _13559_/Y _14110_/A vssd1 vssd1 vccd1 vccd1
+ _13560_/X sky130_fd_sc_hd__a221o_1
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10772_ _12337_/A _20499_/Q _12339_/S0 _20531_/Q vssd1 vssd1 vccd1 vccd1 _10772_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_241_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12511_ _19168_/Q _12511_/B vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__or2_2
X_13491_ _13489_/X _13490_/Y _13552_/A _13488_/X vssd1 vssd1 vccd1 vccd1 _13491_/X
+ sky130_fd_sc_hd__o211a_2
X_15230_ _19706_/Q _15475_/A2 _15475_/B1 _19738_/Q vssd1 vssd1 vccd1 vccd1 _15230_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12442_ _13178_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _12450_/B sky130_fd_sc_hd__or2_1
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15161_ _15161_/A vssd1 vssd1 vccd1 vccd1 _15161_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12373_ _11336_/A _12372_/X _12371_/X vssd1 vssd1 vccd1 vccd1 _12373_/X sky130_fd_sc_hd__o21a_1
XFILLER_193_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14112_ _14112_/A _14112_/B _14112_/C vssd1 vssd1 vccd1 vccd1 _17952_/B sky130_fd_sc_hd__and3_1
X_11324_ _10804_/Y _11319_/X _11323_/Y _10805_/Y vssd1 vssd1 vccd1 vccd1 _11774_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092_ _19703_/Q _15091_/X _15395_/S vssd1 vssd1 vccd1 vccd1 _15092_/X sky130_fd_sc_hd__mux2_2
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043_ _13897_/A _14043_/A2 _14043_/B1 _14042_/X _16129_/B1 vssd1 vssd1 vccd1 vccd1
+ _19181_/D sky130_fd_sc_hd__o221a_1
XFILLER_181_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18920_ _18975_/A _18920_/B vssd1 vssd1 vccd1 vccd1 _18920_/Y sky130_fd_sc_hd__nand2_2
XFILLER_113_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11255_ _20365_/Q _20429_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _11255_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10206_ _10201_/X _10205_/X _10127_/A vssd1 vssd1 vccd1 vccd1 _10206_/Y sky130_fd_sc_hd__o21ai_2
X_18851_ _18968_/A _18851_/B vssd1 vssd1 vccd1 vccd1 _18851_/Y sky130_fd_sc_hd__nand2_1
X_11186_ _11259_/S _11281_/B vssd1 vssd1 vccd1 vccd1 _11186_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17802_ _20579_/Q _17802_/A1 _17806_/S vssd1 vssd1 vccd1 vccd1 _20579_/D sky130_fd_sc_hd__mux2_1
X_10137_ _11336_/A _19443_/Q _10137_/C vssd1 vssd1 vccd1 vccd1 _10137_/X sky130_fd_sc_hd__and3_1
XFILLER_94_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18782_ _18467_/B _18840_/B _18780_/X _18781_/Y vssd1 vssd1 vccd1 vccd1 _18783_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ _20911_/Q _16043_/A2 _15994_/B1 _15993_/X _16043_/C1 vssd1 vssd1 vccd1 vccd1
+ _15994_/X sky130_fd_sc_hd__a221o_1
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17733_ _20514_/Q _17907_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20514_/D sky130_fd_sc_hd__mux2_1
XFILLER_282_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14945_ _14945_/A _14980_/C vssd1 vssd1 vccd1 vccd1 _14945_/Y sky130_fd_sc_hd__nor2_2
X_10068_ _19941_/Q _11680_/C1 _09688_/B _12071_/S vssd1 vssd1 vccd1 vccd1 _10068_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_36_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_205_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20641_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17664_ _20450_/Q _17941_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20450_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14876_ _14841_/X _14875_/X _15612_/S vssd1 vssd1 vccd1 vccd1 _14877_/B sky130_fd_sc_hd__mux2_2
X_19403_ _20694_/CLK _19403_/D vssd1 vssd1 vccd1 vccd1 _19403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16615_ _19874_/Q _17929_/A1 _16632_/S vssd1 vssd1 vccd1 vccd1 _19874_/D sky130_fd_sc_hd__mux2_1
X_13827_ _19997_/Q split1/A _13781_/X split2/A vssd1 vssd1 vccd1 vccd1 _13827_/X sky130_fd_sc_hd__a22o_4
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17595_ _20353_/Q _17906_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20353_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19334_ _20704_/CLK _19334_/D vssd1 vssd1 vccd1 vccd1 _19334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16546_ _19839_/Q _16566_/A2 _16566_/B1 input40/X vssd1 vssd1 vccd1 vccd1 _16547_/B
+ sky130_fd_sc_hd__o22a_1
X_13758_ _13680_/Y _13741_/B _13741_/Y _13681_/Y _13757_/X vssd1 vssd1 vccd1 vccd1
+ _13759_/B sky130_fd_sc_hd__o221a_4
XFILLER_188_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12709_ split6/A _12710_/B vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__and2_4
XFILLER_176_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19265_ _20812_/CLK _19265_/D vssd1 vssd1 vccd1 vccd1 _19265_/Q sky130_fd_sc_hd__dfxtp_1
X_16477_ _19786_/Q _17940_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19786_/D sky130_fd_sc_hd__mux2_1
X_13689_ _13694_/A _14878_/A _13689_/C vssd1 vssd1 vccd1 vccd1 _13689_/X sky130_fd_sc_hd__and3_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18216_ _20797_/Q _18215_/Y _18236_/S vssd1 vssd1 vccd1 vccd1 _18217_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15428_ _16133_/C _15426_/Y _15427_/X _13596_/X _15442_/A vssd1 vssd1 vccd1 vccd1
+ _15428_/X sky130_fd_sc_hd__a32o_1
X_19196_ _19704_/CLK _19196_/D vssd1 vssd1 vccd1 vccd1 _19196_/Q sky130_fd_sc_hd__dfxtp_1
X_18147_ _18157_/A _18156_/B _18156_/C vssd1 vssd1 vccd1 vccd1 _18389_/B sky130_fd_sc_hd__or3_1
XFILLER_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15359_ _15354_/Y _15358_/X _15612_/S vssd1 vssd1 vccd1 vccd1 _15359_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18078_ _18080_/A _18078_/B _18079_/B vssd1 vssd1 vccd1 vccd1 _20766_/D sky130_fd_sc_hd__nor3_1
XFILLER_132_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09920_ _19886_/Q _19787_/Q _09931_/S vssd1 vssd1 vccd1 vccd1 _09920_/X sky130_fd_sc_hd__mux2_1
X_17029_ _20007_/Q input193/X _17040_/S vssd1 vssd1 vccd1 vccd1 _20007_/D sky130_fd_sc_hd__mux2_1
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20040_ _20679_/CLK _20040_/D vssd1 vssd1 vccd1 vccd1 _20040_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout706 _16528_/Y vssd1 vssd1 vccd1 vccd1 _16566_/A2 sky130_fd_sc_hd__buf_4
XFILLER_252_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout717 _16529_/Y vssd1 vssd1 vccd1 vccd1 _16566_/B1 sky130_fd_sc_hd__buf_4
X_09851_ _20323_/Q _11708_/B vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__or2_1
Xfanout728 _13142_/X vssd1 vssd1 vccd1 vccd1 _19661_/D sky130_fd_sc_hd__buf_6
XFILLER_213_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout739 _14204_/A vssd1 vssd1 vccd1 vccd1 _14397_/A sky130_fd_sc_hd__buf_4
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09782_/A vssd1 vssd1 vccd1 vccd1 _09784_/A sky130_fd_sc_hd__clkinv_2
XFILLER_61_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _21008_/CLK _20942_/D vssd1 vssd1 vccd1 vccd1 _20942_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_226_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20873_ _21042_/CLK _20873_/D vssd1 vssd1 vccd1 vccd1 _20873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20307_ _20467_/CLK _20307_/D vssd1 vssd1 vccd1 vccd1 _20307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11040_ _11021_/A _19337_/Q _20692_/Q _11039_/S _11378_/S vssd1 vssd1 vccd1 vccd1
+ _11040_/X sky130_fd_sc_hd__a221o_1
XFILLER_150_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20238_ _20969_/CLK _20238_/D vssd1 vssd1 vccd1 vccd1 _20238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_276_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20169_ _20708_/CLK _20169_/D vssd1 vssd1 vccd1 vccd1 _20169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12991_ _19233_/Q _19224_/Q _13587_/B _12991_/D vssd1 vssd1 vccd1 vccd1 _13296_/B
+ sky130_fd_sc_hd__and4_2
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11942_ _09776_/S _11937_/Y _11941_/Y _12020_/C1 vssd1 vssd1 vccd1 vccd1 _11942_/X
+ sky130_fd_sc_hd__a211o_1
X_14730_ _19487_/Q _17911_/A1 _14732_/S vssd1 vssd1 vccd1 vccd1 _19487_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_600 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_611 _12426_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_622 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _19423_/Q _17805_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19423_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_633 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ _09839_/A _11855_/X _11872_/X vssd1 vssd1 vccd1 vccd1 _11873_/X sky130_fd_sc_hd__o21a_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_644 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_655 input241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16400_ _19745_/Q _16402_/C _16399_/Y vssd1 vssd1 vccd1 vccd1 _19745_/D sky130_fd_sc_hd__o21a_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13612_ _13612_/A _15442_/B vssd1 vssd1 vccd1 vccd1 _13612_/X sky130_fd_sc_hd__and2_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _19934_/Q _12213_/B vssd1 vssd1 vccd1 vccd1 _10824_/X sky130_fd_sc_hd__or2_1
XFILLER_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14592_ _19358_/Q _17944_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19358_/D sky130_fd_sc_hd__mux2_1
X_17380_ _20238_/Q _17390_/A2 _17382_/B1 _20287_/Q _17380_/C1 vssd1 vssd1 vccd1 vccd1
+ _17380_/X sky130_fd_sc_hd__a221o_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16331_ _18821_/A _16331_/B _16332_/B vssd1 vssd1 vccd1 vccd1 _19719_/D sky130_fd_sc_hd__nor3_1
X_13543_ _13544_/A _13544_/B vssd1 vssd1 vccd1 vccd1 _13543_/X sky130_fd_sc_hd__or2_1
XFILLER_111_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10755_ _19804_/Q _19308_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10755_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19050_ _21044_/Q _14112_/A _19050_/S vssd1 vssd1 vccd1 vccd1 _19051_/B sky130_fd_sc_hd__mux2_1
X_16262_ _19678_/Q _17202_/A1 _16274_/S vssd1 vssd1 vccd1 vccd1 _19678_/D sky130_fd_sc_hd__mux2_1
X_13474_ _13462_/B split2/A split1/A _20006_/Q vssd1 vssd1 vccd1 vccd1 _13474_/X sky130_fd_sc_hd__a22o_4
X_10686_ _10692_/A _19904_/Q _12272_/B2 _20029_/Q vssd1 vssd1 vccd1 vccd1 _10686_/X
+ sky130_fd_sc_hd__o22a_1
X_18001_ _20738_/Q _18003_/C _18000_/Y vssd1 vssd1 vccd1 vccd1 _20738_/D sky130_fd_sc_hd__o21a_1
X_15213_ _14817_/X _14855_/X _15357_/S vssd1 vssd1 vccd1 vccd1 _15214_/B sky130_fd_sc_hd__mux2_1
X_12425_ _20148_/Q _20116_/Q _12428_/S vssd1 vssd1 vccd1 vccd1 _12425_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16193_ _16193_/A _16193_/B vssd1 vssd1 vccd1 vccd1 _19620_/D sky130_fd_sc_hd__and2_1
XFILLER_275_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15144_ _17245_/A _15143_/X _15452_/S vssd1 vssd1 vccd1 vccd1 _15144_/X sky130_fd_sc_hd__mux2_2
X_12356_ _12411_/A _20396_/Q _20460_/Q _12352_/S vssd1 vssd1 vccd1 vccd1 _12356_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_275_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput309 _13616_/X vssd1 vssd1 vccd1 vccd1 core_wb_adr_o[13] sky130_fd_sc_hd__buf_4
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11307_ _10356_/A _20365_/Q _20429_/Q _11295_/S vssd1 vssd1 vccd1 vccd1 _11307_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15075_ _15075_/A _15075_/B vssd1 vssd1 vccd1 vccd1 _15075_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19952_ _20480_/CLK _19952_/D vssd1 vssd1 vccd1 vccd1 _19952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12287_ _12288_/B _12288_/C _12288_/A vssd1 vssd1 vccd1 vccd1 _12290_/C sky130_fd_sc_hd__a21oi_1
X_14026_ _14035_/A1 _14038_/A2 _10467_/X _14038_/B1 _19857_/Q vssd1 vssd1 vccd1 vccd1
+ _14097_/C sky130_fd_sc_hd__o32a_1
X_18903_ _21000_/Q _18964_/B vssd1 vssd1 vccd1 vccd1 _18903_/Y sky130_fd_sc_hd__nand2_1
X_11238_ input107/X input132/X _19694_/Q vssd1 vssd1 vccd1 vccd1 _11238_/X sky130_fd_sc_hd__mux2_8
XFILLER_45_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19883_ _20081_/CLK _19883_/D vssd1 vssd1 vccd1 vccd1 _19883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18834_ _18496_/X _18861_/B _18832_/X _18833_/Y vssd1 vssd1 vccd1 vccd1 _18835_/B
+ sky130_fd_sc_hd__o211a_1
X_11169_ _20151_/Q _11169_/B vssd1 vssd1 vccd1 vccd1 _11169_/X sky130_fd_sc_hd__or2_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18765_ _18765_/A _18765_/B _18765_/C _18765_/D vssd1 vssd1 vccd1 vccd1 _18811_/S
+ sky130_fd_sc_hd__or4_4
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15977_ _15977_/A1 _12902_/Y _15976_/X _16062_/B2 vssd1 vssd1 vccd1 vccd1 _15979_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ _20497_/Q _17750_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20497_/D sky130_fd_sc_hd__mux2_1
X_14928_ _14119_/A _12584_/C _18148_/S vssd1 vssd1 vccd1 vccd1 _14955_/B sky130_fd_sc_hd__mux2_8
XFILLER_208_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18696_ _18783_/A _18696_/B vssd1 vssd1 vccd1 vccd1 _20948_/D sky130_fd_sc_hd__nor2_1
XFILLER_282_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17647_ _20433_/Q _17647_/A1 _17657_/S vssd1 vssd1 vccd1 vccd1 _20433_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14859_ _14857_/X _14858_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _14859_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17578_ _20336_/Q _17889_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20336_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19317_ _20692_/CLK _19317_/D vssd1 vssd1 vccd1 vccd1 _19317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16529_ _19863_/Q input9/X _16594_/B _19864_/Q vssd1 vssd1 vccd1 vccd1 _16529_/Y
+ sky130_fd_sc_hd__nand4b_4
XFILLER_188_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ _20268_/CLK _19248_/D vssd1 vssd1 vccd1 vccd1 _19248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19179_ _20426_/CLK _19179_/D vssd1 vssd1 vccd1 vccd1 _19179_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_247_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09903_ _12144_/C1 _09892_/X _09895_/X _09902_/X _12152_/A1 vssd1 vssd1 vccd1 vccd1
+ _09903_/X sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_198_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20649_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout503 _17813_/X vssd1 vssd1 vccd1 vccd1 _17844_/S sky130_fd_sc_hd__buf_6
XFILLER_160_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout514 _17711_/X vssd1 vssd1 vccd1 vccd1 _17743_/S sky130_fd_sc_hd__buf_12
XFILLER_59_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_258_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout525 _17608_/X vssd1 vssd1 vccd1 vccd1 _17635_/S sky130_fd_sc_hd__buf_6
XFILLER_259_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout536 _17212_/S vssd1 vssd1 vccd1 vccd1 _17214_/S sky130_fd_sc_hd__buf_8
X_20023_ _20341_/CLK _20023_/D vssd1 vssd1 vccd1 vccd1 _20023_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout547 _17117_/X vssd1 vssd1 vccd1 vccd1 _17144_/S sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_127_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21022_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09834_ _09834_/A _20679_/Q _09834_/C vssd1 vssd1 vccd1 vccd1 _09834_/X sky130_fd_sc_hd__or3_1
XFILLER_258_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout558 _16673_/X vssd1 vssd1 vccd1 vccd1 _16705_/S sky130_fd_sc_hd__buf_12
Xfanout569 _16490_/X vssd1 vssd1 vccd1 vccd1 _16517_/S sky130_fd_sc_hd__buf_6
XFILLER_59_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09765_ _09752_/A _20388_/Q _20452_/Q _11936_/S _12016_/C1 vssd1 vssd1 vccd1 vccd1
+ _09765_/X sky130_fd_sc_hd__a221o_1
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_273_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_273_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09696_ _11514_/A1 _11983_/A1 _19357_/Q _12129_/S vssd1 vssd1 vccd1 vccd1 _09696_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ _21023_/CLK _20925_/D vssd1 vssd1 vccd1 vccd1 _20925_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20856_ _20856_/CLK _20856_/D vssd1 vssd1 vccd1 vccd1 _20856_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20787_ _20861_/CLK _20787_/D vssd1 vssd1 vccd1 vccd1 _20787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10540_ _10540_/A _10540_/B _10641_/B vssd1 vssd1 vccd1 vccd1 _10540_/X sky130_fd_sc_hd__and3_1
XFILLER_211_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ _10037_/Y _10470_/Y _09669_/X vssd1 vssd1 vccd1 vccd1 _10471_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12210_ _10385_/A _12209_/X _12208_/X vssd1 vssd1 vccd1 vccd1 _12210_/X sky130_fd_sc_hd__a21o_4
XFILLER_182_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13190_ _13481_/A _17041_/B vssd1 vssd1 vccd1 vccd1 _16594_/B sky130_fd_sc_hd__nand2b_4
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12141_ _20425_/Q _20361_/Q _12148_/S vssd1 vssd1 vccd1 vccd1 _12141_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12072_ _12072_/A1 _12071_/X _12068_/X _12072_/C1 vssd1 vssd1 vccd1 vccd1 _12072_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11023_ _19626_/Q _19932_/Q _19270_/Q _20057_/Q _11292_/S0 _11290_/C vssd1 vssd1
+ vccd1 vccd1 _11023_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15900_ _12111_/B _12466_/Y _12468_/X _12109_/Y _15365_/A vssd1 vssd1 vccd1 vccd1
+ _15900_/X sky130_fd_sc_hd__o221a_1
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16880_ _20413_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16880_/X sky130_fd_sc_hd__a21o_2
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_265_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_277_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _16017_/C1 _15830_/X _15826_/X vssd1 vssd1 vccd1 vccd1 _15831_/X sky130_fd_sc_hd__o21a_2
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_265_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _18651_/B _18550_/B vssd1 vssd1 vccd1 vccd1 _18550_/X sky130_fd_sc_hd__or2_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15762_ _15762_/A _15925_/B vssd1 vssd1 vccd1 vccd1 _15762_/Y sky130_fd_sc_hd__nand2_1
X_12974_ _19109_/Q _12974_/B _19112_/Q vssd1 vssd1 vccd1 vccd1 _12975_/D sky130_fd_sc_hd__or3b_4
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _17505_/A1 _17500_/Y _18112_/A vssd1 vssd1 vccd1 vccd1 _20285_/D sky130_fd_sc_hd__a21oi_1
X_14713_ _19470_/Q _17928_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19470_/D sky130_fd_sc_hd__mux2_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18481_ _20887_/Q fanout753/X _18480_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18482_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _12003_/A _19327_/Q _12003_/C vssd1 vssd1 vccd1 vccd1 _11925_/X sky130_fd_sc_hd__or3_1
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15693_ _20932_/Q _15995_/A2 _15692_/X vssd1 vssd1 vccd1 vccd1 _15693_/X sky130_fd_sc_hd__o21a_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_430 _13242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_441 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_452 _14522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17432_ _17432_/A _17432_/B vssd1 vssd1 vccd1 vccd1 _20260_/D sky130_fd_sc_hd__and2_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14644_ _19406_/Q _17788_/A1 _14650_/S vssd1 vssd1 vccd1 vccd1 _19406_/D sky130_fd_sc_hd__mux2_1
X_11856_ _20142_/Q _20110_/Q _11944_/S vssd1 vssd1 vccd1 vccd1 _11856_/X sky130_fd_sc_hd__mux2_1
XANTENNA_463 _19171_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_474 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_485 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10807_ _10373_/A _10119_/Y _09659_/B vssd1 vssd1 vccd1 vccd1 _10807_/X sky130_fd_sc_hd__a21o_1
XANTENNA_496 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14575_ _19341_/Q _17927_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19341_/D sky130_fd_sc_hd__mux2_1
X_17363_ _20230_/Q _17363_/A2 _17362_/X _18396_/A vssd1 vssd1 vccd1 vccd1 _20230_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11787_ _11787_/A _15259_/A _15221_/A _11786_/X vssd1 vssd1 vccd1 vccd1 _11788_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19102_ _19609_/CLK _19102_/D vssd1 vssd1 vccd1 vccd1 _19102_/Q sky130_fd_sc_hd__dfxtp_2
X_16314_ _19712_/Q _19713_/Q _16314_/C vssd1 vssd1 vccd1 vccd1 _16316_/B sky130_fd_sc_hd__and3_1
X_10738_ _10734_/X _10737_/X _12302_/S vssd1 vssd1 vccd1 vccd1 _10738_/X sky130_fd_sc_hd__mux2_1
X_13526_ _13526_/A _13526_/B _13526_/C vssd1 vssd1 vccd1 vccd1 _13526_/X sky130_fd_sc_hd__or3_1
XFILLER_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17294_ _20203_/Q _17327_/A2 _17330_/C1 vssd1 vssd1 vccd1 vccd1 _17294_/X sky130_fd_sc_hd__a21o_1
X_19033_ _21035_/Q _19049_/A2 _19032_/X _18740_/A vssd1 vssd1 vccd1 vccd1 _21035_/D
+ sky130_fd_sc_hd__o211a_1
X_16245_ _17745_/A _17676_/B _16245_/C vssd1 vssd1 vccd1 vccd1 _16245_/X sky130_fd_sc_hd__and3_2
XFILLER_158_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13457_ _13452_/Y _13456_/X _14275_/A1 vssd1 vssd1 vccd1 vccd1 _13457_/X sky130_fd_sc_hd__o21a_1
X_10669_ _19373_/Q _20664_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10669_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12408_ _19653_/Q _19959_/Q _19297_/Q _20084_/Q _11116_/S _12406_/C vssd1 vssd1 vccd1
+ vccd1 _12408_/X sky130_fd_sc_hd__mux4_1
X_16176_ _19612_/Q _15780_/X _16190_/S vssd1 vssd1 vccd1 vccd1 _16177_/B sky130_fd_sc_hd__mux2_1
X_13388_ _13388_/A _13388_/B _13388_/C _13388_/D vssd1 vssd1 vccd1 vccd1 _13412_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12339_ _20428_/Q _20364_/Q _20656_/Q _20620_/Q _12339_/S0 _12254_/C vssd1 vssd1
+ vccd1 vccd1 _12339_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15127_ _15127_/A _15127_/B vssd1 vssd1 vccd1 vccd1 _15127_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19935_ _20061_/CLK _19935_/D vssd1 vssd1 vccd1 vccd1 _19935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15058_ _14812_/X _14821_/X _15058_/S vssd1 vssd1 vccd1 vccd1 _15158_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _19202_/Q _14085_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _14009_/X sky130_fd_sc_hd__mux2_1
X_19866_ _20638_/CLK _19866_/D vssd1 vssd1 vccd1 vccd1 _19866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18817_ _19125_/Q _12533_/B _18880_/B1 vssd1 vssd1 vccd1 vccd1 _18817_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19797_ _20155_/CLK _19797_/D vssd1 vssd1 vccd1 vccd1 _19797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09550_ _12464_/A _11268_/C vssd1 vssd1 vccd1 vccd1 _12468_/C sky130_fd_sc_hd__nand2_8
X_18748_ _18748_/A _18748_/B vssd1 vssd1 vccd1 vccd1 _20974_/D sky130_fd_sc_hd__and2_1
XFILLER_209_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09481_ _20882_/Q vssd1 vssd1 vccd1 vccd1 _09481_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18679_ _19523_/Q _18687_/B vssd1 vssd1 vccd1 vccd1 _18679_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20710_ _20710_/CLK _20710_/D vssd1 vssd1 vccd1 vccd1 _20710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20641_ _20641_/CLK _20641_/D vssd1 vssd1 vccd1 vccd1 _20641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20572_ _20702_/CLK _20572_/D vssd1 vssd1 vccd1 vccd1 _20572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1309 _14836_/S vssd1 vssd1 vccd1 vccd1 _14843_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20006_ _20751_/CLK _20006_/D vssd1 vssd1 vccd1 vccd1 _20006_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09817_ _19820_/Q _19324_/Q _12070_/S vssd1 vssd1 vccd1 vccd1 _09817_/X sky130_fd_sc_hd__mux2_1
XFILLER_247_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09748_ _09748_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09748_/Y sky130_fd_sc_hd__nor2_4
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09679_ _09676_/A _09676_/B _10373_/A vssd1 vssd1 vccd1 vccd1 _09679_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_95_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20428_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _19784_/Q _11718_/S _10622_/S _12023_/S vssd1 vssd1 vccd1 vccd1 _11710_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ _21006_/CLK _20908_/D vssd1 vssd1 vccd1 vccd1 _20908_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _13526_/A _12692_/D vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__nor2_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i _20408_/CLK vssd1 vssd1 vccd1 vccd1 _20668_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11639_/X _11640_/X _11641_/S vssd1 vssd1 vccd1 vccd1 _11641_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20839_ _20969_/CLK _20839_/D vssd1 vssd1 vccd1 vccd1 _20839_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14360_ _19238_/Q _14438_/A2 _14359_/X _18752_/A vssd1 vssd1 vccd1 vccd1 _19238_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11572_ _11574_/A _11735_/B vssd1 vssd1 vccd1 vccd1 _11575_/A sky130_fd_sc_hd__nor2_2
XFILLER_122_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13311_ _19227_/Q _13450_/A vssd1 vssd1 vccd1 vccd1 _13311_/X sky130_fd_sc_hd__or2_1
X_10523_ _10520_/X _10521_/X _10522_/X _09507_/A _12514_/C vssd1 vssd1 vccd1 vccd1
+ _10523_/X sky130_fd_sc_hd__a221o_1
Xinput19 core_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ _14303_/A _14302_/A vssd1 vssd1 vccd1 vccd1 _14293_/A sky130_fd_sc_hd__or2_1
XFILLER_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13242_ _13242_/A _13242_/B _13242_/C _13242_/D vssd1 vssd1 vccd1 vccd1 _13242_/X
+ sky130_fd_sc_hd__or4_2
X_16030_ _15983_/A _15066_/X _16025_/Y _16027_/X _16030_/D1 vssd1 vssd1 vccd1 vccd1
+ _16030_/X sky130_fd_sc_hd__a2111o_1
XFILLER_109_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10454_ _10640_/B _10455_/B vssd1 vssd1 vccd1 vccd1 _10456_/B sky130_fd_sc_hd__nand2_1
XFILLER_183_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13173_ _11961_/B _13433_/B _15887_/S vssd1 vssd1 vccd1 vccd1 _13432_/B sky130_fd_sc_hd__a21oi_4
XFILLER_124_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10385_ _10385_/A _10385_/B vssd1 vssd1 vccd1 vccd1 _10385_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _19426_/Q _20585_/Q _12124_/S vssd1 vssd1 vccd1 vccd1 _12124_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17981_ _20731_/Q _17982_/C _17980_/Y vssd1 vssd1 vccd1 vccd1 _20731_/D sky130_fd_sc_hd__o21a_1
XFILLER_269_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19720_ _21026_/CLK _19720_/D vssd1 vssd1 vccd1 vccd1 _19720_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1810 _19527_/Q vssd1 vssd1 vccd1 vccd1 _11235_/A sky130_fd_sc_hd__buf_6
X_16932_ _16932_/A1 _16931_/X _16932_/B1 vssd1 vssd1 vccd1 vccd1 _16932_/Y sky130_fd_sc_hd__o21ai_2
X_12055_ _12045_/X _12047_/X _12054_/X _12058_/S _12136_/B1 vssd1 vssd1 vccd1 vccd1
+ _12055_/X sky130_fd_sc_hd__o221a_1
Xfanout1821 _19176_/Q vssd1 vssd1 vccd1 vccd1 _12513_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_2_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1832 _12136_/B1 vssd1 vssd1 vccd1 vccd1 _12137_/A1 sky130_fd_sc_hd__buf_6
XFILLER_78_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1843 _19171_/Q vssd1 vssd1 vccd1 vccd1 _12125_/A1 sky130_fd_sc_hd__buf_8
XFILLER_266_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11006_ _19626_/Q _11009_/A2 _11003_/X _11004_/X _11005_/X vssd1 vssd1 vccd1 vccd1
+ _11006_/X sky130_fd_sc_hd__o221a_1
XFILLER_120_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19651_ _20075_/CLK _19651_/D vssd1 vssd1 vccd1 vccd1 _19651_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1854 _12828_/A vssd1 vssd1 vccd1 vccd1 _09776_/S sky130_fd_sc_hd__buf_6
Xfanout1865 _12504_/A vssd1 vssd1 vccd1 vccd1 _11384_/S sky130_fd_sc_hd__buf_8
X_16863_ _16805_/X _16860_/Y _16862_/X _16974_/A1 vssd1 vssd1 vccd1 vccd1 _16863_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1876 _09731_/A vssd1 vssd1 vccd1 vccd1 _12357_/A1 sky130_fd_sc_hd__buf_6
XFILLER_65_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1887 _14802_/C1 vssd1 vssd1 vccd1 vccd1 _17536_/D sky130_fd_sc_hd__buf_2
X_18602_ _18856_/A _18602_/B vssd1 vssd1 vccd1 vccd1 _20923_/D sky130_fd_sc_hd__nor2_1
Xfanout1898 fanout1905/X vssd1 vssd1 vccd1 vccd1 _18736_/A sky130_fd_sc_hd__clkbuf_2
X_15814_ _15814_/A _15814_/B _15814_/C vssd1 vssd1 vccd1 vccd1 _15814_/Y sky130_fd_sc_hd__nand3_1
X_19582_ _19589_/CLK _19582_/D vssd1 vssd1 vccd1 vccd1 _19582_/Q sky130_fd_sc_hd__dfxtp_1
X_16794_ _16869_/A _16794_/B vssd1 vssd1 vccd1 vccd1 _16794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18533_ _20904_/Q fanout750/X _18532_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18534_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_218_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _20870_/Q _16018_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15745_/X sky130_fd_sc_hd__o21ba_1
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _19252_/Q _12964_/A2 _16716_/A _20000_/Q vssd1 vssd1 vccd1 vccd1 _16719_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18464_ _20883_/Q fanout753/X _18463_/X _18509_/B2 vssd1 vssd1 vccd1 vccd1 _18464_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_11908_ _11917_/S _11907_/X _11906_/X _12151_/A1 vssd1 vssd1 vccd1 vccd1 _11908_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_221_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15676_ _15977_/A1 _12846_/Y _15675_/X _15703_/B2 vssd1 vssd1 vccd1 vccd1 _15676_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12888_ _19519_/Q _12884_/B _19520_/Q vssd1 vssd1 vccd1 vccd1 _12889_/B sky130_fd_sc_hd__a21oi_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_271 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_282 _20624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17415_ _17402_/A _17441_/A _17457_/B _20254_/Q vssd1 vssd1 vccd1 vccd1 _17415_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14627_ _19391_/Q _17911_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19391_/D sky130_fd_sc_hd__mux2_1
XANTENNA_293 input223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18395_ _20852_/Q _18170_/Y _18395_/S vssd1 vssd1 vccd1 vccd1 _18396_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11839_ _12140_/C1 _11838_/X _11835_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _11839_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17346_ _20221_/Q _17364_/A2 _17370_/B1 _20270_/Q _17370_/C1 vssd1 vssd1 vccd1 vccd1
+ _17346_/X sky130_fd_sc_hd__a221o_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14558_ _19328_/Q _17178_/A1 _14558_/S vssd1 vssd1 vccd1 vccd1 _19328_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13509_ _16241_/A _13909_/A vssd1 vssd1 vccd1 vccd1 _13509_/Y sky130_fd_sc_hd__nor2_1
X_17277_ _20198_/Q _17280_/A2 _17276_/X _17331_/C1 vssd1 vssd1 vccd1 vccd1 _20198_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14489_ _19267_/Q _17886_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19267_/D sky130_fd_sc_hd__mux2_1
X_19016_ _18235_/Y _18982_/B _19016_/B1 _19015_/X vssd1 vssd1 vccd1 vccd1 _21027_/D
+ sky130_fd_sc_hd__o211a_1
X_16228_ _19651_/Q _17705_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19651_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16159_ _19603_/Q _16178_/S _16158_/Y _16159_/C1 vssd1 vssd1 vccd1 vccd1 _19603_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19918_ _20446_/CLK _19918_/D vssd1 vssd1 vccd1 vccd1 _19918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19849_ _19970_/CLK _19849_/D vssd1 vssd1 vccd1 vccd1 _19849_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09602_ _09609_/A _19093_/Q vssd1 vssd1 vccd1 vccd1 _17709_/C sky130_fd_sc_hd__nand2b_4
XFILLER_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09533_ _19526_/Q _19149_/Q vssd1 vssd1 vccd1 vccd1 _09533_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_243_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20624_ _20624_/CLK _20624_/D vssd1 vssd1 vccd1 vccd1 _20624_/Q sky130_fd_sc_hd__dfxtp_4
X_20555_ _20655_/CLK _20555_/D vssd1 vssd1 vccd1 vccd1 _20555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20486_ _20714_/CLK _20486_/D vssd1 vssd1 vccd1 vccd1 _20486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_142_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19505_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_279_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10170_ _19675_/Q _20163_/Q _12428_/S vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__mux2_1
XFILLER_279_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput470 _19522_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[28] sky130_fd_sc_hd__buf_4
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput481 _19503_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[9] sky130_fd_sc_hd__buf_4
Xfanout1106 _17913_/A1 vssd1 vssd1 vccd1 vccd1 _17111_/A1 sky130_fd_sc_hd__buf_4
XFILLER_248_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1117 _17870_/A1 vssd1 vssd1 vccd1 vccd1 _17938_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_248_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1128 _17592_/A1 vssd1 vssd1 vccd1 vccd1 _17869_/A1 sky130_fd_sc_hd__buf_4
XFILLER_87_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1139 _09947_/X vssd1 vssd1 vccd1 vccd1 _17906_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_259_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21038_ _21041_/CLK _21038_/D vssd1 vssd1 vccd1 vccd1 _21038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13860_ _16066_/B _13860_/B _13860_/C vssd1 vssd1 vccd1 vccd1 _13860_/X sky130_fd_sc_hd__or3_2
XFILLER_270_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _12811_/A _12811_/B vssd1 vssd1 vccd1 vccd1 _12811_/X sky130_fd_sc_hd__or2_1
XFILLER_250_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13791_ _13798_/A1 _13826_/A1 _13666_/B _13826_/B1 input215/X vssd1 vssd1 vccd1 vccd1
+ _13791_/X sky130_fd_sc_hd__a32o_2
XFILLER_234_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15530_ _19715_/Q _15595_/A2 _15595_/B1 _19747_/Q vssd1 vssd1 vccd1 vccd1 _15530_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ split8/A _12847_/A2 _15526_/A _12741_/Y vssd1 vssd1 vccd1 vccd1 _12742_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12673_ _12498_/A _12498_/B _12495_/Y vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__o21ai_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15461_ _10509_/Y _15460_/X _15591_/A vssd1 vssd1 vccd1 vccd1 _15461_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_203_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17200_ _20164_/Q _17657_/A1 _17215_/S vssd1 vssd1 vccd1 vccd1 _20164_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _19523_/Q _14413_/B vssd1 vssd1 vccd1 vccd1 _14426_/A sky130_fd_sc_hd__nor2_1
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11624_ _12003_/A _20544_/Q _20512_/Q _11932_/S0 vssd1 vssd1 vccd1 vccd1 _11624_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_230_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18180_ _18477_/B vssd1 vssd1 vccd1 vccd1 _18180_/Y sky130_fd_sc_hd__clkinv_2
X_15392_ _17296_/A _15482_/A2 _15390_/X _15391_/X vssd1 vssd1 vccd1 vccd1 _15392_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_230_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17131_ _20099_/Q _17199_/A1 _17149_/S vssd1 vssd1 vccd1 vccd1 _20099_/D sky130_fd_sc_hd__mux2_1
XFILLER_156_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14343_ _14343_/A _14343_/B _14343_/C vssd1 vssd1 vccd1 vccd1 _14345_/B sky130_fd_sc_hd__and3_1
X_11555_ _19782_/Q _11563_/S _09931_/S _11945_/S vssd1 vssd1 vccd1 vccd1 _11555_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10506_ _13675_/A _13675_/B _13675_/C _11368_/A1 vssd1 vssd1 vccd1 vccd1 _10540_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14274_ _14269_/B _14273_/Y _14417_/S vssd1 vssd1 vccd1 vccd1 _14274_/X sky130_fd_sc_hd__mux2_1
X_17062_ _20034_/Q _17096_/A1 _17076_/S vssd1 vssd1 vccd1 vccd1 _20034_/D sky130_fd_sc_hd__mux2_1
X_11486_ _11849_/S _11483_/X _11485_/X _12183_/C1 vssd1 vssd1 vccd1 vccd1 _11486_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16013_ _21042_/Q _21010_/Q _16040_/S vssd1 vssd1 vccd1 vccd1 _16013_/X sky130_fd_sc_hd__mux2_1
X_13225_ _13350_/A _13209_/C _13221_/X _13224_/X vssd1 vssd1 vccd1 vccd1 _13229_/B
+ sky130_fd_sc_hd__a31o_1
X_10437_ _10581_/A1 _20668_/Q _12068_/C1 _10585_/S vssd1 vssd1 vccd1 vccd1 _10437_/X
+ sky130_fd_sc_hd__o31a_1
X_13156_ _10456_/A _13155_/A _13155_/B _10455_/B _15473_/A vssd1 vssd1 vccd1 vccd1
+ _13425_/B sky130_fd_sc_hd__a32o_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _13425_/A _13424_/A _13422_/A _13423_/A vssd1 vssd1 vccd1 vccd1 _11409_/A
+ sky130_fd_sc_hd__and4_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12107_ _12107_/A1 _17878_/A1 _12106_/X _12194_/B2 vssd1 vssd1 vccd1 vccd1 _15904_/A
+ sky130_fd_sc_hd__a22o_4
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17964_ _17965_/B _17964_/B vssd1 vssd1 vccd1 vccd1 _20725_/D sky130_fd_sc_hd__nor2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13086_/A _13227_/A _13011_/Y _13012_/X vssd1 vssd1 vccd1 vccd1 _13216_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10299_ _11259_/S _19444_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _10299_/X sky130_fd_sc_hd__and3_1
X_19703_ _21044_/CLK _19703_/D vssd1 vssd1 vccd1 vccd1 _19703_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_238_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1640 _17502_/B vssd1 vssd1 vccd1 vccd1 _17524_/B sky130_fd_sc_hd__clkbuf_4
X_12038_ _19553_/Q _12155_/A2 _12155_/B1 _19617_/Q vssd1 vssd1 vccd1 vccd1 _12038_/X
+ sky130_fd_sc_hd__a22o_2
X_16915_ _16981_/A1 _15753_/X _16879_/X _16914_/X vssd1 vssd1 vccd1 vccd1 _16915_/X
+ sky130_fd_sc_hd__o211a_2
Xfanout1651 _09670_/Y vssd1 vssd1 vccd1 vccd1 _14011_/A2 sky130_fd_sc_hd__buf_6
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17895_ _20666_/Q _17895_/A1 _17912_/S vssd1 vssd1 vccd1 vccd1 _20666_/D sky130_fd_sc_hd__mux2_1
Xfanout1662 _12464_/C vssd1 vssd1 vccd1 vccd1 _11268_/C sky130_fd_sc_hd__clkbuf_16
Xfanout1673 _11228_/A1 vssd1 vssd1 vccd1 vccd1 _11242_/A1 sky130_fd_sc_hd__buf_8
XFILLER_226_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_254_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19634_ _20669_/CLK _19634_/D vssd1 vssd1 vccd1 vccd1 _19634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1684 _12711_/A vssd1 vssd1 vccd1 vccd1 _12102_/A1 sky130_fd_sc_hd__buf_6
Xfanout1695 _12254_/A vssd1 vssd1 vccd1 vccd1 _12427_/A1 sky130_fd_sc_hd__buf_6
X_16846_ _16846_/A input81/X vssd1 vssd1 vccd1 vccd1 _16846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_280_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19565_ _19574_/CLK _19565_/D vssd1 vssd1 vccd1 vccd1 _19565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16777_ _19220_/Q _16996_/A2 _16713_/X _16774_/Y _16776_/X vssd1 vssd1 vccd1 vccd1
+ _16777_/X sky130_fd_sc_hd__o2111a_1
XFILLER_81_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13989_ _19163_/Q _14031_/A2 _14040_/B1 _13988_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1
+ _19163_/D sky130_fd_sc_hd__o221a_1
XFILLER_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18516_ _18891_/A _18516_/B vssd1 vssd1 vccd1 vccd1 _20898_/D sky130_fd_sc_hd__nor2_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15728_ _16024_/A1 _15726_/X _15727_/Y _13428_/C _15975_/B2 vssd1 vssd1 vccd1 vccd1
+ _15728_/X sky130_fd_sc_hd__a32o_1
XFILLER_206_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19496_ _19505_/CLK _19496_/D vssd1 vssd1 vccd1 vccd1 _19496_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_209_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18447_ _20878_/Q _18300_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18448_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15659_ _15659_/A _16009_/B vssd1 vssd1 vccd1 vccd1 _15659_/X sky130_fd_sc_hd__and2_1
XFILLER_178_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18378_ _20844_/Q _18387_/B _18377_/Y _18754_/A vssd1 vssd1 vccd1 vccd1 _20844_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17329_ input8/X input283/X _17329_/S vssd1 vssd1 vccd1 vccd1 _17329_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20340_ _20655_/CLK _20340_/D vssd1 vssd1 vccd1 vccd1 _20340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_1__f_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19552_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20271_ _20818_/CLK _20271_/D vssd1 vssd1 vccd1 vccd1 _20271_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_255_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput209 localMemory_wb_adr_i[5] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09516_ _19660_/Q vssd1 vssd1 vccd1 vccd1 _09516_/Y sky130_fd_sc_hd__inv_6
XFILLER_213_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20607_ _20675_/CLK _20607_/D vssd1 vssd1 vccd1 vccd1 _20607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11340_ _12371_/A1 _19342_/Q _20697_/Q _11342_/S _12304_/C1 vssd1 vssd1 vccd1 vccd1
+ _11340_/X sky130_fd_sc_hd__a221o_1
X_20538_ _20638_/CLK _20538_/D vssd1 vssd1 vccd1 vccd1 _20538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11271_ _19623_/Q _09689_/D _11268_/X _11269_/X _11270_/X vssd1 vssd1 vccd1 vccd1
+ _11275_/B sky130_fd_sc_hd__o221a_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20469_ _20718_/CLK _20469_/D vssd1 vssd1 vccd1 vccd1 _20469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13010_ _20974_/Q _20908_/Q vssd1 vssd1 vccd1 vccd1 _13120_/B sky130_fd_sc_hd__nand2_1
X_10222_ _11345_/S _10210_/X _10214_/X _12310_/C1 vssd1 vssd1 vccd1 vccd1 _10222_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10153_ _09623_/B _10152_/X _10149_/X _11275_/A vssd1 vssd1 vccd1 vccd1 _10153_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_181_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14961_ _15019_/C _15014_/D vssd1 vssd1 vccd1 vccd1 _15021_/B sky130_fd_sc_hd__and2_4
X_10084_ _20473_/Q _11305_/B _09507_/A vssd1 vssd1 vccd1 vccd1 _10084_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16700_ _19955_/Q _17178_/A1 _16701_/S vssd1 vssd1 vccd1 vccd1 _19955_/D sky130_fd_sc_hd__mux2_1
XFILLER_236_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13912_ _19121_/Q _13919_/S _13911_/Y _14758_/C1 vssd1 vssd1 vccd1 vccd1 _19121_/D
+ sky130_fd_sc_hd__o211a_1
X_17680_ _20464_/Q _17923_/A1 _17708_/S vssd1 vssd1 vccd1 vccd1 _20464_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14892_ _14894_/A _12469_/S _15026_/A _12463_/A _13635_/A vssd1 vssd1 vccd1 vccd1
+ _14893_/A sky130_fd_sc_hd__a32o_1
X_16631_ _19890_/Q _17945_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19890_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13843_ _20261_/Q _20260_/Q _13843_/C vssd1 vssd1 vccd1 vccd1 _13844_/B sky130_fd_sc_hd__and3_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19350_ _20710_/CLK _19350_/D vssd1 vssd1 vccd1 vccd1 _19350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16562_ _19847_/Q _16592_/A2 _16592_/B1 input17/X vssd1 vssd1 vccd1 vccd1 _16563_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10986_ _19401_/Q _10986_/B vssd1 vssd1 vccd1 vccd1 _10986_/X sky130_fd_sc_hd__or2_1
X_13774_ _13774_/A _13774_/B vssd1 vssd1 vccd1 vccd1 _13775_/B sky130_fd_sc_hd__nor2_8
XFILLER_262_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18301_ _20814_/Q _18300_/Y _18316_/S vssd1 vssd1 vccd1 vccd1 _18302_/B sky130_fd_sc_hd__mux2_1
X_15513_ input267/X _15013_/Y _15507_/X _15606_/A1 vssd1 vssd1 vccd1 vccd1 _15513_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19281_ _20315_/CLK _19281_/D vssd1 vssd1 vccd1 vccd1 _19281_/Q sky130_fd_sc_hd__dfxtp_1
X_12725_ _12726_/C _12726_/D vssd1 vssd1 vccd1 vccd1 _13377_/A sky130_fd_sc_hd__or2_1
X_16493_ _19800_/Q _17679_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19800_/D sky130_fd_sc_hd__mux2_1
XFILLER_231_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18232_ _18708_/A _18232_/B vssd1 vssd1 vccd1 vccd1 _20800_/D sky130_fd_sc_hd__and2_1
X_15444_ _19712_/Q _15475_/A2 _15475_/B1 _19744_/Q vssd1 vssd1 vccd1 vccd1 _15444_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12656_ _12680_/B _12656_/B vssd1 vssd1 vccd1 vccd1 _12656_/X sky130_fd_sc_hd__or2_1
XFILLER_169_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18163_ _18163_/A _18163_/B vssd1 vssd1 vccd1 vccd1 _18163_/Y sky130_fd_sc_hd__nand2_1
X_11607_ _12151_/A1 _11606_/X _11603_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _11607_/X
+ sky130_fd_sc_hd__o211a_1
X_12587_ _12587_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _12589_/C sky130_fd_sc_hd__nor2_1
X_15375_ _12468_/X _15374_/X _11401_/B vssd1 vssd1 vccd1 vccd1 _15378_/B sky130_fd_sc_hd__a21oi_1
XFILLER_184_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17114_ _20084_/Q _17114_/A1 _17114_/S vssd1 vssd1 vccd1 vccd1 _20084_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14326_ _14325_/A _14322_/B _14325_/X vssd1 vssd1 vccd1 vccd1 _14326_/X sky130_fd_sc_hd__a21bo_1
X_18094_ _18094_/A _18094_/B _18095_/B vssd1 vssd1 vccd1 vccd1 _20772_/D sky130_fd_sc_hd__nor3_1
X_11538_ _20166_/Q _11616_/B vssd1 vssd1 vccd1 vccd1 _11538_/X sky130_fd_sc_hd__or2_1
XFILLER_239_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17045_ input252/X _17015_/C _17015_/B vssd1 vssd1 vccd1 vccd1 _17045_/X sky130_fd_sc_hd__o21ba_1
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11469_ _12189_/A _11468_/X _11467_/X _11851_/C vssd1 vssd1 vccd1 vccd1 _11469_/X
+ sky130_fd_sc_hd__o211a_1
X_14257_ _20280_/Q _14267_/A2 _14267_/B1 input220/X vssd1 vssd1 vccd1 vccd1 _14259_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13208_ _13221_/B _13221_/C _13221_/A vssd1 vssd1 vccd1 vccd1 _13209_/C sky130_fd_sc_hd__o21ai_2
XFILLER_171_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14188_ _19501_/Q _14188_/B vssd1 vssd1 vccd1 vccd1 _14189_/B sky130_fd_sc_hd__nand2_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _13139_/A _19244_/Q vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__and2_1
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18996_ _18185_/Y _18983_/B _19002_/B1 _18995_/X vssd1 vssd1 vccd1 vccd1 _21017_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _20716_/Q _17947_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20716_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1470 _10630_/C1 vssd1 vssd1 vccd1 vccd1 _12082_/S sky130_fd_sc_hd__buf_4
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1481 _10629_/A vssd1 vssd1 vccd1 vccd1 _12023_/S sky130_fd_sc_hd__buf_6
X_17878_ _20651_/Q _17878_/A1 _17878_/S vssd1 vssd1 vccd1 vccd1 _20651_/D sky130_fd_sc_hd__mux2_1
Xfanout1492 _09728_/X vssd1 vssd1 vccd1 vccd1 _12342_/A sky130_fd_sc_hd__buf_12
XFILLER_226_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16829_ _16846_/A _09523_/Y _16809_/X _16828_/Y vssd1 vssd1 vccd1 vccd1 _16829_/X
+ sky130_fd_sc_hd__o211a_4
X_19617_ _19617_/CLK _19617_/D vssd1 vssd1 vccd1 vccd1 _19617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19548_ _20263_/CLK _19548_/D vssd1 vssd1 vccd1 vccd1 _19548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19479_ _20574_/CLK _19479_/D vssd1 vssd1 vccd1 vccd1 _19479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20323_ _20579_/CLK _20323_/D vssd1 vssd1 vccd1 vccd1 _20323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20254_ _20261_/CLK _20254_/D vssd1 vssd1 vccd1 vccd1 _20254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20185_ _20428_/CLK _20185_/D vssd1 vssd1 vccd1 vccd1 _20185_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09996_ _19885_/Q _19786_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _09996_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10840_ _19803_/Q _19307_/Q _12323_/S vssd1 vssd1 vccd1 vccd1 _10840_/X sky130_fd_sc_hd__mux2_1
XFILLER_272_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_260_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10771_ _10769_/X _10770_/X _12345_/S vssd1 vssd1 vccd1 vccd1 _10771_/X sky130_fd_sc_hd__mux2_1
XFILLER_241_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12510_ _12510_/A _14808_/A _12510_/C _15095_/B vssd1 vssd1 vccd1 vccd1 _12516_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_158_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13490_ _20948_/Q _09481_/Y _13564_/B _18570_/B vssd1 vssd1 vccd1 vccd1 _13490_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_200_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12441_ _12284_/A _12284_/B _13182_/A _12279_/Y _12282_/A vssd1 vssd1 vccd1 vccd1
+ _12442_/B sky130_fd_sc_hd__o32a_1
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12372_ _19428_/Q _20587_/Q _12375_/S vssd1 vssd1 vccd1 vccd1 _12372_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15160_ _15055_/X _15061_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _15161_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14111_ _16193_/A _14111_/B vssd1 vssd1 vccd1 vccd1 _14111_/Y sky130_fd_sc_hd__nand2_1
X_11323_ _11778_/B _11323_/B vssd1 vssd1 vccd1 vccd1 _11323_/Y sky130_fd_sc_hd__nand2_2
X_15091_ _19735_/Q _15453_/A2 _15080_/X _15019_/A _15090_/X vssd1 vssd1 vccd1 vccd1
+ _15091_/X sky130_fd_sc_hd__a221o_1
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14042_ _19213_/Q _14107_/C _14042_/S vssd1 vssd1 vccd1 vccd1 _14042_/X sky130_fd_sc_hd__mux2_1
X_11254_ _20461_/Q _20301_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _11254_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10205_ _09638_/Y _10202_/Y _10204_/X _10035_/Y vssd1 vssd1 vccd1 vccd1 _10205_/X
+ sky130_fd_sc_hd__o211a_1
X_18850_ _12967_/B _18864_/A2 _18864_/B1 _13426_/C vssd1 vssd1 vccd1 vccd1 _18851_/B
+ sky130_fd_sc_hd__a22o_1
X_11185_ _12569_/A _13644_/B _11184_/Y _11281_/B vssd1 vssd1 vccd1 vccd1 _11185_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_133_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17801_ _20578_/Q _17801_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20578_/D sky130_fd_sc_hd__mux2_1
XFILLER_268_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ _19878_/Q _19779_/Q _10137_/C vssd1 vssd1 vccd1 vccd1 _10136_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18781_ _20982_/Q _18819_/B vssd1 vssd1 vccd1 vccd1 _18781_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15993_ _21041_/Q _21009_/Q _15993_/S vssd1 vssd1 vccd1 vccd1 _15993_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ _20513_/Q _17906_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20513_/D sky130_fd_sc_hd__mux2_1
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14944_ _15133_/B _15012_/B vssd1 vssd1 vccd1 vccd1 _14980_/C sky130_fd_sc_hd__or2_2
X_10067_ _19279_/Q _09688_/B _11684_/A1 vssd1 vssd1 vccd1 vccd1 _10067_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17663_ _20449_/Q _17800_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20449_/D sky130_fd_sc_hd__mux2_1
XFILLER_48_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14875_ _14856_/X _14874_/X _15611_/S vssd1 vssd1 vccd1 vccd1 _14875_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19402_ _20561_/CLK _19402_/D vssd1 vssd1 vccd1 vccd1 _19402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16614_ _19873_/Q _17928_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19873_/D sky130_fd_sc_hd__mux2_1
X_13826_ _13826_/A1 _16239_/B _13826_/B1 _20624_/Q vssd1 vssd1 vccd1 vccd1 _13826_/X
+ sky130_fd_sc_hd__a22o_4
X_17594_ _20352_/Q _17871_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20352_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19333_ _20085_/CLK _19333_/D vssd1 vssd1 vccd1 vccd1 _19333_/Q sky130_fd_sc_hd__dfxtp_1
X_16545_ _16557_/A _16545_/B vssd1 vssd1 vccd1 vccd1 _19838_/D sky130_fd_sc_hd__or2_1
XFILLER_232_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ _13777_/A _13757_/B vssd1 vssd1 vccd1 vccd1 _13757_/X sky130_fd_sc_hd__or2_1
X_10969_ _15578_/S _10969_/B vssd1 vssd1 vccd1 vccd1 _15226_/A sky130_fd_sc_hd__nand2_2
XFILLER_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19264_ _20812_/CLK _19264_/D vssd1 vssd1 vccd1 vccd1 _19264_/Q sky130_fd_sc_hd__dfxtp_1
X_12708_ _12708_/A _12708_/B vssd1 vssd1 vccd1 vccd1 _12710_/B sky130_fd_sc_hd__or2_4
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16476_ _19785_/Q _17939_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19785_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13688_ _13688_/A _13698_/B vssd1 vssd1 vccd1 vccd1 _13688_/X sky130_fd_sc_hd__or2_4
X_18215_ _18499_/B vssd1 vssd1 vccd1 vccd1 _18215_/Y sky130_fd_sc_hd__inv_4
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15427_ _15283_/A _15413_/Y _16002_/B1 vssd1 vssd1 vccd1 vccd1 _15427_/X sky130_fd_sc_hd__a21o_1
X_19195_ _20665_/CLK _19195_/D vssd1 vssd1 vccd1 vccd1 _19195_/Q sky130_fd_sc_hd__dfxtp_1
X_12639_ _12639_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _12639_/X sky130_fd_sc_hd__or2_2
XFILLER_31_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18146_ _18148_/S _19111_/Q _14921_/X vssd1 vssd1 vccd1 vccd1 _18156_/C sky130_fd_sc_hd__a21o_1
XFILLER_102_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15358_ _15356_/A _15357_/X _15611_/S vssd1 vssd1 vccd1 vccd1 _15358_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14309_ _14301_/B _14304_/B _14301_/A vssd1 vssd1 vccd1 vccd1 _14314_/A sky130_fd_sc_hd__a21boi_1
X_18077_ _20766_/Q _20765_/Q _18077_/C vssd1 vssd1 vccd1 vccd1 _18079_/B sky130_fd_sc_hd__and3_1
XFILLER_172_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15289_ _15104_/X _15107_/X _15292_/S vssd1 vssd1 vccd1 vccd1 _15289_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17028_ _20006_/Q input192/X _17040_/S vssd1 vssd1 vccd1 vccd1 _20006_/D sky130_fd_sc_hd__mux2_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_236_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout707 _13802_/A1 vssd1 vssd1 vccd1 vccd1 _13826_/A1 sky130_fd_sc_hd__clkbuf_4
X_09850_ _12103_/A1 _09849_/X _09848_/X vssd1 vssd1 vccd1 vccd1 _09850_/X sky130_fd_sc_hd__o21a_1
Xfanout718 _13775_/A vssd1 vssd1 vccd1 vccd1 _13765_/A sky130_fd_sc_hd__buf_6
Xfanout729 _13142_/X vssd1 vssd1 vccd1 vccd1 _13478_/B sky130_fd_sc_hd__buf_8
XFILLER_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09781_ _09783_/A _11799_/B vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__or2_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _18560_/X _18978_/B _18977_/X _18978_/Y vssd1 vssd1 vccd1 vccd1 _18980_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20941_ _21011_/CLK _20941_/D vssd1 vssd1 vccd1 vccd1 _20941_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20872_ _21042_/CLK _20872_/D vssd1 vssd1 vccd1 vccd1 _20872_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20306_ _20630_/CLK _20306_/D vssd1 vssd1 vccd1 vccd1 _20306_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_49_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20180_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20237_ _21043_/CLK _20237_/D vssd1 vssd1 vccd1 vccd1 _20237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_276_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20168_ _20715_/CLK _20168_/D vssd1 vssd1 vccd1 vccd1 _20168_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09979_ _12140_/C1 _09978_/X _09975_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _09979_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20099_ _20718_/CLK _20099_/D vssd1 vssd1 vccd1 vccd1 _20099_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _19225_/Q _12990_/B _12990_/C vssd1 vssd1 vccd1 vccd1 _12991_/D sky130_fd_sc_hd__and3_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_268_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _11938_/X _11940_/X _11949_/S vssd1 vssd1 vccd1 vccd1 _11941_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_601 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_612 _12464_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_623 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _19422_/Q _17804_/A1 _14664_/S vssd1 vssd1 vccd1 vccd1 _19422_/D sky130_fd_sc_hd__mux2_1
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_634 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11872_/A _11872_/B _11871_/X vssd1 vssd1 vccd1 vccd1 _11872_/X sky130_fd_sc_hd__or3b_4
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_645 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13611_/A _13611_/B vssd1 vssd1 vccd1 vccd1 _15442_/B sky130_fd_sc_hd__xnor2_4
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ _20530_/Q _12323_/S vssd1 vssd1 vccd1 vccd1 _10823_/X sky130_fd_sc_hd__or2_1
X_14591_ _19357_/Q _17666_/A1 _14596_/S vssd1 vssd1 vccd1 vccd1 _19357_/D sky130_fd_sc_hd__mux2_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16330_ _19718_/Q _19719_/Q _16330_/C vssd1 vssd1 vccd1 vccd1 _16332_/B sky130_fd_sc_hd__and3_2
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13542_ _13612_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _13542_/X sky130_fd_sc_hd__and2_1
X_10754_ _19629_/Q _19935_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10754_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _19677_/Q _17692_/A1 _16277_/S vssd1 vssd1 vccd1 vccd1 _19677_/D sky130_fd_sc_hd__mux2_1
XFILLER_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ _19501_/Q _11189_/B vssd1 vssd1 vccd1 vccd1 _10685_/Y sky130_fd_sc_hd__nor2_1
X_13473_ split2/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13473_/X sky130_fd_sc_hd__and2b_2
XFILLER_186_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18000_ _20738_/Q _18003_/C _18094_/A vssd1 vssd1 vccd1 vccd1 _18000_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_145_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15212_ _15180_/X _15211_/X _15577_/S vssd1 vssd1 vccd1 vccd1 _15212_/X sky130_fd_sc_hd__mux2_4
X_12424_ _19692_/Q _20180_/Q _12428_/S vssd1 vssd1 vccd1 vccd1 _12424_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16192_ _19620_/Q _16000_/X _16196_/S vssd1 vssd1 vccd1 vccd1 _16193_/B sky130_fd_sc_hd__mux2_1
XFILLER_185_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15143_ input272/X _15482_/A2 _15142_/X vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__a21o_1
X_12355_ _20332_/Q _11213_/B _12354_/X vssd1 vssd1 vccd1 vccd1 _12355_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_154_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11306_ _20461_/Q _11295_/S _11304_/S vssd1 vssd1 vccd1 vccd1 _11306_/X sky130_fd_sc_hd__o21a_1
XFILLER_141_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15074_ _15468_/A _15066_/X _15072_/X _15073_/Y vssd1 vssd1 vccd1 vccd1 _15074_/X
+ sky130_fd_sc_hd__a211o_1
X_12286_ _12286_/A _13182_/A _12286_/C vssd1 vssd1 vccd1 vccd1 _15982_/B sky130_fd_sc_hd__and3_2
X_19951_ _20479_/CLK _19951_/D vssd1 vssd1 vccd1 vccd1 _19951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14025_ _12513_/B _14031_/A2 _14043_/B1 _14024_/X _16127_/B1 vssd1 vssd1 vccd1 vccd1
+ _19175_/D sky130_fd_sc_hd__o221a_1
X_11237_ _11246_/A1 _11235_/X _11236_/Y _11226_/X vssd1 vssd1 vccd1 vccd1 _11237_/X
+ sky130_fd_sc_hd__a31o_1
X_18902_ _18902_/A _18902_/B vssd1 vssd1 vccd1 vccd1 _18902_/Y sky130_fd_sc_hd__nand2_1
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19882_ _20574_/CLK _19882_/D vssd1 vssd1 vccd1 vccd1 _19882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11168_ _11359_/S _11166_/X _11167_/X vssd1 vssd1 vccd1 vccd1 _11168_/X sky130_fd_sc_hd__o21a_1
X_18833_ _20990_/Q _18861_/B vssd1 vssd1 vccd1 vccd1 _18833_/Y sky130_fd_sc_hd__nand2_1
XFILLER_268_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_256_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _10119_/A _10465_/A vssd1 vssd1 vccd1 vccd1 _10119_/Y sky130_fd_sc_hd__nand2_1
XFILLER_267_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18764_ _19084_/Q _12589_/B _12591_/X _13637_/A vssd1 vssd1 vccd1 vccd1 _18764_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ _19159_/Q _12569_/A vssd1 vssd1 vccd1 vccd1 _11099_/Y sky130_fd_sc_hd__nor2_1
X_15976_ _15526_/B _15959_/X _15975_/X _15976_/B2 vssd1 vssd1 vccd1 vccd1 _15976_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_95_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ _20496_/Q _17855_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20496_/D sky130_fd_sc_hd__mux2_1
X_14927_ _14927_/A _14960_/B vssd1 vssd1 vccd1 vccd1 _15019_/B sky130_fd_sc_hd__nor2_8
XFILLER_64_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18695_ _09480_/Y _18466_/B _18707_/S vssd1 vssd1 vccd1 vccd1 _18696_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17646_ _20432_/Q _17923_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20432_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14858_ _10802_/B _11958_/B _14870_/S vssd1 vssd1 vccd1 vccd1 _14858_/X sky130_fd_sc_hd__mux2_1
XFILLER_263_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13809_ _13816_/A1 _13715_/Y _13816_/B1 input224/X vssd1 vssd1 vccd1 vccd1 _13809_/X
+ sky130_fd_sc_hd__a22o_1
X_17577_ _20335_/Q _17888_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20335_/D sky130_fd_sc_hd__mux2_1
XFILLER_211_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ _19519_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14789_/X sky130_fd_sc_hd__or2_1
XFILLER_205_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19316_ _20315_/CLK _19316_/D vssd1 vssd1 vccd1 vccd1 _19316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16528_ _19864_/Q _16527_/Y _19863_/Q vssd1 vssd1 vccd1 vccd1 _16528_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_232_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19247_ _20621_/CLK _19247_/D vssd1 vssd1 vccd1 vccd1 _19247_/Q sky130_fd_sc_hd__dfxtp_1
X_16459_ _19768_/Q _17922_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19768_/D sky130_fd_sc_hd__mux2_1
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19178_ _19704_/CLK _19178_/D vssd1 vssd1 vccd1 vccd1 _19178_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_129_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18129_ _20785_/Q _18126_/B _18128_/Y vssd1 vssd1 vccd1 vccd1 _20785_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _12140_/C1 _09901_/X _09898_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _09902_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout504 _17779_/X vssd1 vssd1 vccd1 vccd1 _17808_/S sky130_fd_sc_hd__buf_12
Xfanout515 _17711_/X vssd1 vssd1 vccd1 vccd1 _17742_/S sky130_fd_sc_hd__buf_6
XFILLER_116_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout526 _17623_/S vssd1 vssd1 vccd1 vccd1 _17640_/S sky130_fd_sc_hd__buf_12
X_20022_ _20315_/CLK _20022_/D vssd1 vssd1 vccd1 vccd1 _20022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_263_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout537 _17215_/S vssd1 vssd1 vccd1 vccd1 _17217_/S sky130_fd_sc_hd__buf_12
X_09833_ _12102_/A1 _20515_/Q _10621_/S _20547_/Q vssd1 vssd1 vccd1 vccd1 _09833_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout548 _17083_/X vssd1 vssd1 vccd1 vccd1 _17112_/S sky130_fd_sc_hd__buf_12
XFILLER_113_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout559 _16673_/X vssd1 vssd1 vccd1 vccd1 _16704_/S sky130_fd_sc_hd__buf_6
XFILLER_259_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09764_ _11948_/A1 _09763_/X _09762_/X vssd1 vssd1 vccd1 vccd1 _09764_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_167_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20812_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09695_ _09695_/A _13192_/A vssd1 vssd1 vccd1 vccd1 _09695_/Y sky130_fd_sc_hd__nor2_8
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20924_ _20990_/CLK _20924_/D vssd1 vssd1 vccd1 vccd1 _20924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _21020_/CLK _20855_/D vssd1 vssd1 vccd1 vccd1 _20855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20786_ _20856_/CLK _20786_/D vssd1 vssd1 vccd1 vccd1 _20786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ _11236_/B _10470_/B vssd1 vssd1 vccd1 vccd1 _10470_/Y sky130_fd_sc_hd__nand2_1
XFILLER_167_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12140_ _12150_/S _12139_/X _12138_/X _12140_/C1 vssd1 vssd1 vccd1 vccd1 _12140_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_194_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12071_ _12069_/X _12070_/X _12071_/S vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _19801_/Q _11192_/A2 _11020_/X _11291_/B2 _11021_/X vssd1 vssd1 vccd1 vccd1
+ _11022_/X sky130_fd_sc_hd__o221a_1
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_249_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _20969_/Q _16045_/A2 _16016_/S _20841_/Q _15829_/X vssd1 vssd1 vccd1 vccd1
+ _15830_/X sky130_fd_sc_hd__a221o_1
XFILLER_49_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _19547_/Q _15980_/A2 _15760_/Y _16187_/A vssd1 vssd1 vccd1 vccd1 _19547_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_264_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12973_ _19103_/Q _19102_/Q _19101_/Q _19100_/Q vssd1 vssd1 vccd1 vccd1 _12974_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_252_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _20285_/Q _17502_/B vssd1 vssd1 vccd1 vccd1 _17500_/Y sky130_fd_sc_hd__nand2_1
X_14712_ _19469_/Q _17684_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19469_/D sky130_fd_sc_hd__mux2_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_261_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18480_ _18760_/B _18480_/B vssd1 vssd1 vccd1 vccd1 _18480_/X sky130_fd_sc_hd__or2_2
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _12003_/A _19922_/Q _11932_/S0 _20047_/Q vssd1 vssd1 vccd1 vccd1 _11924_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_233_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _20900_/Q _15937_/A2 _15994_/B1 _15691_/X _15937_/C1 vssd1 vssd1 vccd1 vccd1
+ _15692_/X sky130_fd_sc_hd__a221o_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_420 _09728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_431 _13777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _20260_/Q _20253_/Q _17433_/S vssd1 vssd1 vccd1 vccd1 _17432_/B sky130_fd_sc_hd__mux2_1
XANTENNA_442 _13725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _19405_/Q _17927_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19405_/D sky130_fd_sc_hd__mux2_1
XANTENNA_453 _19104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _11849_/X _11854_/X _12012_/S vssd1 vssd1 vccd1 vccd1 _11855_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_464 _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_475 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_486 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ _19532_/Q _09613_/A _18152_/C _19596_/Q vssd1 vssd1 vccd1 vccd1 _10806_/X
+ sky130_fd_sc_hd__a22o_1
X_17362_ _20229_/Q _17364_/A2 _17362_/B1 _20278_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17362_/X sky130_fd_sc_hd__a221o_1
XANTENNA_497 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14574_ _19340_/Q _17926_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19340_/D sky130_fd_sc_hd__mux2_1
XFILLER_198_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ _13636_/A _11786_/B _11786_/C _13637_/A vssd1 vssd1 vccd1 vccd1 _11786_/X
+ sky130_fd_sc_hd__and4_1
X_19101_ _19609_/CLK _19101_/D vssd1 vssd1 vccd1 vccd1 _19101_/Q sky130_fd_sc_hd__dfxtp_1
X_16313_ _19712_/Q _16314_/C _19713_/Q vssd1 vssd1 vccd1 vccd1 _16315_/B sky130_fd_sc_hd__a21oi_1
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13525_ _19661_/D _13522_/Y _13524_/Y _13624_/B2 vssd1 vssd1 vccd1 vccd1 _13525_/X
+ sky130_fd_sc_hd__a22o_4
X_17293_ _17293_/A _17329_/S _17305_/C vssd1 vssd1 vccd1 vccd1 _17293_/X sky130_fd_sc_hd__and3_1
X_10737_ _10735_/X _10736_/X _12376_/S vssd1 vssd1 vccd1 vccd1 _10737_/X sky130_fd_sc_hd__mux2_1
X_19032_ _18275_/Y _19046_/A2 _18760_/X _12553_/A _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19032_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16244_ _17850_/A _17184_/A vssd1 vssd1 vccd1 vccd1 _16245_/C sky130_fd_sc_hd__nor2_1
X_13456_ _13607_/B _13453_/X _13454_/Y _13455_/Y _18604_/B vssd1 vssd1 vccd1 vccd1
+ _13456_/X sky130_fd_sc_hd__o311a_2
X_10668_ _20404_/Q _12323_/S _10656_/X _12324_/S vssd1 vssd1 vccd1 vccd1 _10668_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ _19828_/Q _12412_/A2 _12405_/X _12412_/B2 _12406_/X vssd1 vssd1 vccd1 vccd1
+ _12407_/X sky130_fd_sc_hd__o221a_1
XFILLER_173_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16175_ _16187_/A _16175_/B vssd1 vssd1 vccd1 vccd1 _19611_/D sky130_fd_sc_hd__and2_1
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13387_ _14275_/A1 _19229_/Q _14772_/C1 _13386_/Y vssd1 vssd1 vccd1 vccd1 _13388_/D
+ sky130_fd_sc_hd__o211a_1
X_10599_ _10596_/X _10597_/X _10598_/Y vssd1 vssd1 vccd1 vccd1 _10642_/B sky130_fd_sc_hd__o21ai_4
XFILLER_154_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15126_ _11140_/B _12468_/X _15119_/Y _15125_/X vssd1 vssd1 vccd1 vccd1 _15126_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12338_ _19397_/Q _12412_/A2 _12336_/X _09738_/A _12337_/X vssd1 vssd1 vccd1 vccd1
+ _12338_/X sky130_fd_sc_hd__o221a_1
XFILLER_142_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19934_ _20085_/CLK _19934_/D vssd1 vssd1 vccd1 vccd1 _19934_/Q sky130_fd_sc_hd__dfxtp_1
X_15057_ _15053_/A _15056_/X _15254_/S vssd1 vssd1 vccd1 vccd1 _15057_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12269_ _12420_/B1 _12268_/X _12267_/X vssd1 vssd1 vccd1 vccd1 _12269_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_142_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_269_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14008_ _14029_/A1 _09672_/B _09943_/X _14041_/B1 _19851_/Q vssd1 vssd1 vccd1 vccd1
+ _14085_/C sky130_fd_sc_hd__o32a_1
X_19865_ _20704_/CLK _19865_/D vssd1 vssd1 vccd1 vccd1 _19865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18816_ _18830_/A _18816_/B vssd1 vssd1 vccd1 vccd1 _18816_/Y sky130_fd_sc_hd__nand2_1
X_19796_ _20719_/CLK _19796_/D vssd1 vssd1 vccd1 vccd1 _19796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18747_ _20974_/Q _18300_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18748_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15959_ _15219_/Y _15954_/Y _15955_/Y _15958_/X vssd1 vssd1 vccd1 vccd1 _15959_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_283_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09480_ _20948_/Q vssd1 vssd1 vccd1 vccd1 _09480_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18678_ _20943_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18678_/Y sky130_fd_sc_hd__nand2_1
XFILLER_224_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17629_ _20385_/Q _17800_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20385_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20640_ _20672_/CLK _20640_/D vssd1 vssd1 vccd1 vccd1 _20640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20571_ _20701_/CLK _20571_/D vssd1 vssd1 vccd1 vccd1 _20571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20005_ _20751_/CLK _20005_/D vssd1 vssd1 vccd1 vccd1 _20005_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09816_ _19645_/Q _12070_/S _09801_/X _12071_/S vssd1 vssd1 vccd1 vccd1 _09816_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_274_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09747_ _09747_/A _09747_/B _09747_/C _09632_/B vssd1 vssd1 vccd1 vccd1 _09750_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_274_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09678_ _09678_/A _09678_/B _09678_/C _09678_/D vssd1 vssd1 vccd1 vccd1 _09678_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_199_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _21009_/CLK _20907_/D vssd1 vssd1 vccd1 vccd1 _20907_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11640_ _12007_/A1 _19817_/Q _19321_/Q _11932_/S0 vssd1 vssd1 vccd1 vccd1 _11640_/X
+ sky130_fd_sc_hd__a22o_1
X_20838_ _21041_/CLK _20838_/D vssd1 vssd1 vccd1 vccd1 _20838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11571_ _19510_/Q _11570_/Y _11726_/S vssd1 vssd1 vccd1 vccd1 _11735_/B sky130_fd_sc_hd__mux2_4
X_20769_ _20796_/CLK _20769_/D vssd1 vssd1 vccd1 vccd1 _20769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_64_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20085_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13310_ _13281_/B _13309_/X _13107_/A vssd1 vssd1 vccd1 vccd1 _13310_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10522_ _10356_/A _20375_/Q _20439_/Q _11295_/S vssd1 vssd1 vccd1 vccd1 _10522_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14290_ _19511_/Q _14294_/B vssd1 vssd1 vccd1 vccd1 _14302_/A sky130_fd_sc_hd__and2_1
XFILLER_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13241_ _13230_/X _13240_/X _14794_/C1 vssd1 vssd1 vccd1 vccd1 _13242_/D sky130_fd_sc_hd__o21a_1
XFILLER_108_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10453_ _10453_/A vssd1 vssd1 vccd1 vccd1 _10456_/A sky130_fd_sc_hd__inv_2
XFILLER_182_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10384_ _10035_/Y _10378_/X _10383_/X _10373_/X _10024_/X vssd1 vssd1 vccd1 vccd1
+ _10385_/B sky130_fd_sc_hd__a32o_2
XFILLER_163_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13172_ _11880_/B _13434_/B _11878_/B vssd1 vssd1 vccd1 vccd1 _13433_/B sky130_fd_sc_hd__o21bai_4
XFILLER_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12123_ _12138_/A1 _19362_/Q _20717_/Q _12124_/S _12123_/C1 vssd1 vssd1 vccd1 vccd1
+ _12123_/X sky130_fd_sc_hd__a221o_1
XFILLER_272_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17980_ _18080_/A _17985_/C vssd1 vssd1 vccd1 vccd1 _17980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16931_ _17006_/A1 _15807_/X _16879_/X _16930_/X vssd1 vssd1 vccd1 vccd1 _16931_/X
+ sky130_fd_sc_hd__o211a_1
Xfanout1800 _16769_/S vssd1 vssd1 vccd1 vccd1 _16846_/A sky130_fd_sc_hd__clkbuf_8
X_12054_ _12052_/X _12053_/X _12056_/S vssd1 vssd1 vccd1 vccd1 _12054_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1811 _19527_/Q vssd1 vssd1 vccd1 vccd1 _09659_/B sky130_fd_sc_hd__buf_8
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1822 _19175_/Q vssd1 vssd1 vccd1 vccd1 _12513_/B sky130_fd_sc_hd__buf_12
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1833 _19172_/Q vssd1 vssd1 vccd1 vccd1 _12136_/B1 sky130_fd_sc_hd__buf_6
Xfanout1844 _12584_/C vssd1 vssd1 vccd1 vccd1 _11336_/A sky130_fd_sc_hd__clkbuf_8
X_11005_ _19932_/Q _11008_/A3 _11169_/B _11250_/S vssd1 vssd1 vccd1 vccd1 _11005_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_237_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16862_ _19229_/Q _16862_/A2 _17005_/A2 _19098_/Q _16861_/X vssd1 vssd1 vccd1 vccd1
+ _16862_/X sky130_fd_sc_hd__o221a_1
Xfanout1855 _18765_/B vssd1 vssd1 vccd1 vccd1 _12828_/A sky130_fd_sc_hd__clkbuf_16
X_19650_ _19956_/CLK _19650_/D vssd1 vssd1 vccd1 vccd1 _19650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_266_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1866 _15678_/A1 vssd1 vssd1 vccd1 vccd1 _12504_/A sky130_fd_sc_hd__buf_12
XFILLER_277_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1877 _19166_/Q vssd1 vssd1 vccd1 vccd1 _09731_/A sky130_fd_sc_hd__buf_6
XFILLER_226_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout890 _18563_/X vssd1 vssd1 vccd1 vccd1 _18621_/A2 sky130_fd_sc_hd__buf_6
X_18601_ _18493_/X _18621_/A2 _18599_/Y _18600_/Y vssd1 vssd1 vccd1 vccd1 _18602_/B
+ sky130_fd_sc_hd__o211a_1
Xfanout1888 _14802_/C1 vssd1 vssd1 vccd1 vccd1 _16191_/A sky130_fd_sc_hd__buf_4
X_15813_ _19172_/Q _15978_/A2 _13414_/Y _15895_/S vssd1 vssd1 vccd1 vccd1 _15814_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_19581_ _19589_/CLK _19581_/D vssd1 vssd1 vccd1 vccd1 _19581_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1899 fanout1905/X vssd1 vssd1 vccd1 vccd1 _14794_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_253_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16793_ _19967_/Q _16849_/A _16792_/Y _16451_/A vssd1 vssd1 vccd1 vccd1 _19967_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_219_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18532_ _18651_/B _18532_/B vssd1 vssd1 vccd1 vccd1 _18532_/X sky130_fd_sc_hd__or2_2
XFILLER_218_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15744_ _20742_/Q _15934_/A2 _15934_/B1 _20774_/Q vssd1 vssd1 vccd1 vccd1 _15744_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12956_ _16945_/C _17219_/A vssd1 vssd1 vccd1 vccd1 _18136_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _18490_/A _18463_/B vssd1 vssd1 vccd1 vccd1 _18463_/X sky130_fd_sc_hd__or2_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _20650_/Q _20614_/Q _11915_/S vssd1 vssd1 vccd1 vccd1 _11907_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15675_ _15890_/B _15658_/X _15674_/X _15544_/A vssd1 vssd1 vccd1 vccd1 _15675_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ _12917_/A _12887_/B vssd1 vssd1 vccd1 vccd1 _13233_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_261 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_272 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17414_ _17402_/Y _17413_/X _17412_/X _17434_/A vssd1 vssd1 vccd1 vccd1 _20253_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _19390_/Q _17910_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19390_/D sky130_fd_sc_hd__mux2_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _18414_/A _18394_/B vssd1 vssd1 vccd1 vccd1 _20851_/D sky130_fd_sc_hd__and2_1
XANTENNA_283 _20624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ _11836_/X _11837_/X _12150_/S vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_294 input224/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17345_ _20221_/Q _17363_/A2 _17344_/X _18700_/A vssd1 vssd1 vccd1 vccd1 _20221_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _19327_/Q _17911_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19327_/D sky130_fd_sc_hd__mux2_1
XFILLER_202_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11769_ _11319_/A _13523_/A _11779_/B _11323_/Y vssd1 vssd1 vccd1 vccd1 _11775_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13508_ _12584_/A _19218_/Q _13507_/X vssd1 vssd1 vccd1 vccd1 _13909_/A sky130_fd_sc_hd__a21oi_4
X_17276_ _20197_/Q _17330_/A2 _17279_/C1 _17275_/X vssd1 vssd1 vccd1 vccd1 _17276_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14488_ _17851_/A _17676_/B _14488_/C vssd1 vssd1 vccd1 vccd1 _14488_/X sky130_fd_sc_hd__and3_4
XFILLER_228_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_0__f_wb_clk_i clkbuf_3_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_4_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
X_19015_ _21027_/Q _19015_/B vssd1 vssd1 vccd1 vccd1 _19015_/X sky130_fd_sc_hd__or2_1
X_16227_ _19650_/Q _17111_/A1 _16227_/S vssd1 vssd1 vccd1 vccd1 _19650_/D sky130_fd_sc_hd__mux2_1
XFILLER_162_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13439_ _15949_/B _15898_/A _13439_/C vssd1 vssd1 vccd1 vccd1 _13440_/A sky130_fd_sc_hd__or3_1
XFILLER_127_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16158_ _16842_/B _16178_/S vssd1 vssd1 vccd1 vccd1 _16158_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15109_ _15105_/X _15108_/X _15577_/S vssd1 vssd1 vccd1 vccd1 _15109_/X sky130_fd_sc_hd__mux2_2
XFILLER_115_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16089_ _19569_/Q _16081_/B _16143_/A vssd1 vssd1 vccd1 vccd1 _16089_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19917_ _20677_/CLK _19917_/D vssd1 vssd1 vccd1 vccd1 _19917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_256_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19848_ _20014_/CLK _19848_/D vssd1 vssd1 vccd1 vccd1 _19848_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09601_ _09609_/A _19094_/Q vssd1 vssd1 vccd1 vccd1 _17538_/C sky130_fd_sc_hd__nand2b_4
XFILLER_84_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19779_ _20570_/CLK _19779_/D vssd1 vssd1 vccd1 vccd1 _19779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_260_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09532_ _19526_/Q _19149_/Q vssd1 vssd1 vccd1 vccd1 _09532_/X sky130_fd_sc_hd__and2b_1
XFILLER_25_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20623_ _20624_/CLK _20623_/D vssd1 vssd1 vccd1 vccd1 _20623_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20554_ _20686_/CLK _20554_/D vssd1 vssd1 vccd1 vccd1 _20554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20485_ _21046_/A _20485_/D vssd1 vssd1 vccd1 vccd1 _20485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_285_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput460 _19513_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[19] sky130_fd_sc_hd__buf_4
Xoutput471 _19523_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[29] sky130_fd_sc_hd__buf_4
Xoutput482 output482/A vssd1 vssd1 vccd1 vccd1 probe_state sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_182_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20421_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xfanout1107 _11964_/X vssd1 vssd1 vccd1 vccd1 _17913_/A1 sky130_fd_sc_hd__buf_4
Xfanout1118 _17904_/A1 vssd1 vssd1 vccd1 vccd1 _17870_/A1 sky130_fd_sc_hd__buf_4
XFILLER_114_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1129 _17592_/A1 vssd1 vssd1 vccd1 vccd1 _17903_/A1 sky130_fd_sc_hd__buf_4
XFILLER_219_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_111_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20862_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_21037_ _21041_/CLK _21037_/D vssd1 vssd1 vccd1 vccd1 _21037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12810_ _19513_/Q _12835_/A _19514_/Q vssd1 vssd1 vccd1 vccd1 _12811_/B sky130_fd_sc_hd__a21oi_1
XFILLER_90_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_274_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13790_ _13790_/A split1/A vssd1 vssd1 vccd1 vccd1 _13790_/X sky130_fd_sc_hd__and2_4
XFILLER_263_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12741_/A vssd1 vssd1 vccd1 vccd1 _12741_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _12578_/B _12762_/Y _15459_/X _15589_/S vssd1 vssd1 vccd1 vccd1 _15460_/X
+ sky130_fd_sc_hd__o211a_1
X_12672_ _12674_/B _12674_/C _12674_/A vssd1 vssd1 vccd1 vccd1 _12675_/A sky130_fd_sc_hd__a21o_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _20295_/Q _14431_/A2 _14431_/B1 input236/X vssd1 vssd1 vccd1 vccd1 _14413_/B
+ sky130_fd_sc_hd__a22o_4
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11641_/S _11620_/X _11622_/X vssd1 vssd1 vccd1 vccd1 _11623_/X sky130_fd_sc_hd__a21o_1
X_15391_ _20794_/Q _15016_/Y _15334_/B _15142_/S vssd1 vssd1 vccd1 vccd1 _15391_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17130_ _20098_/Q _17689_/A1 _17132_/S vssd1 vssd1 vccd1 vccd1 _20098_/D sky130_fd_sc_hd__mux2_1
X_14342_ _19516_/Q _14342_/B vssd1 vssd1 vccd1 vccd1 _14343_/C sky130_fd_sc_hd__xnor2_1
XFILLER_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11554_ _19414_/Q _09931_/S _11553_/X _09986_/C vssd1 vssd1 vccd1 vccd1 _11554_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10505_ _09689_/A _10488_/X _10504_/X _11012_/A vssd1 vssd1 vccd1 vccd1 _13675_/C
+ sky130_fd_sc_hd__a211o_4
X_17061_ _20033_/Q _17095_/A1 _17076_/S vssd1 vssd1 vccd1 vccd1 _20033_/D sky130_fd_sc_hd__mux2_1
XFILLER_7_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14273_ _14273_/A _14278_/B vssd1 vssd1 vccd1 vccd1 _14273_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ _12189_/A _11485_/B vssd1 vssd1 vccd1 vccd1 _11485_/X sky130_fd_sc_hd__or2_1
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _19764_/Q _14948_/Y _16011_/X _16049_/A1 _16048_/C1 vssd1 vssd1 vccd1 vccd1
+ _16012_/X sky130_fd_sc_hd__a221o_1
X_13224_ _13323_/C _12996_/Y _13222_/X _13223_/X vssd1 vssd1 vccd1 vccd1 _13224_/X
+ sky130_fd_sc_hd__a31o_1
X_10436_ _10581_/A1 _20504_/Q _12064_/S _20536_/Q vssd1 vssd1 vccd1 vccd1 _10436_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13155_ _13155_/A _13155_/B vssd1 vssd1 vccd1 vccd1 _13459_/B sky130_fd_sc_hd__nand2_2
X_10367_ _13423_/A vssd1 vssd1 vccd1 vccd1 _10367_/Y sky130_fd_sc_hd__inv_2
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12106_ _09728_/X _12088_/X _12105_/X vssd1 vssd1 vccd1 vccd1 _12106_/X sky130_fd_sc_hd__o21a_2
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17963_ _20725_/Q _17961_/A _17963_/B1 vssd1 vssd1 vccd1 vccd1 _17964_/B sky130_fd_sc_hd__o21ai_1
X_10298_ _19879_/Q _19780_/Q _10303_/S vssd1 vssd1 vccd1 vccd1 _10298_/X sky130_fd_sc_hd__mux2_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _13086_/A _13086_/B _13086_/C vssd1 vssd1 vccd1 vccd1 _13227_/A sky130_fd_sc_hd__nor3_2
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19702_ _19704_/CLK _19702_/D vssd1 vssd1 vccd1 vccd1 _19702_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1630 _09617_/Y vssd1 vssd1 vccd1 vccd1 fanout1630/X sky130_fd_sc_hd__buf_12
X_12037_ _13431_/A vssd1 vssd1 vccd1 vccd1 _12288_/A sky130_fd_sc_hd__inv_2
X_16914_ _19235_/Q _16980_/A2 _16980_/B1 _19104_/Q _16913_/X vssd1 vssd1 vccd1 vccd1
+ _16914_/X sky130_fd_sc_hd__o221a_1
XFILLER_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1641 _12922_/X vssd1 vssd1 vccd1 vccd1 _17502_/B sky130_fd_sc_hd__clkbuf_8
X_17894_ _20665_/Q _17894_/A1 _17916_/S vssd1 vssd1 vccd1 vccd1 _20665_/D sky130_fd_sc_hd__mux2_1
Xfanout1652 _09670_/Y vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__buf_2
Xfanout1663 _11261_/C vssd1 vssd1 vccd1 vccd1 _10979_/C sky130_fd_sc_hd__buf_12
Xfanout1674 _09672_/A vssd1 vssd1 vccd1 vccd1 _11228_/A1 sky130_fd_sc_hd__buf_6
X_19633_ _20667_/CLK _19633_/D vssd1 vssd1 vccd1 vccd1 _19633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1685 _12711_/A vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__buf_4
XFILLER_238_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16845_ _16805_/X _16842_/Y _16844_/X _16932_/A1 vssd1 vssd1 vccd1 vccd1 _16845_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_254_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1696 _12254_/A vssd1 vssd1 vccd1 vccd1 _12347_/A1 sky130_fd_sc_hd__buf_4
XFILLER_225_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19564_ _19574_/CLK _19564_/D vssd1 vssd1 vccd1 vccd1 _19564_/Q sky130_fd_sc_hd__dfxtp_1
X_16776_ _19089_/Q _16996_/B1 _16775_/X vssd1 vssd1 vccd1 vccd1 _16776_/X sky130_fd_sc_hd__o21a_1
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13988_ _19195_/Q _14071_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _13988_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15727_ _16051_/A1 _15713_/Y _16051_/B1 vssd1 vssd1 vccd1 vccd1 _15727_/Y sky130_fd_sc_hd__o21ai_1
X_18515_ _20898_/Q _18559_/B _18514_/X _18458_/B vssd1 vssd1 vccd1 vccd1 _18516_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12939_ _19257_/Q _12964_/A2 _16945_/B _20005_/Q vssd1 vssd1 vccd1 vccd1 _12944_/C
+ sky130_fd_sc_hd__a22o_2
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _21004_/CLK _19495_/D vssd1 vssd1 vccd1 vccd1 _19495_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_280_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18446_ _18754_/A _18446_/B vssd1 vssd1 vccd1 vccd1 _20877_/D sky130_fd_sc_hd__and2_1
X_15658_ _15652_/X _15653_/X _15657_/X vssd1 vssd1 vccd1 vccd1 _15658_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14609_ _19373_/Q _17893_/A1 _14632_/S vssd1 vssd1 vccd1 vccd1 _19373_/D sky130_fd_sc_hd__mux2_1
XFILLER_222_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18377_ _18544_/B _18387_/B vssd1 vssd1 vccd1 vccd1 _18377_/Y sky130_fd_sc_hd__nand2_1
XFILLER_194_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15589_ _13426_/B _15588_/X _15589_/S vssd1 vssd1 vccd1 vccd1 _15589_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17328_ _20215_/Q _17328_/A2 _17327_/X _17974_/B1 vssd1 vssd1 vccd1 vccd1 _20215_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17259_ _20192_/Q _17268_/A2 _17257_/X _17258_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1
+ _20192_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20270_ _21013_/CLK _20270_/D vssd1 vssd1 vccd1 vccd1 _20270_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09515_ _17998_/A vssd1 vssd1 vccd1 vccd1 _09515_/Y sky130_fd_sc_hd__clkinv_8
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_262_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20606_ _20685_/CLK _20606_/D vssd1 vssd1 vccd1 vccd1 _20606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20537_ _20669_/CLK _20537_/D vssd1 vssd1 vccd1 vccd1 _20537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20468_ _20468_/CLK _20468_/D vssd1 vssd1 vccd1 vccd1 _20468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ _19929_/Q _11270_/A2 _09688_/B _11250_/S vssd1 vssd1 vccd1 vccd1 _11270_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10221_ _10219_/X _10220_/X _12377_/S vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20399_ _20428_/CLK _20399_/D vssd1 vssd1 vccd1 vccd1 _20399_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_106_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10152_ _10150_/X _10151_/X _10152_/S vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput290 _13832_/X vssd1 vssd1 vccd1 vccd1 addr0[5] sky130_fd_sc_hd__buf_4
X_14960_ _14927_/A _14960_/B vssd1 vssd1 vccd1 vccd1 _15014_/D sky130_fd_sc_hd__and2b_1
X_10083_ _09829_/A _20377_/Q _20441_/Q _10400_/S _11304_/S vssd1 vssd1 vccd1 vccd1
+ _10083_/X sky130_fd_sc_hd__a221o_1
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13911_ _13911_/A _13919_/S vssd1 vssd1 vccd1 vccd1 _13911_/Y sky130_fd_sc_hd__nand2_1
XFILLER_275_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_275_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14891_ _13694_/A _12466_/Y _14815_/S _16053_/B _14878_/Y vssd1 vssd1 vccd1 vccd1
+ _14891_/X sky130_fd_sc_hd__o221a_1
XFILLER_247_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16630_ _19889_/Q _17804_/A1 _16634_/S vssd1 vssd1 vccd1 vccd1 _19889_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13842_ _20259_/Q _20258_/Q _20257_/Q vssd1 vssd1 vccd1 vccd1 _13843_/C sky130_fd_sc_hd__and3_1
XFILLER_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_262_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16561_ _16593_/A _16561_/B vssd1 vssd1 vccd1 vccd1 _19846_/D sky130_fd_sc_hd__or2_1
XFILLER_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13773_ _13693_/X _13741_/B _13741_/Y _13694_/X _13772_/X vssd1 vssd1 vccd1 vccd1
+ _13774_/B sky130_fd_sc_hd__o221a_4
X_10985_ _09618_/A _10983_/X _10984_/X _11345_/S vssd1 vssd1 vccd1 vccd1 _10985_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15512_ _20862_/Q _15511_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15512_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18300_ _18550_/B vssd1 vssd1 vccd1 vccd1 _18300_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19280_ _20694_/CLK _19280_/D vssd1 vssd1 vccd1 vccd1 _19280_/Q sky130_fd_sc_hd__dfxtp_1
X_12724_ _12709_/X _12716_/Y _12721_/Y _12722_/X vssd1 vssd1 vccd1 vccd1 _12726_/D
+ sky130_fd_sc_hd__a211oi_2
X_16492_ _19799_/Q _17051_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19799_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18231_ _20800_/Q _18230_/Y _18311_/S vssd1 vssd1 vccd1 vccd1 _18232_/B sky130_fd_sc_hd__mux2_1
XFILLER_95_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15443_ _15443_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _15443_/Y sky130_fd_sc_hd__nand2_1
X_12655_ _19497_/Q _12665_/A vssd1 vssd1 vccd1 vccd1 _12656_/B sky130_fd_sc_hd__nor2_1
X_18162_ _18418_/A _18162_/B vssd1 vssd1 vccd1 vccd1 _20786_/D sky130_fd_sc_hd__and2_1
X_11606_ _11604_/X _11605_/X _11917_/S vssd1 vssd1 vccd1 vccd1 _11606_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15374_ _12471_/X _12466_/Y _15374_/S vssd1 vssd1 vccd1 vccd1 _15374_/X sky130_fd_sc_hd__mux2_1
X_12586_ _13193_/B vssd1 vssd1 vccd1 vccd1 _12592_/A sky130_fd_sc_hd__inv_2
XFILLER_157_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17113_ _20083_/Q _17915_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20083_/D sky130_fd_sc_hd__mux2_1
X_14325_ _14325_/A _14325_/B _14333_/B vssd1 vssd1 vccd1 vccd1 _14325_/X sky130_fd_sc_hd__or3b_1
X_18093_ _20772_/Q _20771_/Q _18093_/C vssd1 vssd1 vccd1 vccd1 _18095_/B sky130_fd_sc_hd__and3_4
X_11537_ _11537_/A1 _15922_/B2 _11536_/X vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__a21oi_2
XFILLER_117_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17044_ _18985_/A _17044_/B _17044_/C vssd1 vssd1 vccd1 vccd1 _20020_/D sky130_fd_sc_hd__and3_1
X_14256_ _19228_/Q _14256_/A2 _14255_/X _18352_/C1 vssd1 vssd1 vccd1 vccd1 _19228_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11468_ _19284_/Q _20071_/Q _12182_/S vssd1 vssd1 vccd1 vccd1 _11468_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13207_ _12871_/A _12871_/B _12896_/A vssd1 vssd1 vccd1 vccd1 _13221_/C sky130_fd_sc_hd__a21oi_1
X_10419_ _20129_/Q _20097_/Q _10428_/S vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__mux2_1
X_14187_ _19501_/Q _14188_/B vssd1 vssd1 vccd1 vccd1 _14189_/A sky130_fd_sc_hd__or2_2
XFILLER_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11399_ _11400_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _15374_/S sky130_fd_sc_hd__and2_2
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _18767_/A _13137_/X _13133_/Y _13373_/A vssd1 vssd1 vccd1 vccd1 _13138_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _21017_/Q _18997_/B vssd1 vssd1 vccd1 vccd1 _18995_/X sky130_fd_sc_hd__or2_1
XFILLER_135_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13069_ _13043_/Y _13605_/A _13604_/B vssd1 vssd1 vccd1 vccd1 _13453_/C sky130_fd_sc_hd__o21ai_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _20715_/Q _17946_/A1 _17946_/S vssd1 vssd1 vccd1 vccd1 _20715_/D sky130_fd_sc_hd__mux2_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1460 _09733_/Y vssd1 vssd1 vccd1 vccd1 _12012_/S sky130_fd_sc_hd__buf_8
Xfanout1471 _11204_/S vssd1 vssd1 vccd1 vccd1 _10630_/C1 sky130_fd_sc_hd__buf_4
XFILLER_239_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17877_ _20650_/Q _17877_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20650_/D sky130_fd_sc_hd__mux2_1
Xfanout1482 _12426_/S vssd1 vssd1 vccd1 vccd1 _10629_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_253_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1493 _11895_/B vssd1 vssd1 vccd1 vccd1 _11897_/B sky130_fd_sc_hd__buf_8
XFILLER_54_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19616_ _20649_/CLK _19616_/D vssd1 vssd1 vccd1 vccd1 _19616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_285_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16828_ _16846_/A input79/X vssd1 vssd1 vccd1 vccd1 _16828_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19547_ _20263_/CLK _19547_/D vssd1 vssd1 vccd1 vccd1 _19547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16759_ input76/X input71/X _16799_/S vssd1 vssd1 vccd1 vccd1 _16760_/A sky130_fd_sc_hd__mux2_2
XFILLER_206_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19478_ _20677_/CLK _19478_/D vssd1 vssd1 vccd1 vccd1 _19478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18429_ _20869_/Q _18255_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18430_/B sky130_fd_sc_hd__mux2_1
XFILLER_210_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20322_ _20482_/CLK _20322_/D vssd1 vssd1 vccd1 vccd1 _20322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20253_ _20261_/CLK _20253_/D vssd1 vssd1 vccd1 vccd1 _20253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_282_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20184_ _20184_/CLK _20184_/D vssd1 vssd1 vccd1 vccd1 _20184_/Q sky130_fd_sc_hd__dfxtp_1
X_09995_ _09989_/X _09994_/X _12012_/S vssd1 vssd1 vccd1 vccd1 _09995_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10770_ _19629_/Q _19935_/Q _19273_/Q _20060_/Q _11116_/S _12406_/C vssd1 vssd1 vccd1
+ vccd1 _10770_/X sky130_fd_sc_hd__mux4_1
XFILLER_198_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ _12440_/A _14882_/A vssd1 vssd1 vccd1 vccd1 _12447_/B sky130_fd_sc_hd__and2_2
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _12371_/A1 _19364_/Q _20719_/Q _12375_/S _12371_/C1 vssd1 vssd1 vccd1 vccd1
+ _12371_/X sky130_fd_sc_hd__a221o_1
XFILLER_197_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14110_ _14110_/A _14110_/B _14110_/C vssd1 vssd1 vccd1 vccd1 _14111_/B sky130_fd_sc_hd__or3_2
XFILLER_153_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11322_ _10884_/A _11322_/B vssd1 vssd1 vccd1 vccd1 _11323_/B sky130_fd_sc_hd__nand2b_1
XFILLER_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15090_ _17242_/A _15089_/X _15452_/S vssd1 vssd1 vccd1 vccd1 _15090_/X sky130_fd_sc_hd__mux2_2
XFILLER_181_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14041_ _14041_/A1 _14041_/A2 _09647_/X _14041_/B1 _19862_/Q vssd1 vssd1 vccd1 vccd1
+ _14107_/C sky130_fd_sc_hd__o32a_1
X_11253_ _11259_/S _11251_/X _11252_/X vssd1 vssd1 vccd1 vccd1 _11253_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10204_ _10037_/Y _10203_/Y _09669_/X vssd1 vssd1 vccd1 vccd1 _10204_/X sky130_fd_sc_hd__a21o_1
X_11184_ _19158_/Q _12569_/A vssd1 vssd1 vccd1 vccd1 _11184_/Y sky130_fd_sc_hd__nor2_1
XFILLER_267_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17800_ _20577_/Q _17800_/A1 _17808_/S vssd1 vssd1 vccd1 vccd1 _20577_/D sky130_fd_sc_hd__mux2_1
X_10135_ _10133_/X _10134_/X _10235_/S vssd1 vssd1 vccd1 vccd1 _10135_/X sky130_fd_sc_hd__mux2_1
X_18780_ _18574_/Y _18867_/A2 _18779_/Y _18901_/S vssd1 vssd1 vccd1 vccd1 _18780_/X
+ sky130_fd_sc_hd__a22o_1
X_15992_ _20879_/Q _16042_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15992_/X sky130_fd_sc_hd__o21ba_1
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_283_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14943_ _15133_/B _15012_/B vssd1 vssd1 vccd1 vccd1 _15308_/B sky130_fd_sc_hd__nor2_2
XFILLER_236_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10066_ _11281_/A _20066_/Q _11268_/C vssd1 vssd1 vccd1 vccd1 _10066_/X sky130_fd_sc_hd__and3_1
X_17731_ _20512_/Q _17871_/A1 _17740_/S vssd1 vssd1 vccd1 vccd1 _20512_/D sky130_fd_sc_hd__mux2_1
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17662_ _20448_/Q _17696_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20448_/D sky130_fd_sc_hd__mux2_1
X_14874_ _14865_/X _14873_/X _15357_/S vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19401_ _20692_/CLK _19401_/D vssd1 vssd1 vccd1 vccd1 _19401_/Q sky130_fd_sc_hd__dfxtp_1
X_16613_ _19872_/Q _17684_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19872_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13825_ _13826_/A1 _16237_/B _13826_/B1 _20623_/Q vssd1 vssd1 vccd1 vccd1 _13825_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_211_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17593_ _20351_/Q _17904_/A1 _17601_/S vssd1 vssd1 vccd1 vccd1 _20351_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19332_ _20084_/CLK _19332_/D vssd1 vssd1 vccd1 vccd1 _19332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16544_ _19838_/Q _16578_/A2 _16578_/B1 input39/X vssd1 vssd1 vccd1 vccd1 _16545_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13756_ _11999_/Y _13742_/B _13663_/A vssd1 vssd1 vccd1 vccd1 _13759_/A sky130_fd_sc_hd__o21a_2
X_10968_ _15578_/S _10969_/B vssd1 vssd1 vccd1 vccd1 _10968_/Y sky130_fd_sc_hd__nor2_1
X_12707_ _19509_/Q _12758_/B vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__and2_1
X_19263_ _20990_/CLK _19263_/D vssd1 vssd1 vccd1 vccd1 _19263_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16475_ _19784_/Q _17938_/A1 _16483_/S vssd1 vssd1 vccd1 vccd1 _19784_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13687_ _13765_/A _13687_/B vssd1 vssd1 vccd1 vccd1 _13687_/X sky130_fd_sc_hd__and2_1
X_10899_ _11008_/A1 _20497_/Q _10986_/B _20529_/Q vssd1 vssd1 vccd1 vccd1 _10899_/X
+ sky130_fd_sc_hd__o22a_1
X_18214_ _18213_/B _14229_/B _18213_/Y vssd1 vssd1 vccd1 vccd1 _18499_/B sky130_fd_sc_hd__o21ai_4
XFILLER_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15426_ _15644_/A1 _16815_/B _15413_/Y vssd1 vssd1 vccd1 vccd1 _15426_/Y sky130_fd_sc_hd__o21ai_1
X_19194_ _20670_/CLK _19194_/D vssd1 vssd1 vccd1 vccd1 _19194_/Q sky130_fd_sc_hd__dfxtp_1
X_12638_ _19500_/Q _12647_/A vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__nor2_1
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18145_ _18148_/S _19109_/Q _14915_/X vssd1 vssd1 vccd1 vccd1 _18156_/B sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_214_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20573_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15357_ _15166_/Y _15172_/B _15357_/S vssd1 vssd1 vccd1 vccd1 _15357_/X sky130_fd_sc_hd__mux2_1
X_12569_ _12569_/A _12587_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _12589_/A sky130_fd_sc_hd__nor3_1
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14308_ _19233_/Q _14398_/A2 _14307_/X _14776_/C1 vssd1 vssd1 vccd1 vccd1 _19233_/D
+ sky130_fd_sc_hd__o211a_1
X_18076_ _20765_/Q _18077_/C _20766_/Q vssd1 vssd1 vccd1 vccd1 _18078_/B sky130_fd_sc_hd__a21oi_1
XFILLER_102_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15288_ _19532_/Q _15402_/A _15287_/Y _15288_/C1 vssd1 vssd1 vccd1 vccd1 _19532_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17027_ _20005_/Q input191/X _17040_/S vssd1 vssd1 vccd1 vccd1 _20005_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14239_ _19506_/Q _14239_/B vssd1 vssd1 vccd1 vccd1 _14240_/C sky130_fd_sc_hd__xnor2_1
XFILLER_113_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout708 _13810_/A1 vssd1 vssd1 vccd1 vccd1 _13802_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout719 _13624_/B2 vssd1 vssd1 vccd1 vccd1 _13626_/B2 sky130_fd_sc_hd__buf_4
XFILLER_213_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09780_ _19517_/Q _15822_/A _15895_/S vssd1 vssd1 vccd1 vccd1 _11799_/B sky130_fd_sc_hd__mux2_8
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18978_ _21011_/Q _18978_/B vssd1 vssd1 vccd1 vccd1 _18978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _20698_/Q _17929_/A1 _17946_/S vssd1 vssd1 vccd1 vccd1 _20698_/D sky130_fd_sc_hd__mux2_1
XFILLER_252_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1290 _09541_/Y vssd1 vssd1 vccd1 vccd1 _12832_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_282_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20940_ _21011_/CLK _20940_/D vssd1 vssd1 vccd1 vccd1 _20940_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20871_ _21042_/CLK _20871_/D vssd1 vssd1 vccd1 vccd1 _20871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20305_ _20465_/CLK _20305_/D vssd1 vssd1 vccd1 vccd1 _20305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20236_ _21043_/CLK _20236_/D vssd1 vssd1 vccd1 vccd1 _20236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19574_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20167_ _20641_/CLK _20167_/D vssd1 vssd1 vccd1 vccd1 _20167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_276_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09978_ _09976_/X _09977_/X _11528_/S vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__mux2_1
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20479_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_276_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20098_ _20711_/CLK _20098_/D vssd1 vssd1 vccd1 vccd1 _20098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _20326_/Q _11947_/S _11939_/X vssd1 vssd1 vccd1 vccd1 _11940_/X sky130_fd_sc_hd__a21o_1
XFILLER_268_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_602 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_613 _12464_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ _11949_/S _11866_/Y _11868_/Y _11870_/Y _12020_/C1 vssd1 vssd1 vccd1 vccd1
+ _11871_/X sky130_fd_sc_hd__a221o_1
XFILLER_72_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_624 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_635 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_646 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ _14244_/A1 _19225_/Q _14758_/C1 _13609_/Y vssd1 vssd1 vccd1 vccd1 _13610_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _20338_/Q _12295_/B vssd1 vssd1 vccd1 vccd1 _10822_/X sky130_fd_sc_hd__or2_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _19356_/Q _17942_/A1 _14594_/S vssd1 vssd1 vccd1 vccd1 _19356_/D sky130_fd_sc_hd__mux2_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13541_ _13541_/A _13541_/B vssd1 vssd1 vccd1 vccd1 _15303_/B sky130_fd_sc_hd__xnor2_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10753_ _12399_/A1 _10752_/X _10749_/X _12392_/C1 vssd1 vssd1 vccd1 vccd1 _10753_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_213_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16260_ _19676_/Q _17657_/A1 _16275_/S vssd1 vssd1 vccd1 vccd1 _19676_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13472_ _13472_/A vssd1 vssd1 vccd1 vccd1 _13472_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _11368_/A1 _13661_/B _10683_/X _11189_/B vssd1 vssd1 vccd1 vccd1 _10718_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_40_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _14832_/X _14824_/X _15215_/S vssd1 vssd1 vccd1 vccd1 _15211_/X sky130_fd_sc_hd__mux2_1
X_12423_ _11118_/A _12418_/Y _12422_/Y _12431_/A1 vssd1 vssd1 vccd1 vccd1 _12423_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_185_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16191_ _16191_/A _16191_/B vssd1 vssd1 vccd1 vccd1 _19619_/D sky130_fd_sc_hd__and2_1
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15142_ _15133_/X _15141_/X _15142_/S vssd1 vssd1 vccd1 vccd1 _15142_/X sky130_fd_sc_hd__mux2_1
X_12354_ _20492_/Q _12352_/S _11212_/S vssd1 vssd1 vccd1 vccd1 _12354_/X sky130_fd_sc_hd__o21a_1
XFILLER_193_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11305_ _20301_/Q _11305_/B vssd1 vssd1 vccd1 vccd1 _11305_/X sky130_fd_sc_hd__or2_1
XFILLER_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15073_ _14882_/B _16025_/B _15220_/A vssd1 vssd1 vccd1 vccd1 _15073_/Y sky130_fd_sc_hd__o21ai_1
X_19950_ _20075_/CLK _19950_/D vssd1 vssd1 vccd1 vccd1 _19950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12285_ _12286_/A _12286_/C _13182_/A vssd1 vssd1 vccd1 vccd1 _15982_/A sky130_fd_sc_hd__a21oi_2
XFILLER_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ _19207_/Q _14095_/C _14042_/S vssd1 vssd1 vccd1 vccd1 _14024_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18901_ _19514_/Q _18900_/X _18901_/S vssd1 vssd1 vccd1 vccd1 _18902_/B sky130_fd_sc_hd__mux2_1
X_11236_ _11236_/A _11236_/B _11236_/C vssd1 vssd1 vccd1 vccd1 _11236_/Y sky130_fd_sc_hd__nand3_1
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_268_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19881_ _20673_/CLK _19881_/D vssd1 vssd1 vccd1 vccd1 _19881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18832_ _18604_/Y _18867_/A2 _18830_/Y _18831_/Y vssd1 vssd1 vccd1 vccd1 _18832_/X
+ sky130_fd_sc_hd__a22o_1
X_11167_ _12371_/A1 _20366_/Q _20430_/Q _12296_/S _12301_/S vssd1 vssd1 vccd1 vccd1
+ _11167_/X sky130_fd_sc_hd__a221o_1
XFILLER_95_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xsplit1 split1/A vssd1 vssd1 vccd1 vccd1 split1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_268_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10118_ _10373_/A _11234_/B _10117_/X vssd1 vssd1 vccd1 vccd1 _10118_/X sky130_fd_sc_hd__or3b_2
X_18763_ _18763_/A1 _12982_/C _18762_/X _18476_/A vssd1 vssd1 vccd1 vccd1 _20979_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11098_ _12245_/A1 _17782_/A1 _11097_/X vssd1 vssd1 vccd1 vccd1 _13646_/B sky130_fd_sc_hd__o21ai_4
X_15975_ _16024_/A1 _15973_/X _15974_/Y _15954_/A _15975_/B2 vssd1 vssd1 vccd1 vccd1
+ _15975_/X sky130_fd_sc_hd__a32o_1
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ _20495_/Q _17888_/A1 _17742_/S vssd1 vssd1 vccd1 vccd1 _20495_/D sky130_fd_sc_hd__mux2_1
X_14926_ _12959_/B _12584_/B _18148_/S vssd1 vssd1 vccd1 vccd1 _14960_/B sky130_fd_sc_hd__mux2_4
X_10049_ _19410_/Q _20569_/Q _10485_/S vssd1 vssd1 vccd1 vccd1 _10049_/X sky130_fd_sc_hd__mux2_1
X_18694_ _18694_/A _18694_/B vssd1 vssd1 vccd1 vccd1 _20947_/D sky130_fd_sc_hd__and2_1
XFILLER_270_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17645_ _20431_/Q _17922_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20431_/D sky130_fd_sc_hd__mux2_1
XFILLER_223_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14857_ _10803_/B _12115_/B _14870_/S vssd1 vssd1 vccd1 vccd1 _14857_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13808_ _13816_/A1 _13711_/B _13816_/B1 input223/X vssd1 vssd1 vccd1 vccd1 _13808_/X
+ sky130_fd_sc_hd__a22o_1
X_17576_ _20334_/Q _17887_/A1 _17606_/S vssd1 vssd1 vccd1 vccd1 _20334_/D sky130_fd_sc_hd__mux2_1
X_14788_ _19141_/Q _14802_/A2 _14787_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _19518_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19315_ _20633_/CLK _19315_/D vssd1 vssd1 vccd1 vccd1 _19315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16527_ input9/X _16594_/B vssd1 vssd1 vccd1 vccd1 _16527_/Y sky130_fd_sc_hd__nand2_1
X_13739_ _11842_/Y _13742_/B _13663_/A vssd1 vssd1 vccd1 vccd1 _13744_/A sky130_fd_sc_hd__o21a_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19246_ _19246_/CLK _19246_/D vssd1 vssd1 vccd1 vccd1 _19246_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_220_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16458_ _19767_/Q _17921_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19767_/D sky130_fd_sc_hd__mux2_1
XFILLER_176_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15409_ _15468_/A _15409_/B vssd1 vssd1 vccd1 vccd1 _15409_/Y sky130_fd_sc_hd__nand2_1
X_16389_ _18064_/A _16394_/C vssd1 vssd1 vccd1 vccd1 _16389_/Y sky130_fd_sc_hd__nor2_1
X_19177_ _20665_/CLK _19177_/D vssd1 vssd1 vccd1 vccd1 _19177_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_145_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18128_ _20785_/Q _18126_/B _18126_/A vssd1 vssd1 vccd1 vccd1 _18128_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_247_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18059_ _20759_/Q _18061_/C _18058_/Y vssd1 vssd1 vccd1 vccd1 _20759_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _09899_/X _09900_/X _09901_/S vssd1 vssd1 vccd1 vccd1 _09901_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout505 _17779_/X vssd1 vssd1 vccd1 vccd1 _17806_/S sky130_fd_sc_hd__clkbuf_8
X_20021_ _20621_/CLK _20021_/D vssd1 vssd1 vccd1 vccd1 _20021_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_141_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout516 _17676_/X vssd1 vssd1 vccd1 vccd1 _17705_/S sky130_fd_sc_hd__clkbuf_16
Xfanout527 _17608_/X vssd1 vssd1 vccd1 vccd1 _17623_/S sky130_fd_sc_hd__buf_12
XFILLER_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09832_ _09830_/X _09831_/X _12082_/S vssd1 vssd1 vccd1 vccd1 _09832_/X sky130_fd_sc_hd__mux2_1
Xfanout538 _17212_/S vssd1 vssd1 vccd1 vccd1 _17215_/S sky130_fd_sc_hd__buf_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout549 _17083_/X vssd1 vssd1 vccd1 vccd1 _17111_/S sky130_fd_sc_hd__buf_6
XFILLER_140_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09763_ _19888_/Q _19789_/Q _11936_/S vssd1 vssd1 vccd1 vccd1 _09763_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09694_ _19421_/Q _11599_/S _09693_/X _12123_/C1 vssd1 vssd1 vccd1 vccd1 _09694_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_227_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_273_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20923_ _21023_/CLK _20923_/D vssd1 vssd1 vccd1 vccd1 _20923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20854_ _20863_/CLK _20854_/D vssd1 vssd1 vccd1 vccd1 _20854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20785_ _21020_/CLK _20785_/D vssd1 vssd1 vccd1 vccd1 _20785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_259_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12070_ _19293_/Q _20080_/Q _12070_/S vssd1 vssd1 vccd1 vccd1 _12070_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11021_ _11021_/A _19305_/Q _11021_/C vssd1 vssd1 vccd1 vccd1 _11021_/X sky130_fd_sc_hd__or3_1
XFILLER_150_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20219_ _20268_/CLK _20219_/D vssd1 vssd1 vccd1 vccd1 _20219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _15814_/A _15760_/B _15760_/C vssd1 vssd1 vccd1 vccd1 _15760_/Y sky130_fd_sc_hd__nand3_1
X_12972_ _19114_/Q _12972_/B _12972_/C _12972_/D vssd1 vssd1 vccd1 vccd1 _12975_/C
+ sky130_fd_sc_hd__or4_2
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14711_ _19468_/Q _17683_/A1 _14736_/S vssd1 vssd1 vccd1 vccd1 _19468_/D sky130_fd_sc_hd__mux2_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11923_ _12513_/B _11649_/S _11922_/Y vssd1 vssd1 vccd1 vccd1 _11955_/A sky130_fd_sc_hd__o21a_2
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_273_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15691_ _21030_/Q _20998_/Q _15993_/S vssd1 vssd1 vccd1 vccd1 _15691_/X sky130_fd_sc_hd__mux2_1
XANTENNA_410 _18205_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_421 _09889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _19404_/Q _17926_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19404_/D sky130_fd_sc_hd__mux2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17430_ _17430_/A _17430_/B vssd1 vssd1 vccd1 vccd1 _20259_/D sky130_fd_sc_hd__or2_1
XANTENNA_432 _13666_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11854_ _11852_/X _11853_/X _12011_/S vssd1 vssd1 vccd1 vccd1 _11854_/X sky130_fd_sc_hd__mux2_1
XANTENNA_443 _13725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_454 _19104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_465 _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_476 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10805_ _13567_/A _13541_/A _10804_/Y vssd1 vssd1 vccd1 vccd1 _10805_/Y sky130_fd_sc_hd__o21bai_2
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14573_ _19339_/Q _17925_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19339_/D sky130_fd_sc_hd__mux2_1
X_17361_ _20229_/Q _17363_/A2 _17360_/X _18700_/A vssd1 vssd1 vccd1 vccd1 _20229_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_487 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_498 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ _13694_/A _14878_/A vssd1 vssd1 vccd1 vccd1 _11785_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19100_ _19609_/CLK _19100_/D vssd1 vssd1 vccd1 vccd1 _19100_/Q sky130_fd_sc_hd__dfxtp_1
X_16312_ _19712_/Q _16314_/C _16311_/Y vssd1 vssd1 vccd1 vccd1 _19712_/D sky130_fd_sc_hd__o21a_1
X_13524_ _13524_/A vssd1 vssd1 vccd1 vccd1 _13524_/Y sky130_fd_sc_hd__inv_2
X_17292_ _20203_/Q _17331_/A2 _17290_/X _17291_/X _17331_/C1 vssd1 vssd1 vccd1 vccd1
+ _20203_/D sky130_fd_sc_hd__o221a_1
X_10736_ _20124_/Q _20092_/Q _11074_/S vssd1 vssd1 vccd1 vccd1 _10736_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16243_ _19095_/Q _16243_/B _17538_/C vssd1 vssd1 vccd1 vccd1 _17184_/A sky130_fd_sc_hd__or3_2
XFILLER_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19031_ _21034_/Q _19049_/A2 _19030_/X _18734_/A vssd1 vssd1 vccd1 vccd1 _21034_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13455_ _20957_/Q _13607_/B vssd1 vssd1 vccd1 vccd1 _13455_/Y sky130_fd_sc_hd__nand2_1
X_10667_ _11094_/S _10666_/X _10665_/X _12398_/C1 vssd1 vssd1 vccd1 vccd1 _10667_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12406_ _12411_/A _19332_/Q _12406_/C vssd1 vssd1 vccd1 vccd1 _12406_/X sky130_fd_sc_hd__or3_1
X_16174_ _19611_/Q _15753_/X _16190_/S vssd1 vssd1 vccd1 vccd1 _16175_/B sky130_fd_sc_hd__mux2_1
XFILLER_63_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13386_ _13381_/X _13385_/Y _14275_/A1 vssd1 vssd1 vccd1 vccd1 _13386_/Y sky130_fd_sc_hd__o21ai_1
X_10598_ _12517_/C _12577_/A _12581_/A vssd1 vssd1 vccd1 vccd1 _10598_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_126_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15125_ _13482_/A _12471_/X _14837_/S _15123_/X _15124_/Y vssd1 vssd1 vccd1 vccd1
+ _15125_/X sky130_fd_sc_hd__o221a_1
X_12337_ _12337_/A _20688_/Q _12337_/C vssd1 vssd1 vccd1 vccd1 _12337_/X sky130_fd_sc_hd__or3_1
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19933_ _20690_/CLK _19933_/D vssd1 vssd1 vccd1 vccd1 _19933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15056_ _15054_/X _15055_/X _15155_/S vssd1 vssd1 vccd1 vccd1 _15056_/X sky130_fd_sc_hd__mux2_1
X_12268_ _19894_/Q _19795_/Q _12268_/S vssd1 vssd1 vccd1 vccd1 _12268_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14007_ _10866_/A _14031_/A2 _14040_/B1 _14006_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1
+ _19169_/D sky130_fd_sc_hd__o221a_1
XFILLER_269_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11219_ _12433_/A1 _17921_/A1 _11218_/Y _09750_/Y vssd1 vssd1 vccd1 vccd1 _11219_/X
+ sky130_fd_sc_hd__o2bb2a_4
X_19864_ _20812_/CLK _19864_/D vssd1 vssd1 vccd1 vccd1 _19864_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12199_ _12197_/Y _12199_/B vssd1 vssd1 vccd1 vccd1 _12200_/A sky130_fd_sc_hd__nand2b_2
XFILLER_228_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18815_ _19092_/Q _12589_/B _12592_/C _15369_/A vssd1 vssd1 vccd1 vccd1 _18816_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19795_ _20179_/CLK _19795_/D vssd1 vssd1 vccd1 vccd1 _19795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18746_ _18746_/A _18746_/B vssd1 vssd1 vccd1 vccd1 _20973_/D sky130_fd_sc_hd__and2_1
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15958_ _12200_/A _16054_/B _15956_/X _15957_/X vssd1 vssd1 vccd1 vccd1 _15958_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_255_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput190 localMemory_wb_adr_i[0] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14909_ _14973_/A vssd1 vssd1 vccd1 vccd1 _14958_/A sky130_fd_sc_hd__inv_2
XFILLER_224_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_252_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18677_ _18960_/A _18677_/B vssd1 vssd1 vccd1 vccd1 _20942_/D sky130_fd_sc_hd__nor2_1
XFILLER_36_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15889_ _14870_/S _15294_/X _15297_/Y _15468_/A _15888_/X vssd1 vssd1 vccd1 vccd1
+ _15890_/C sky130_fd_sc_hd__a221o_4
XFILLER_263_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17628_ _20384_/Q _17696_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20384_/D sky130_fd_sc_hd__mux2_1
XFILLER_197_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17559_ _20319_/Q _17870_/A1 _17567_/S vssd1 vssd1 vccd1 vccd1 _20319_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20570_ _20570_/CLK _20570_/D vssd1 vssd1 vccd1 vccd1 _20570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19229_ _19695_/CLK _19229_/D vssd1 vssd1 vccd1 vccd1 _19229_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_177_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_279_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20004_ _20004_/CLK _20004_/D vssd1 vssd1 vccd1 vccd1 _20004_/Q sky130_fd_sc_hd__dfxtp_4
X_09815_ _10585_/S _09814_/X _09813_/X _11680_/C1 vssd1 vssd1 vccd1 vccd1 _09815_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09746_ _09746_/A _09746_/B _09746_/C _09743_/X vssd1 vssd1 vccd1 vccd1 _09747_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09676_/A _09676_/B _09669_/X vssd1 vssd1 vccd1 vccd1 _09678_/D sky130_fd_sc_hd__a21oi_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20906_ _21010_/CLK _20906_/D vssd1 vssd1 vccd1 vccd1 _20906_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ _21043_/CLK _20837_/D vssd1 vssd1 vccd1 vccd1 _20837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11570_ _15630_/A vssd1 vssd1 vccd1 vccd1 _11570_/Y sky130_fd_sc_hd__inv_2
X_20768_ _20796_/CLK _20768_/D vssd1 vssd1 vccd1 vccd1 _20768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ _20471_/Q _11295_/S _11304_/S vssd1 vssd1 vccd1 vccd1 _10521_/X sky130_fd_sc_hd__o21a_1
XFILLER_210_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20699_ _20701_/CLK _20699_/D vssd1 vssd1 vccd1 vccd1 _20699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13240_ _13139_/A _19240_/Q _13239_/X vssd1 vssd1 vccd1 vccd1 _13240_/X sky130_fd_sc_hd__a21o_2
X_10452_ _10640_/B _10455_/B vssd1 vssd1 vccd1 vccd1 _10453_/A sky130_fd_sc_hd__nor2_1
XFILLER_183_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ _09782_/A _13413_/B _09784_/B vssd1 vssd1 vccd1 vccd1 _13434_/B sky130_fd_sc_hd__a21oi_4
X_10383_ _10037_/Y _10382_/Y _09669_/X vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__a21o_1
XFILLER_272_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20379_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12122_ _12125_/A1 _12121_/X _12120_/X vssd1 vssd1 vccd1 vccd1 _12122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12053_ _20144_/Q _20112_/Q _12053_/S vssd1 vssd1 vccd1 vccd1 _12053_/X sky130_fd_sc_hd__mux2_1
X_16930_ _19237_/Q _17003_/B _16964_/B1 _19106_/Q _16929_/X vssd1 vssd1 vccd1 vccd1
+ _16930_/X sky130_fd_sc_hd__o221a_2
Xfanout1801 _16769_/S vssd1 vssd1 vccd1 vccd1 _16884_/S sky130_fd_sc_hd__buf_4
XFILLER_78_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1812 _09666_/B vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__buf_4
Xfanout1823 _12135_/A vssd1 vssd1 vccd1 vccd1 _11904_/S sky130_fd_sc_hd__buf_6
Xfanout1834 _11101_/A vssd1 vssd1 vccd1 vccd1 _09502_/A sky130_fd_sc_hd__buf_8
X_11004_ _19270_/Q _09688_/B _11009_/B2 vssd1 vssd1 vccd1 vccd1 _11004_/X sky130_fd_sc_hd__a21o_1
XFILLER_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1845 _12584_/C vssd1 vssd1 vccd1 vccd1 _09503_/A sky130_fd_sc_hd__buf_8
X_16861_ _20411_/Q _17004_/A2 _17004_/B1 vssd1 vssd1 vccd1 vccd1 _16861_/X sky130_fd_sc_hd__a21o_1
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1856 _18765_/B vssd1 vssd1 vccd1 vccd1 _12514_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_78_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1867 _19167_/Q vssd1 vssd1 vccd1 vccd1 _15678_/A1 sky130_fd_sc_hd__buf_12
XFILLER_237_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout880 _15395_/S vssd1 vssd1 vccd1 vccd1 _15454_/S sky130_fd_sc_hd__buf_6
Xfanout1878 _12510_/A vssd1 vssd1 vccd1 vccd1 _14895_/A sky130_fd_sc_hd__buf_8
X_18600_ _19503_/Q _18604_/B vssd1 vssd1 vccd1 vccd1 _18600_/Y sky130_fd_sc_hd__nand2_1
Xfanout891 _18563_/X vssd1 vssd1 vccd1 vccd1 _18564_/A sky130_fd_sc_hd__clkbuf_4
Xfanout1889 _13887_/C1 vssd1 vssd1 vccd1 vccd1 _14802_/C1 sky130_fd_sc_hd__clkbuf_4
X_15812_ _15948_/A1 _12804_/Y _15811_/X _12832_/B vssd1 vssd1 vccd1 vccd1 _15814_/B
+ sky130_fd_sc_hd__a22o_1
X_19580_ _20665_/CLK _19580_/D vssd1 vssd1 vccd1 vccd1 _19580_/Q sky130_fd_sc_hd__dfxtp_1
X_16792_ _16788_/Y _16791_/X _17011_/B1 vssd1 vssd1 vccd1 vccd1 _16792_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_65_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_265_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18531_ _18932_/A _18531_/B vssd1 vssd1 vccd1 vccd1 _20903_/D sky130_fd_sc_hd__nor2_1
XFILLER_234_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12955_ _17461_/A _12930_/B _13790_/A _14237_/A2 vssd1 vssd1 vccd1 vccd1 _17219_/A
+ sky130_fd_sc_hd__a31o_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15743_ _19722_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15743_/X sky130_fd_sc_hd__or2_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11906_ _11983_/A1 _20518_/Q _11513_/S _11896_/X vssd1 vssd1 vccd1 vccd1 _11906_/X
+ sky130_fd_sc_hd__o211a_1
X_18462_ _18462_/A _18462_/B _12592_/B vssd1 vssd1 vccd1 vccd1 _18462_/X sky130_fd_sc_hd__or3b_2
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _19519_/Q _12916_/A2 _12885_/X _12916_/B2 vssd1 vssd1 vccd1 vccd1 _12887_/B
+ sky130_fd_sc_hd__o22a_2
X_15674_ _16052_/A1 _15672_/X _15673_/Y _13427_/B _16052_/B2 vssd1 vssd1 vccd1 vccd1
+ _15674_/X sky130_fd_sc_hd__a32o_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_251 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_262 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17413_ _20260_/Q _20252_/Q _17442_/A vssd1 vssd1 vccd1 vccd1 _17413_/X sky130_fd_sc_hd__mux2_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_273 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ _19291_/Q _20078_/Q _11987_/S vssd1 vssd1 vccd1 vccd1 _11837_/X sky130_fd_sc_hd__mux2_1
X_14625_ _19389_/Q _17909_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19389_/D sky130_fd_sc_hd__mux2_1
X_18393_ _20851_/Q _18165_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18394_/B sky130_fd_sc_hd__mux2_1
XFILLER_221_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_284 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 input225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17344_ _20220_/Q _17364_/A2 _17370_/B1 _20269_/Q _17370_/C1 vssd1 vssd1 vccd1 vccd1
+ _17344_/X sky130_fd_sc_hd__a221o_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14556_ _19326_/Q _17910_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19326_/D sky130_fd_sc_hd__mux2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11768_ _11754_/B _11768_/B vssd1 vssd1 vccd1 vccd1 _11768_/X sky130_fd_sc_hd__and2b_1
XFILLER_186_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13507_ _13552_/A _13507_/B _13507_/C vssd1 vssd1 vccd1 vccd1 _13507_/X sky130_fd_sc_hd__and3_2
X_10719_ _10720_/B vssd1 vssd1 vccd1 vccd1 _10719_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17275_ _17275_/A _17275_/B _17290_/C vssd1 vssd1 vccd1 vccd1 _17275_/X sky130_fd_sc_hd__and3_1
X_14487_ _17850_/A _17082_/A vssd1 vssd1 vccd1 vccd1 _14488_/C sky130_fd_sc_hd__nor2_1
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11699_ _09834_/C _11698_/X _12091_/S vssd1 vssd1 vccd1 vccd1 _11699_/X sky130_fd_sc_hd__a21o_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19014_ _18230_/Y _18982_/B _19016_/B1 _19013_/X vssd1 vssd1 vccd1 vccd1 _21026_/D
+ sky130_fd_sc_hd__o211a_1
X_13438_ _13245_/A _13245_/B _16242_/B vssd1 vssd1 vccd1 vccd1 _13438_/Y sky130_fd_sc_hd__a21oi_4
X_16226_ _19649_/Q _17178_/A1 _16227_/S vssd1 vssd1 vccd1 vccd1 _19649_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16157_ _19602_/Q _16164_/B _16156_/Y _16143_/A vssd1 vssd1 vccd1 vccd1 _19602_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_142_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13369_ _13368_/A _13368_/B _13370_/B vssd1 vssd1 vccd1 vccd1 _13369_/X sky130_fd_sc_hd__a21o_1
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15108_ _15107_/X _15106_/X _15292_/S vssd1 vssd1 vccd1 vccd1 _15108_/X sky130_fd_sc_hd__mux2_1
X_16088_ _10546_/X _16106_/A2 _16087_/X vssd1 vssd1 vccd1 vccd1 _19568_/D sky130_fd_sc_hd__o21a_1
XFILLER_142_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15039_ _15039_/A _15039_/B vssd1 vssd1 vccd1 vccd1 _15039_/Y sky130_fd_sc_hd__nor2_1
X_19916_ _20480_/CLK _19916_/D vssd1 vssd1 vccd1 vccd1 _19916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19847_ _20014_/CLK _19847_/D vssd1 vssd1 vccd1 vccd1 _19847_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_284_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09600_ _09609_/A _19095_/Q vssd1 vssd1 vccd1 vccd1 _14668_/B sky130_fd_sc_hd__nand2b_4
XFILLER_272_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19778_ _20451_/CLK _19778_/D vssd1 vssd1 vccd1 vccd1 _19778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_216_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09531_ _19864_/Q _19863_/Q vssd1 vssd1 vccd1 vccd1 _09531_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18729_ _20965_/Q _18255_/Y _18749_/S vssd1 vssd1 vccd1 vccd1 _18730_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_280_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20622_ _20624_/CLK _20622_/D vssd1 vssd1 vccd1 vccd1 _20622_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_177_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20553_ _20685_/CLK _20553_/D vssd1 vssd1 vccd1 vccd1 _20553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20484_ _20580_/CLK _20484_/D vssd1 vssd1 vccd1 vccd1 _20484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_285_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput450 _19494_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[0] sky130_fd_sc_hd__buf_4
Xoutput461 _19495_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[1] sky130_fd_sc_hd__buf_4
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput472 _19496_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[2] sky130_fd_sc_hd__buf_4
XFILLER_78_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput483 _13469_/Y vssd1 vssd1 vccd1 vccd1 web0 sky130_fd_sc_hd__buf_4
Xfanout1108 _17911_/A1 vssd1 vssd1 vccd1 vccd1 _17945_/A1 sky130_fd_sc_hd__buf_4
XFILLER_133_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1119 _11689_/X vssd1 vssd1 vccd1 vccd1 _17904_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_87_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21036_ _21042_/CLK _21036_/D vssd1 vssd1 vccd1 vccd1 _21036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09729_ _19168_/Q _13863_/A vssd1 vssd1 vccd1 vccd1 _09729_/Y sky130_fd_sc_hd__nand2_8
XFILLER_216_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_151_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20959_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12740_ _19507_/Q _12740_/B vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__xnor2_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ _12674_/B _12674_/C _12674_/A vssd1 vssd1 vccd1 vccd1 _12676_/A sky130_fd_sc_hd__a21oi_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _19243_/Q _14438_/A2 _14409_/X _14794_/C1 vssd1 vssd1 vccd1 vccd1 _19243_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11622_ _12003_/C _11621_/X _11933_/S vssd1 vssd1 vccd1 vccd1 _11622_/X sky130_fd_sc_hd__a21o_1
X_15390_ _15140_/S _15383_/X _15389_/X _15384_/Y vssd1 vssd1 vccd1 vccd1 _15390_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ _19516_/Q _14342_/B vssd1 vssd1 vccd1 vccd1 _14354_/A sky130_fd_sc_hd__nand2_1
X_11553_ _20573_/Q _11616_/B vssd1 vssd1 vccd1 vccd1 _11553_/X sky130_fd_sc_hd__or2_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10504_ _09689_/C _10492_/X _10495_/X _10503_/X vssd1 vssd1 vccd1 vccd1 _10504_/X
+ sky130_fd_sc_hd__o31a_1
X_17060_ _20032_/Q _17060_/A1 _17081_/S vssd1 vssd1 vccd1 vccd1 _20032_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14272_ _14271_/A _14271_/B _14271_/C vssd1 vssd1 vccd1 vccd1 _14278_/B sky130_fd_sc_hd__a21oi_2
X_11484_ _20478_/Q _20318_/Q _12188_/S vssd1 vssd1 vccd1 vccd1 _11485_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16011_ _20752_/Q _16011_/A2 _16011_/B1 _20784_/Q vssd1 vssd1 vccd1 vccd1 _16011_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13223_ _20940_/Q _13366_/C1 _18667_/B vssd1 vssd1 vccd1 vccd1 _13223_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10435_ _20408_/Q _10502_/A2 _10432_/X _10433_/X _10434_/X vssd1 vssd1 vccd1 vccd1
+ _10435_/X sky130_fd_sc_hd__o221a_1
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ _13596_/A _13596_/B _10540_/X _15410_/S vssd1 vssd1 vccd1 vccd1 _13155_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10366_ _10366_/A _15580_/S vssd1 vssd1 vccd1 vccd1 _13423_/A sky130_fd_sc_hd__nand2_8
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12105_/A _12105_/B _12104_/X vssd1 vssd1 vccd1 vccd1 _12105_/X sky130_fd_sc_hd__or3b_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _20725_/Q _20724_/Q _17962_/C vssd1 vssd1 vccd1 vccd1 _17965_/B sky130_fd_sc_hd__and3_2
X_13085_ _13015_/X _13084_/Y _13016_/Y vssd1 vssd1 vccd1 vccd1 _13086_/C sky130_fd_sc_hd__a21boi_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10297_ _10295_/X _10296_/X _11256_/S vssd1 vssd1 vccd1 vccd1 _10297_/X sky130_fd_sc_hd__mux2_1
X_19701_ _19701_/CLK _19701_/D vssd1 vssd1 vccd1 vccd1 _19701_/Q sky130_fd_sc_hd__dfxtp_4
Xfanout1620 _10322_/S vssd1 vssd1 vccd1 vccd1 _11256_/S sky130_fd_sc_hd__buf_8
X_16913_ _20417_/Q _16979_/A2 _16979_/B1 vssd1 vssd1 vccd1 vccd1 _16913_/X sky130_fd_sc_hd__a21o_2
X_12036_ _12034_/Y _12036_/B vssd1 vssd1 vccd1 vccd1 _13431_/A sky130_fd_sc_hd__and2b_4
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1631 _09615_/Y vssd1 vssd1 vccd1 vccd1 _12137_/C1 sky130_fd_sc_hd__buf_8
X_17893_ _20664_/Q _17893_/A1 _17916_/S vssd1 vssd1 vccd1 vccd1 _20664_/D sky130_fd_sc_hd__mux2_1
XFILLER_239_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1642 _17494_/B vssd1 vssd1 vccd1 vccd1 _17486_/B sky130_fd_sc_hd__buf_6
Xfanout1653 _13978_/A2 vssd1 vssd1 vccd1 vccd1 _09664_/B sky130_fd_sc_hd__buf_4
XFILLER_238_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1664 _13863_/A vssd1 vssd1 vccd1 vccd1 _11261_/C sky130_fd_sc_hd__buf_6
X_19632_ _20438_/CLK _19632_/D vssd1 vssd1 vccd1 vccd1 _19632_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1675 _11239_/A1 vssd1 vssd1 vccd1 vccd1 _09672_/A sky130_fd_sc_hd__buf_8
X_16844_ _19227_/Q _16862_/A2 _16964_/B1 _19096_/Q _16843_/X vssd1 vssd1 vccd1 vccd1
+ _16844_/X sky130_fd_sc_hd__o221a_1
XFILLER_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1686 _12711_/A vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__buf_6
XFILLER_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1697 _10692_/A vssd1 vssd1 vccd1 vccd1 _12411_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_281_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19563_ _19574_/CLK _19563_/D vssd1 vssd1 vccd1 vccd1 _19563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16775_ _20402_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16775_/X sky130_fd_sc_hd__a21o_1
XFILLER_281_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13987_ _14035_/A1 _09664_/B _10115_/X _14035_/B1 _19844_/Q vssd1 vssd1 vccd1 vccd1
+ _14071_/C sky130_fd_sc_hd__o32a_1
XFILLER_218_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _18628_/B _18514_/B vssd1 vssd1 vccd1 vccd1 _18514_/X sky130_fd_sc_hd__or2_1
XFILLER_206_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15726_ _15973_/A1 _15725_/X _15713_/Y vssd1 vssd1 vccd1 vccd1 _15726_/X sky130_fd_sc_hd__a21o_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _19258_/Q _12964_/A2 _16945_/B _20006_/Q vssd1 vssd1 vccd1 vccd1 _14906_/B
+ sky130_fd_sc_hd__a22o_1
X_19494_ _21004_/CLK _19494_/D vssd1 vssd1 vccd1 vccd1 _19494_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18445_ _20877_/Q _18295_/Y _18449_/S vssd1 vssd1 vccd1 vccd1 _18446_/B sky130_fd_sc_hd__mux2_1
XFILLER_233_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15657_ _11497_/A _16057_/A2 _15654_/Y _15656_/X vssd1 vssd1 vccd1 vccd1 _15657_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _13389_/B _12869_/B vssd1 vssd1 vccd1 vccd1 _12869_/Y sky130_fd_sc_hd__nor2_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14608_ _19372_/Q _17892_/A1 _14632_/S vssd1 vssd1 vccd1 vccd1 _19372_/D sky130_fd_sc_hd__mux2_1
X_18376_ _20843_/Q _18375_/B _18375_/Y _18754_/A vssd1 vssd1 vccd1 vccd1 _20843_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15588_ _16005_/A1 _12718_/X _15587_/X _12716_/B vssd1 vssd1 vccd1 vccd1 _15588_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17327_ _20214_/Q _17327_/A2 _17302_/C _17326_/X _17330_/C1 vssd1 vssd1 vccd1 vccd1
+ _17327_/X sky130_fd_sc_hd__a221o_1
XFILLER_239_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14539_ _19309_/Q _17859_/A1 _14562_/S vssd1 vssd1 vccd1 vccd1 _19309_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17258_ _20191_/Q _17235_/Y _17279_/C1 vssd1 vssd1 vccd1 vccd1 _17258_/X sky130_fd_sc_hd__a21o_1
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16209_ _19632_/Q _17861_/A1 _16227_/S vssd1 vssd1 vccd1 vccd1 _19632_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17189_ _20153_/Q _17189_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20153_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_271_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_272_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _19086_/Q vssd1 vssd1 vccd1 vccd1 _09583_/B sky130_fd_sc_hd__inv_2
XFILLER_25_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20605_ _20641_/CLK _20605_/D vssd1 vssd1 vccd1 vccd1 _20605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20536_ _20668_/CLK _20536_/D vssd1 vssd1 vccd1 vccd1 _20536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20467_ _20467_/CLK _20467_/D vssd1 vssd1 vccd1 vccd1 _20467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ _10215_/X _10216_/X _10235_/S vssd1 vssd1 vccd1 vccd1 _10220_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20398_ _20759_/CLK _20398_/D vssd1 vssd1 vccd1 vccd1 _20398_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_161_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10151_ _19379_/Q _20670_/Q _11174_/S vssd1 vssd1 vccd1 vccd1 _10151_/X sky130_fd_sc_hd__mux2_1
XFILLER_267_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput291 _13833_/X vssd1 vssd1 vccd1 vccd1 addr0[6] sky130_fd_sc_hd__buf_4
XFILLER_248_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10082_ _10079_/X _10080_/X _10081_/X _12103_/A1 _10516_/S vssd1 vssd1 vccd1 vccd1
+ _10082_/X sky130_fd_sc_hd__a221o_1
XFILLER_181_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_275_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21019_ _21019_/CLK _21019_/D vssd1 vssd1 vccd1 vccd1 _21019_/Q sky130_fd_sc_hd__dfxtp_1
X_13910_ _19120_/Q _13919_/S _13909_/Y _18714_/A vssd1 vssd1 vccd1 vccd1 _19120_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14890_ _15610_/A1 _14889_/X _15610_/B1 vssd1 vssd1 vccd1 vccd1 _16053_/B sky130_fd_sc_hd__o21ai_4
XFILLER_236_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13841_ _20260_/Q _13840_/X _13839_/X vssd1 vssd1 vccd1 vccd1 _17226_/B sky130_fd_sc_hd__o21a_2
XFILLER_90_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16560_ _19846_/Q _16576_/A2 _16576_/B1 input16/X vssd1 vssd1 vccd1 vccd1 _16561_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13772_ _13777_/A _13772_/B vssd1 vssd1 vccd1 vccd1 _13772_/X sky130_fd_sc_hd__or2_1
XFILLER_250_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10984_ _12371_/A1 _19465_/Q _19433_/Q _11342_/S _11338_/A1 vssd1 vssd1 vccd1 vccd1
+ _10984_/X sky130_fd_sc_hd__a221o_1
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15511_ _20958_/Q _15568_/A2 _15568_/B1 _20830_/Q _15510_/X vssd1 vssd1 vccd1 vccd1
+ _15511_/X sky130_fd_sc_hd__a221o_4
XFILLER_271_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12723_ _12721_/Y _12722_/X _12709_/X _12716_/Y vssd1 vssd1 vccd1 vccd1 _12726_/C
+ sky130_fd_sc_hd__o211a_2
X_16491_ _19798_/Q _17886_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19798_/D sky130_fd_sc_hd__mux2_1
XFILLER_31_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18230_ _18508_/B vssd1 vssd1 vccd1 vccd1 _18230_/Y sky130_fd_sc_hd__clkinv_4
X_12654_ _19160_/Q _12479_/X _16005_/A1 _12513_/D vssd1 vssd1 vccd1 vccd1 _12662_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_31_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15442_ _15442_/A _15442_/B vssd1 vssd1 vccd1 vccd1 _15442_/Y sky130_fd_sc_hd__nand2_1
XFILLER_203_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _19286_/Q _20073_/Q _11965_/B vssd1 vssd1 vccd1 vccd1 _11605_/X sky130_fd_sc_hd__mux2_1
X_18161_ _20786_/Q _18160_/Y _18236_/S vssd1 vssd1 vccd1 vccd1 _18162_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12585_ _12588_/A _18765_/C _12585_/C _12588_/D vssd1 vssd1 vccd1 vccd1 _13193_/B
+ sky130_fd_sc_hd__or4_4
X_15373_ _15362_/Y _15372_/Y _15612_/S vssd1 vssd1 vccd1 vccd1 _15373_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17112_ _20082_/Q _17112_/A1 _17112_/S vssd1 vssd1 vccd1 vccd1 _20082_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14324_ _14323_/A _14323_/B _14323_/C vssd1 vssd1 vccd1 vccd1 _14333_/B sky130_fd_sc_hd__a21o_1
X_11536_ _12403_/A1 _13742_/A _12403_/B1 vssd1 vssd1 vccd1 vccd1 _11536_/X sky130_fd_sc_hd__o21a_1
X_18092_ _20771_/Q _18093_/C _20772_/Q vssd1 vssd1 vccd1 vccd1 _18094_/B sky130_fd_sc_hd__a21oi_1
XFILLER_239_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17043_ _17014_/A _17014_/B input252/X _17015_/B vssd1 vssd1 vccd1 vccd1 _17044_/C
+ sky130_fd_sc_hd__a31o_1
X_14255_ _14255_/A _16068_/B _14255_/C vssd1 vssd1 vccd1 vccd1 _14255_/X sky130_fd_sc_hd__or3_1
X_11467_ _11851_/A _20039_/Q _12011_/S _11458_/X vssd1 vssd1 vccd1 vccd1 _11467_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_137_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13206_ _13205_/A _19239_/Q _18752_/A _13205_/Y vssd1 vssd1 vccd1 vccd1 _13242_/C
+ sky130_fd_sc_hd__o211a_4
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10418_ _19505_/Q _15473_/A _11398_/S vssd1 vssd1 vccd1 vccd1 _10640_/B sky130_fd_sc_hd__mux2_8
X_14186_ _20273_/Q _14237_/A2 _14216_/B1 input244/X vssd1 vssd1 vccd1 vccd1 _14188_/B
+ sky130_fd_sc_hd__a22o_4
X_11398_ _19502_/Q _15380_/A _11398_/S vssd1 vssd1 vccd1 vccd1 _11404_/B sky130_fd_sc_hd__mux2_2
XFILLER_180_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13137_ _13135_/Y _13136_/X _20975_/Q _13370_/B vssd1 vssd1 vccd1 vccd1 _13137_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10349_ _11290_/A _20507_/Q _11292_/S0 _20539_/Q vssd1 vssd1 vccd1 vccd1 _10349_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18994_ _18180_/Y _18983_/B _19002_/B1 _18993_/X vssd1 vssd1 vccd1 vccd1 _21016_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13068_ _13590_/A _13591_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13605_/A sky130_fd_sc_hd__o21ba_2
X_17945_ _20714_/Q _17945_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20714_/D sky130_fd_sc_hd__mux2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1450 _09734_/Y vssd1 vssd1 vccd1 vccd1 _10611_/B sky130_fd_sc_hd__buf_6
X_12019_ _12016_/X _12018_/X _09776_/S vssd1 vssd1 vccd1 vccd1 _12019_/Y sky130_fd_sc_hd__a21oi_1
Xfanout1461 _09733_/Y vssd1 vssd1 vccd1 vccd1 _12088_/S sky130_fd_sc_hd__buf_6
XFILLER_238_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1472 _11033_/S vssd1 vssd1 vccd1 vccd1 _11297_/S sky130_fd_sc_hd__clkbuf_16
X_17876_ _20649_/Q _17876_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20649_/D sky130_fd_sc_hd__mux2_1
XFILLER_266_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1483 _09730_/Y vssd1 vssd1 vccd1 vccd1 _12426_/S sky130_fd_sc_hd__buf_12
X_19615_ _20425_/CLK _19615_/D vssd1 vssd1 vccd1 vccd1 _19615_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1494 _11895_/B vssd1 vssd1 vccd1 vccd1 _12131_/B sky130_fd_sc_hd__buf_6
X_16827_ _16805_/X _16824_/Y _16826_/X _16932_/A1 vssd1 vssd1 vccd1 vccd1 _16827_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_253_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19546_ _19617_/CLK _19546_/D vssd1 vssd1 vccd1 vccd1 _19546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16758_ _17008_/A1 _16757_/X _17008_/B1 vssd1 vssd1 vccd1 vccd1 _16758_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_253_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_253_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15709_ _13167_/A _15984_/A2 _15984_/B1 _13166_/A _15890_/A vssd1 vssd1 vccd1 vccd1
+ _15709_/X sky130_fd_sc_hd__a221o_1
X_19477_ _20702_/CLK _19477_/D vssd1 vssd1 vccd1 vccd1 _19477_/Q sky130_fd_sc_hd__dfxtp_1
X_16689_ _19944_/Q _17099_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19944_/D sky130_fd_sc_hd__mux2_1
XFILLER_181_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18428_ _18728_/A _18428_/B vssd1 vssd1 vccd1 vccd1 _20868_/D sky130_fd_sc_hd__and2_1
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18359_ _18517_/B _18363_/B vssd1 vssd1 vccd1 vccd1 _18359_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20321_ _20481_/CLK _20321_/D vssd1 vssd1 vccd1 vccd1 _20321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20252_ _20261_/CLK _20252_/D vssd1 vssd1 vccd1 vccd1 _20252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_135_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20183_ _20184_/CLK _20183_/D vssd1 vssd1 vccd1 vccd1 _20183_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09994_ _09992_/X _09993_/X _11849_/S vssd1 vssd1 vccd1 vccd1 _09994_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12370_ _09503_/A _12368_/X _12369_/X vssd1 vssd1 vccd1 vccd1 _12370_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_176_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11321_ _15264_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__or2_1
XFILLER_193_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20519_ _20683_/CLK _20519_/D vssd1 vssd1 vccd1 vccd1 _20519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14040_ _12512_/B _14040_/A2 _14040_/B1 _14039_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1
+ _19180_/D sky130_fd_sc_hd__o221a_1
X_11252_ _11258_/A1 _19334_/Q _20689_/Q _11257_/S _12519_/C vssd1 vssd1 vccd1 vccd1
+ _11252_/X sky130_fd_sc_hd__a221o_1
XFILLER_107_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10203_ _10203_/A _11236_/B vssd1 vssd1 vccd1 vccd1 _10203_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11183_ _12402_/A1 _17921_/A1 _11182_/X _13675_/A vssd1 vssd1 vccd1 vccd1 _13644_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10134_ _20378_/Q _20442_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _10134_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_267_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _20751_/Q _16011_/A2 _16011_/B1 _20783_/Q vssd1 vssd1 vccd1 vccd1 _15991_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17730_ _20511_/Q _17870_/A1 _17738_/S vssd1 vssd1 vccd1 vccd1 _20511_/D sky130_fd_sc_hd__mux2_1
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14942_ _15019_/B _14955_/B vssd1 vssd1 vccd1 vccd1 _15012_/B sky130_fd_sc_hd__nand2_4
X_10065_ _19378_/Q _10502_/A2 _10063_/X _11684_/A1 _10064_/X vssd1 vssd1 vccd1 vccd1
+ _10065_/X sky130_fd_sc_hd__o221a_1
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17661_ _20447_/Q _17695_/A1 _17669_/S vssd1 vssd1 vccd1 vccd1 _20447_/D sky130_fd_sc_hd__mux2_1
XFILLER_236_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14873_ _14868_/X _14872_/Y _15167_/S vssd1 vssd1 vccd1 vccd1 _14873_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19400_ _20559_/CLK _19400_/D vssd1 vssd1 vccd1 vccd1 _19400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16612_ _19871_/Q _17683_/A1 _16637_/S vssd1 vssd1 vccd1 vccd1 _19871_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13824_ _13826_/A1 _16235_/B _13826_/B1 _20622_/Q vssd1 vssd1 vccd1 vccd1 _13824_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_251_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17592_ _20350_/Q _17592_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20350_/D sky130_fd_sc_hd__mux2_1
XFILLER_245_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19331_ _20662_/CLK _19331_/D vssd1 vssd1 vccd1 vccd1 _19331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16543_ _16557_/A _16543_/B vssd1 vssd1 vccd1 vccd1 _19837_/D sky130_fd_sc_hd__or2_1
X_10967_ _10969_/B vssd1 vssd1 vccd1 vccd1 _11320_/B sky130_fd_sc_hd__inv_2
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13755_ _13780_/A _13755_/B vssd1 vssd1 vccd1 vccd1 _13755_/X sky130_fd_sc_hd__and2_1
XFILLER_189_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12706_ _12704_/X _12705_/Y _15703_/B2 vssd1 vssd1 vccd1 vccd1 _12706_/Y sky130_fd_sc_hd__a21oi_2
X_19262_ _20990_/CLK _19262_/D vssd1 vssd1 vccd1 vccd1 _19262_/Q sky130_fd_sc_hd__dfxtp_2
X_16474_ _19783_/Q _17937_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19783_/D sky130_fd_sc_hd__mux2_1
X_10898_ _20401_/Q _09689_/D _10895_/X _10896_/X _10897_/X vssd1 vssd1 vccd1 vccd1
+ _10898_/X sky130_fd_sc_hd__o221a_1
X_13686_ _13685_/A _13684_/Y _13685_/Y _13655_/A vssd1 vssd1 vccd1 vccd1 _13687_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_204_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18213_ _19538_/Q _18213_/B vssd1 vssd1 vccd1 vccd1 _18213_/Y sky130_fd_sc_hd__nand2b_4
X_15425_ _15019_/A _15414_/X _15424_/X vssd1 vssd1 vccd1 vccd1 _16815_/B sky130_fd_sc_hd__a21oi_4
XPHY_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19193_ _20341_/CLK _19193_/D vssd1 vssd1 vccd1 vccd1 _19193_/Q sky130_fd_sc_hd__dfxtp_1
X_12637_ _12519_/A _13589_/A1 _12633_/Y _12634_/Y vssd1 vssd1 vccd1 vccd1 _12698_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18144_ _18144_/A _18144_/B vssd1 vssd1 vccd1 vccd1 _18157_/A sky130_fd_sc_hd__nand2_2
X_12568_ _13730_/B _13776_/B1 _12567_/X _13740_/A vssd1 vssd1 vccd1 vccd1 _13443_/B
+ sky130_fd_sc_hd__o22a_4
X_15356_ _15356_/A vssd1 vssd1 vccd1 vccd1 _15356_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11519_ _11528_/S _11518_/X _11517_/X _12140_/C1 vssd1 vssd1 vccd1 vccd1 _11519_/X
+ sky130_fd_sc_hd__a211o_1
X_14307_ _14397_/A _14397_/B _14307_/C vssd1 vssd1 vccd1 vccd1 _14307_/X sky130_fd_sc_hd__or3_1
X_18075_ _20765_/Q _18077_/C _18074_/Y vssd1 vssd1 vccd1 vccd1 _20765_/D sky130_fd_sc_hd__o21a_1
X_15287_ _15402_/A _15287_/B vssd1 vssd1 vccd1 vccd1 _15287_/Y sky130_fd_sc_hd__nand2_1
X_12499_ _12664_/C _12498_/Y _13334_/A vssd1 vssd1 vccd1 vccd1 _12533_/A sky130_fd_sc_hd__a21oi_2
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17026_ _20004_/Q input213/X _17026_/S vssd1 vssd1 vccd1 vccd1 _20004_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14238_ _19506_/Q _14239_/B vssd1 vssd1 vccd1 vccd1 _14250_/A sky130_fd_sc_hd__nand2_1
XFILLER_160_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ _14157_/Y _14162_/B _14159_/B vssd1 vssd1 vccd1 vccd1 _14170_/B sky130_fd_sc_hd__o21ai_2
XFILLER_124_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout709 _13810_/A1 vssd1 vssd1 vccd1 vccd1 _13816_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_252_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18977_ _18687_/Y _18977_/A2 _18975_/Y _18976_/Y vssd1 vssd1 vccd1 vccd1 _18977_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _20697_/Q _17928_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20697_/D sky130_fd_sc_hd__mux2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1280 _09547_/X vssd1 vssd1 vccd1 vccd1 _16034_/S sky130_fd_sc_hd__buf_8
XFILLER_227_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1291 _15921_/B2 vssd1 vssd1 vccd1 vccd1 _12916_/B2 sky130_fd_sc_hd__buf_4
XFILLER_67_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17859_ _20632_/Q _17859_/A1 _17882_/S vssd1 vssd1 vccd1 vccd1 _20632_/D sky130_fd_sc_hd__mux2_1
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20870_ _21040_/CLK _20870_/D vssd1 vssd1 vccd1 vccd1 _20870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19529_ _19560_/CLK _19529_/D vssd1 vssd1 vccd1 vccd1 _19529_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_241_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_277_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20304_ _20565_/CLK _20304_/D vssd1 vssd1 vccd1 vccd1 _20304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20235_ _21043_/CLK _20235_/D vssd1 vssd1 vccd1 vccd1 _20235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20166_ _20573_/CLK _20166_/D vssd1 vssd1 vccd1 vccd1 _20166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09977_ _19287_/Q _20074_/Q _11965_/B vssd1 vssd1 vccd1 vccd1 _09977_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20097_ _20711_/CLK _20097_/D vssd1 vssd1 vccd1 vccd1 _20097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_217_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_58_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20559_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_603 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _11948_/A1 _11869_/X _11949_/S vssd1 vssd1 vccd1 vccd1 _11870_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_217_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_614 _13775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_625 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10821_ _12306_/A1 _20694_/Q _12300_/S _10820_/X vssd1 vssd1 vccd1 vccd1 _10821_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_232_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_636 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_647 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_260_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20999_ _21011_/CLK _20999_/D vssd1 vssd1 vccd1 vccd1 _20999_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ _10750_/X _10751_/X _12317_/S vssd1 vssd1 vccd1 vccd1 _10752_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13540_ _19661_/D _13537_/Y _13539_/Y _13663_/B vssd1 vssd1 vccd1 vccd1 _13540_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_214_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13471_ _19701_/Q _16279_/C vssd1 vssd1 vccd1 vccd1 _13472_/A sky130_fd_sc_hd__or2_4
X_10683_ _19177_/Q _11367_/B vssd1 vssd1 vccd1 vccd1 _10683_/X sky130_fd_sc_hd__or2_1
XFILLER_9_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12422_ _12419_/X _12421_/X _11118_/A vssd1 vssd1 vccd1 vccd1 _12422_/Y sky130_fd_sc_hd__a21oi_1
X_15210_ _19530_/Q _15402_/A _15209_/Y _16197_/A vssd1 vssd1 vccd1 vccd1 _19530_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16190_ _19619_/Q _15972_/X _16190_/S vssd1 vssd1 vccd1 vccd1 _16191_/B sky130_fd_sc_hd__mux2_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15141_ _20788_/Q _16047_/A2 _15021_/X input3/X _15140_/X vssd1 vssd1 vccd1 vccd1
+ _15141_/X sky130_fd_sc_hd__a221o_1
X_12353_ _12357_/A1 _12352_/X _12351_/X vssd1 vssd1 vccd1 vccd1 _12353_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_139_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11304_ _11302_/X _11303_/X _11304_/S vssd1 vssd1 vccd1 vccd1 _11304_/X sky130_fd_sc_hd__mux2_1
X_15072_ _15067_/S _11223_/B _14878_/B _15071_/X vssd1 vssd1 vccd1 vccd1 _15072_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12284_ _12284_/A _12284_/B vssd1 vssd1 vccd1 vccd1 _12286_/C sky130_fd_sc_hd__or2_1
X_14023_ _14029_/A1 _14038_/A2 _10555_/X _14035_/B1 _19856_/Q vssd1 vssd1 vccd1 vccd1
+ _14095_/C sky130_fd_sc_hd__o32a_1
X_18900_ _19137_/Q _18899_/X _18975_/A vssd1 vssd1 vccd1 vccd1 _18900_/X sky130_fd_sc_hd__mux2_1
X_11235_ _11235_/A _11326_/C vssd1 vssd1 vccd1 vccd1 _11235_/X sky130_fd_sc_hd__and2_1
XFILLER_84_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19880_ _20180_/CLK _19880_/D vssd1 vssd1 vccd1 vccd1 _19880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_268_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18831_ _19127_/Q _18949_/A2 _18949_/B1 vssd1 vssd1 vccd1 vccd1 _18831_/Y sky130_fd_sc_hd__a21oi_1
X_11166_ _20462_/Q _20302_/Q _12296_/S vssd1 vssd1 vccd1 vccd1 _11166_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xsplit2 split2/A vssd1 vssd1 vccd1 vccd1 split2/X sky130_fd_sc_hd__clkbuf_4
X_10117_ _19572_/Q _10116_/X _11243_/S vssd1 vssd1 vccd1 vccd1 _10117_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18762_ _20979_/Q _18756_/Y _18761_/X vssd1 vssd1 vccd1 vccd1 _18762_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11097_ _11012_/A _11096_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _11097_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15974_ _16051_/A1 _15960_/X _16051_/B1 vssd1 vssd1 vccd1 vccd1 _15974_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ _20494_/Q _17887_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20494_/D sky130_fd_sc_hd__mux2_1
XFILLER_212_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14925_ _18148_/S _12513_/D _18322_/A vssd1 vssd1 vccd1 vccd1 _14927_/A sky130_fd_sc_hd__a21o_2
X_10048_ _10046_/X _10047_/X _12071_/S vssd1 vssd1 vccd1 vccd1 _10048_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18693_ _20947_/Q _18165_/Y _18707_/S vssd1 vssd1 vccd1 vccd1 _18694_/B sky130_fd_sc_hd__mux2_1
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _20430_/Q _17678_/A1 _17674_/S vssd1 vssd1 vccd1 vccd1 _20430_/D sky130_fd_sc_hd__mux2_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14856_ _14855_/X _14848_/X _15215_/S vssd1 vssd1 vccd1 vccd1 _14856_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13807_ _13822_/A1 _13706_/B _13790_/X input222/X vssd1 vssd1 vccd1 vccd1 _13807_/X
+ sky130_fd_sc_hd__a22o_2
X_17575_ _20333_/Q _17852_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20333_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14787_ _19518_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14787_/X sky130_fd_sc_hd__or2_1
XFILLER_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _12157_/A1 _17913_/A1 _11998_/X vssd1 vssd1 vccd1 vccd1 _11999_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19314_ _20472_/CLK _19314_/D vssd1 vssd1 vccd1 vccd1 _19314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16526_ _16598_/A _16594_/C _16524_/Y _16567_/A vssd1 vssd1 vccd1 vccd1 _19830_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_91_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13738_ _13780_/A _13738_/B vssd1 vssd1 vccd1 vccd1 _13738_/X sky130_fd_sc_hd__and2_1
XFILLER_220_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19245_ _19246_/CLK _19245_/D vssd1 vssd1 vccd1 vccd1 _19245_/Q sky130_fd_sc_hd__dfxtp_4
X_16457_ _19766_/Q _17920_/A1 _16471_/S vssd1 vssd1 vccd1 vccd1 _19766_/D sky130_fd_sc_hd__mux2_1
XFILLER_188_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13669_ _16598_/C _13669_/B vssd1 vssd1 vccd1 vccd1 _13669_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15408_ _15295_/X _15407_/X _15578_/S vssd1 vssd1 vccd1 vccd1 _15409_/B sky130_fd_sc_hd__mux2_2
X_19176_ _19590_/CLK _19176_/D vssd1 vssd1 vccd1 vccd1 _19176_/Q sky130_fd_sc_hd__dfxtp_4
X_16388_ _19741_/Q _16388_/B vssd1 vssd1 vccd1 vccd1 _16394_/C sky130_fd_sc_hd__and2_2
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18127_ _20784_/Q _18125_/B _18126_/Y vssd1 vssd1 vccd1 vccd1 _20784_/D sky130_fd_sc_hd__o21a_1
XFILLER_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15339_ _20857_/Q _15338_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15339_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18058_ _20759_/Q _18061_/C _18056_/A vssd1 vssd1 vccd1 vccd1 _18058_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17009_ input67/X input102/X _17009_/S vssd1 vssd1 vccd1 vccd1 _17009_/X sky130_fd_sc_hd__mux2_8
X_09900_ _19288_/Q _20075_/Q _12149_/S vssd1 vssd1 vccd1 vccd1 _09900_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout506 _17794_/S vssd1 vssd1 vccd1 vccd1 _17811_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_98_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20020_ _20621_/CLK _20020_/D vssd1 vssd1 vccd1 vccd1 _20020_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_263_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09831_ _19645_/Q _19951_/Q _19289_/Q _20076_/Q _10621_/S _09834_/C vssd1 vssd1 vccd1
+ vccd1 _09831_/X sky130_fd_sc_hd__mux4_1
Xfanout517 _17676_/X vssd1 vssd1 vccd1 vccd1 _17703_/S sky130_fd_sc_hd__buf_4
Xfanout528 _17574_/X vssd1 vssd1 vccd1 vccd1 _17603_/S sky130_fd_sc_hd__buf_12
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout539 _17185_/X vssd1 vssd1 vccd1 vccd1 _17212_/S sky130_fd_sc_hd__buf_12
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09762_ _09752_/A _19485_/Q _19453_/Q _11936_/S _11946_/C1 vssd1 vssd1 vccd1 vccd1
+ _09762_/X sky130_fd_sc_hd__a221o_1
XFILLER_274_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_273_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09693_ _20580_/Q _11897_/B vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__or2_1
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20922_ _21019_/CLK _20922_/D vssd1 vssd1 vccd1 vccd1 _20922_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_254_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20853_ _20856_/CLK _20853_/D vssd1 vssd1 vccd1 vccd1 _20853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20784_ _21020_/CLK _20784_/D vssd1 vssd1 vccd1 vccd1 _20784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_176_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21009_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_105_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20861_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_175_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11020_ _11021_/A _19900_/Q _11035_/S _20025_/Q vssd1 vssd1 vccd1 vccd1 _11020_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20218_ _21022_/CLK _20218_/D vssd1 vssd1 vccd1 vccd1 _20218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20149_ _20720_/CLK _20149_/D vssd1 vssd1 vccd1 vccd1 _20149_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12971_ _19108_/Q _12971_/B _19113_/Q vssd1 vssd1 vccd1 vccd1 _12972_/D sky130_fd_sc_hd__or3b_1
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14710_ _19467_/Q _17857_/A1 _14719_/S vssd1 vssd1 vccd1 vccd1 _19467_/D sky130_fd_sc_hd__mux2_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11922_/A1 _11921_/Y _12158_/B1 vssd1 vssd1 vccd1 vccd1 _11922_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_218_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _20868_/Q _16042_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15690_/X sky130_fd_sc_hd__o21ba_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_400 _16811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_411 _18205_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_422 _10379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14641_ _19403_/Q _17925_/A1 _14667_/S vssd1 vssd1 vccd1 vccd1 _19403_/D sky130_fd_sc_hd__mux2_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_433 _13735_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11853_ _20421_/Q _20357_/Q _20649_/Q _20613_/Q _12165_/S _11846_/C vssd1 vssd1 vccd1
+ vccd1 _11853_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_444 _13755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_261_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_455 _19105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_466 _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _20228_/Q _17364_/A2 _17362_/B1 _20277_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17360_/X sky130_fd_sc_hd__a221o_1
XANTENNA_477 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ _13567_/A _10803_/Y _10802_/Y vssd1 vssd1 vccd1 vccd1 _10804_/Y sky130_fd_sc_hd__o21ai_4
X_14572_ _19338_/Q _17647_/A1 _14599_/S vssd1 vssd1 vccd1 vccd1 _19338_/D sky130_fd_sc_hd__mux2_1
XANTENNA_488 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11784_ _13694_/A _14878_/A vssd1 vssd1 vccd1 vccd1 _13658_/A sky130_fd_sc_hd__and2_4
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_499 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16311_ _19712_/Q _16314_/C _18086_/A vssd1 vssd1 vccd1 vccd1 _16311_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_213_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13523_ _13523_/A _13523_/B vssd1 vssd1 vccd1 vccd1 _13524_/A sky130_fd_sc_hd__xor2_4
X_17291_ _20202_/Q _17327_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17291_/X sky130_fd_sc_hd__a21o_1
X_10735_ _19668_/Q _20156_/Q _11074_/S vssd1 vssd1 vccd1 vccd1 _10735_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19030_ _18270_/Y _19046_/A2 _19048_/B1 _12551_/D _19046_/C1 vssd1 vssd1 vccd1 vccd1
+ _19030_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16242_ _18048_/A _16242_/B vssd1 vssd1 vccd1 vccd1 _19660_/D sky130_fd_sc_hd__nor2_1
X_10666_ _20632_/Q _20596_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _10666_/X sky130_fd_sc_hd__mux2_1
X_13454_ _13453_/A _13453_/B _13453_/C vssd1 vssd1 vccd1 vccd1 _13454_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_185_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12405_ _12411_/A _19927_/Q _11116_/S _20052_/Q vssd1 vssd1 vccd1 vccd1 _12405_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16173_ _16187_/A _16173_/B vssd1 vssd1 vccd1 vccd1 _19610_/D sky130_fd_sc_hd__and2_1
X_13385_ _20960_/Q _13607_/B _13383_/X _13384_/Y _18462_/A vssd1 vssd1 vccd1 vccd1
+ _13385_/Y sky130_fd_sc_hd__a221oi_4
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10597_ _19179_/Q _13653_/A _12577_/A vssd1 vssd1 vccd1 vccd1 _10597_/X sky130_fd_sc_hd__a21o_1
XFILLER_182_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15124_ _11140_/A _12465_/X _16030_/D1 vssd1 vssd1 vccd1 vccd1 _15124_/Y sky130_fd_sc_hd__a21oi_1
X_12336_ _12337_/A _20524_/Q _12339_/S0 _20556_/Q vssd1 vssd1 vccd1 vccd1 _12336_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_154_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12267_ _10692_/A _19491_/Q _19459_/Q _12268_/S _12419_/C1 vssd1 vssd1 vccd1 vccd1
+ _12267_/X sky130_fd_sc_hd__a221o_1
X_19932_ _20379_/CLK _19932_/D vssd1 vssd1 vccd1 vccd1 _19932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15055_ _14826_/X _14830_/X _15062_/S vssd1 vssd1 vccd1 vccd1 _15055_/X sky130_fd_sc_hd__mux2_2
XFILLER_268_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14006_ _19201_/Q _14083_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _14006_/X sky130_fd_sc_hd__mux2_1
X_11218_ _12275_/A _11209_/X _11217_/X _11201_/X vssd1 vssd1 vccd1 vccd1 _11218_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_268_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19863_ _20812_/CLK _19863_/D vssd1 vssd1 vccd1 vccd1 _19863_/Q sky130_fd_sc_hd__dfxtp_2
X_12198_ _12284_/A _12198_/B vssd1 vssd1 vccd1 vccd1 _12199_/B sky130_fd_sc_hd__nand2_2
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_269_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11149_ _09643_/A _09686_/D _11148_/Y _09586_/Y vssd1 vssd1 vccd1 vccd1 _11149_/X
+ sky130_fd_sc_hd__o211a_1
X_18814_ _18814_/A _18814_/B vssd1 vssd1 vccd1 vccd1 _20987_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19794_ _20677_/CLK _19794_/D vssd1 vssd1 vccd1 vccd1 _19794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18745_ _20973_/Q _18295_/Y _18749_/S vssd1 vssd1 vccd1 vccd1 _18746_/B sky130_fd_sc_hd__mux2_1
XFILLER_49_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15957_ _14882_/B _15177_/X _15182_/Y _12463_/B vssd1 vssd1 vccd1 vccd1 _15957_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput180 irq[3] vssd1 vssd1 vccd1 vccd1 _12549_/C sky130_fd_sc_hd__clkbuf_2
Xinput191 localMemory_wb_adr_i[10] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_hd__clkbuf_2
XFILLER_252_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14908_ _12944_/A _19176_/Q _14917_/A vssd1 vssd1 vccd1 vccd1 _14973_/A sky130_fd_sc_hd__mux2_2
XFILLER_236_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18676_ _18550_/X _18684_/A2 _18674_/Y _18675_/Y vssd1 vssd1 vccd1 vccd1 _18677_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _11955_/A _12115_/B _15984_/B1 _15887_/X vssd1 vssd1 vccd1 vccd1 _15888_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17627_ _20383_/Q _17695_/A1 _17635_/S vssd1 vssd1 vccd1 vccd1 _20383_/D sky130_fd_sc_hd__mux2_1
XFILLER_263_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14839_ _14835_/X _14838_/X _15067_/S vssd1 vssd1 vccd1 vccd1 _14839_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17558_ _20318_/Q _17903_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20318_/D sky130_fd_sc_hd__mux2_1
XFILLER_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20708_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_189_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16509_ _19816_/Q _17938_/A1 _16517_/S vssd1 vssd1 vccd1 vccd1 _19816_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17489_ _17495_/A1 _17488_/Y _18821_/A vssd1 vssd1 vccd1 vccd1 _20279_/D sky130_fd_sc_hd__a21oi_1
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19228_ _19228_/CLK _19228_/D vssd1 vssd1 vccd1 vccd1 _19228_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19159_ _19560_/CLK _19159_/D vssd1 vssd1 vccd1 vccd1 _19159_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_178_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20003_ _20004_/CLK _20003_/D vssd1 vssd1 vccd1 vccd1 _20003_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_143_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09814_ _19388_/Q _20679_/Q _11682_/S vssd1 vssd1 vccd1 vccd1 _09814_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09745_ _17538_/C _12342_/A _11305_/B _16454_/A vssd1 vssd1 vccd1 vccd1 _09746_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_274_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09676_/A _09676_/B vssd1 vssd1 vccd1 vccd1 _09676_/Y sky130_fd_sc_hd__nand2_2
XFILLER_215_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20905_ _21010_/CLK _20905_/D vssd1 vssd1 vccd1 vccd1 _20905_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20836_ _20998_/CLK _20836_/D vssd1 vssd1 vccd1 vccd1 _20836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20767_ _20796_/CLK _20767_/D vssd1 vssd1 vccd1 vccd1 _20767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10520_ _20311_/Q _11305_/B vssd1 vssd1 vccd1 vccd1 _10520_/X sky130_fd_sc_hd__or2_1
XFILLER_211_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20698_ _20698_/CLK _20698_/D vssd1 vssd1 vccd1 vccd1 _20698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_182_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10451_ _11368_/A1 _13680_/A _10450_/X _11398_/S vssd1 vssd1 vccd1 vccd1 _10455_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_148_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ _09863_/A _13414_/B _09862_/A vssd1 vssd1 vccd1 vccd1 _13413_/B sky130_fd_sc_hd__a21o_4
X_10382_ _11230_/A _10382_/B vssd1 vssd1 vccd1 vccd1 _10382_/Y sky130_fd_sc_hd__nand2_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12121_ _19893_/Q _19794_/Q _12121_/S vssd1 vssd1 vccd1 vccd1 _12121_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12052_ _19688_/Q _20176_/Q _12053_/S vssd1 vssd1 vccd1 vccd1 _12052_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1802 _16769_/S vssd1 vssd1 vccd1 vccd1 _16975_/S sky130_fd_sc_hd__buf_12
XFILLER_89_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1813 _14524_/B1 vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__clkbuf_4
X_11003_ _11268_/A _20057_/Q _11261_/C vssd1 vssd1 vccd1 vccd1 _11003_/X sky130_fd_sc_hd__and3_1
XFILLER_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1824 _12058_/S vssd1 vssd1 vccd1 vccd1 _12135_/A sky130_fd_sc_hd__buf_6
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1835 _11101_/A vssd1 vssd1 vccd1 vccd1 _12311_/A1 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_73_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20181_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_16860_ _16878_/A _16860_/B vssd1 vssd1 vccd1 vccd1 _16860_/Y sky130_fd_sc_hd__nand2_1
Xfanout1846 _11259_/S vssd1 vssd1 vccd1 vccd1 _09618_/A sky130_fd_sc_hd__buf_8
Xfanout1857 _10866_/A vssd1 vssd1 vccd1 vccd1 _12430_/S sky130_fd_sc_hd__buf_6
XFILLER_77_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout870 _15937_/A2 vssd1 vssd1 vccd1 vccd1 _16043_/A2 sky130_fd_sc_hd__buf_6
Xfanout1868 _12015_/A1 vssd1 vssd1 vccd1 vccd1 _11948_/A1 sky130_fd_sc_hd__buf_6
X_15811_ _15526_/B _15794_/Y _15810_/X _15526_/Y vssd1 vssd1 vccd1 vccd1 _15811_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout881 _16039_/B vssd1 vssd1 vccd1 vccd1 _15395_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_237_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1879 _19164_/Q vssd1 vssd1 vccd1 vccd1 _12510_/A sky130_fd_sc_hd__buf_6
XFILLER_120_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16791_ _16726_/X _16790_/Y _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16791_/X sky130_fd_sc_hd__a21o_2
Xfanout892 _18449_/S vssd1 vssd1 vccd1 vccd1 _18453_/S sky130_fd_sc_hd__buf_8
XFILLER_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18530_ _20903_/Q fanout750/X _18529_/X _18557_/B2 vssd1 vssd1 vccd1 vccd1 _18531_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_218_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15742_ _19722_/Q _15961_/A2 _15961_/B1 _19754_/Q vssd1 vssd1 vccd1 vccd1 _15742_/X
+ sky130_fd_sc_hd__a22o_1
X_12954_ _20021_/Q _20020_/Q vssd1 vssd1 vccd1 vccd1 _16716_/B sky130_fd_sc_hd__nand2b_4
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18461_ _18455_/X _18460_/X _18694_/A vssd1 vssd1 vccd1 vccd1 _20882_/D sky130_fd_sc_hd__o21a_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _11981_/C1 _11904_/X _11901_/X _12137_/C1 vssd1 vssd1 vccd1 vccd1 _11905_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_93_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15673_ _15026_/Y _15659_/X _15673_/B1 vssd1 vssd1 vccd1 vccd1 _15673_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_230 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12885_ _12483_/Y _12884_/Y _15870_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12885_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_252 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17412_ _17460_/A2 _17446_/A _17457_/B _20253_/Q vssd1 vssd1 vccd1 vccd1 _17412_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_263 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14624_ _19388_/Q _17908_/A1 _14628_/S vssd1 vssd1 vccd1 vccd1 _19388_/D sky130_fd_sc_hd__mux2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _18422_/A _18392_/B vssd1 vssd1 vccd1 vccd1 _20850_/D sky130_fd_sc_hd__and2_1
XFILLER_221_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11836_ _20046_/Q _19921_/Q _12139_/S vssd1 vssd1 vccd1 vccd1 _11836_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_274 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_296 input225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17343_ _20220_/Q _17363_/A2 _17342_/X _18702_/A vssd1 vssd1 vccd1 vccd1 _20220_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14555_ _19325_/Q _17107_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19325_/D sky130_fd_sc_hd__mux2_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _10645_/A _11772_/A _11408_/X _13425_/A vssd1 vssd1 vccd1 vccd1 _11768_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_14_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _20949_/Q _13519_/S _13504_/X _13505_/Y _18462_/A vssd1 vssd1 vccd1 vccd1
+ _13507_/C sky130_fd_sc_hd__a221o_1
XFILLER_147_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17274_ _20197_/Q _17280_/A2 _17272_/X _17273_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1
+ _20197_/D sky130_fd_sc_hd__o221a_1
XFILLER_202_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10718_ _10718_/A _10802_/B vssd1 vssd1 vccd1 vccd1 _10720_/B sky130_fd_sc_hd__nor2_4
X_14486_ _19094_/Q _16243_/B _14668_/B vssd1 vssd1 vccd1 vccd1 _17082_/A sky130_fd_sc_hd__or3_2
XFILLER_158_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11698_ _12102_/A1 _20136_/Q _20104_/Q _11698_/B2 vssd1 vssd1 vccd1 vccd1 _11698_/X
+ sky130_fd_sc_hd__a22o_1
X_19013_ _21026_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _19013_/X sky130_fd_sc_hd__or2_1
X_16225_ _19648_/Q _17911_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19648_/D sky130_fd_sc_hd__mux2_1
X_13437_ _13437_/A _13437_/B vssd1 vssd1 vccd1 vccd1 _16242_/B sky130_fd_sc_hd__or2_4
X_10649_ _12371_/A1 _19341_/Q _20696_/Q _12368_/S _12371_/C1 vssd1 vssd1 vccd1 vccd1
+ _10649_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16156_ _16833_/B _16164_/B vssd1 vssd1 vccd1 vccd1 _16156_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ _13368_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13368_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15107_ _14820_/X _14831_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15107_/X sky130_fd_sc_hd__mux2_1
X_12319_ _19654_/Q _12323_/S _12295_/X _12324_/S vssd1 vssd1 vccd1 vccd1 _12319_/X
+ sky130_fd_sc_hd__o211a_1
X_16087_ _19568_/Q _16081_/B _16087_/B1 vssd1 vssd1 vccd1 vccd1 _16087_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13299_ _13321_/B _13321_/C _13321_/A vssd1 vssd1 vccd1 vccd1 _13300_/C sky130_fd_sc_hd__a21o_1
XFILLER_170_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15038_ _14860_/X _14870_/X _15062_/S vssd1 vssd1 vccd1 vccd1 _15038_/X sky130_fd_sc_hd__mux2_1
X_19915_ _20679_/CLK _19915_/D vssd1 vssd1 vccd1 vccd1 _19915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19846_ _20014_/CLK _19846_/D vssd1 vssd1 vccd1 vccd1 _19846_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16989_ _17006_/A1 _16000_/X _16987_/X _16988_/X vssd1 vssd1 vccd1 vccd1 _16989_/X
+ sky130_fd_sc_hd__o211a_1
X_19777_ _20472_/CLK _19777_/D vssd1 vssd1 vccd1 vccd1 _19777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_271_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09530_ _18667_/B vssd1 vssd1 vccd1 vccd1 _09530_/Y sky130_fd_sc_hd__inv_2
X_18728_ _18728_/A _18728_/B vssd1 vssd1 vccd1 vccd1 _20964_/D sky130_fd_sc_hd__and2_1
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18659_ _19518_/Q _18683_/B vssd1 vssd1 vccd1 vccd1 _18659_/Y sky130_fd_sc_hd__nand2_1
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_280_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_269_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20621_ _20621_/CLK _20621_/D vssd1 vssd1 vccd1 vccd1 _20621_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20552_ _20706_/CLK _20552_/D vssd1 vssd1 vccd1 vccd1 _20552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20483_ _20579_/CLK _20483_/D vssd1 vssd1 vccd1 vccd1 _20483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput440 _19969_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[8] sky130_fd_sc_hd__buf_4
XFILLER_279_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput451 _19504_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[10] sky130_fd_sc_hd__buf_4
XFILLER_154_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput462 _19514_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[20] sky130_fd_sc_hd__buf_4
Xoutput473 _19524_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[30] sky130_fd_sc_hd__buf_4
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput484 _13823_/X vssd1 vssd1 vccd1 vccd1 wmask0[0] sky130_fd_sc_hd__buf_6
XFILLER_114_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1109 _17877_/A1 vssd1 vssd1 vccd1 vccd1 _17911_/A1 sky130_fd_sc_hd__buf_4
XFILLER_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21035_ _21042_/CLK _21035_/D vssd1 vssd1 vccd1 vccd1 _21035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_275_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_275_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ _19168_/Q _13863_/A vssd1 vssd1 vccd1 vccd1 _09728_/X sky130_fd_sc_hd__and2_4
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09659_ _10284_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _09659_/X sky130_fd_sc_hd__or2_4
XFILLER_216_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12670_ _19496_/Q _12758_/B vssd1 vssd1 vccd1 vccd1 _12674_/C sky130_fd_sc_hd__nand2_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_191_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19618_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _09752_/A _20137_/Q _20105_/Q _12013_/S vssd1 vssd1 vccd1 vccd1 _11621_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_120_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20816_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_20819_ _21013_/CLK _20819_/D vssd1 vssd1 vccd1 vccd1 _20819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14340_ _20288_/Q _14431_/A2 _14431_/B1 input229/X vssd1 vssd1 vccd1 vccd1 _14342_/B
+ sky130_fd_sc_hd__a22o_4
X_11552_ _12192_/A1 _11541_/X _11545_/X _11551_/X vssd1 vssd1 vccd1 vccd1 _11568_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ _11275_/A _10499_/X _10502_/X _12311_/C1 vssd1 vssd1 vccd1 vccd1 _10503_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11483_ _20382_/Q _20446_/Q _12188_/S vssd1 vssd1 vccd1 vccd1 _11483_/X sky130_fd_sc_hd__mux2_1
X_14271_ _14271_/A _14271_/B _14271_/C vssd1 vssd1 vccd1 vccd1 _14273_/A sky130_fd_sc_hd__and3_1
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16010_ _19732_/Q _14933_/Y _14935_/Y _19764_/Q vssd1 vssd1 vccd1 vccd1 _16010_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13222_ _19240_/Q _13231_/B _19241_/Q vssd1 vssd1 vccd1 vccd1 _13222_/X sky130_fd_sc_hd__a21o_1
X_10434_ _20344_/Q _11680_/C1 _12043_/B _12063_/C1 vssd1 vssd1 vccd1 vccd1 _10434_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_137_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10365_ _10365_/A _11414_/B vssd1 vssd1 vccd1 vccd1 _15580_/S sky130_fd_sc_hd__nand2_4
X_13153_ _13596_/A _13596_/B _15410_/S vssd1 vssd1 vccd1 vccd1 _13611_/B sky130_fd_sc_hd__a21oi_4
XFILLER_163_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12104_ _12828_/A _12099_/Y _12101_/Y _12103_/Y _12850_/A1 vssd1 vssd1 vccd1 vccd1
+ _12104_/X sky130_fd_sc_hd__a221o_1
X_17961_ _17961_/A _17961_/B vssd1 vssd1 vccd1 vccd1 _20724_/D sky130_fd_sc_hd__nor2_1
X_13084_ _13017_/Y _13195_/A _13194_/B vssd1 vssd1 vccd1 vccd1 _13084_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10296_ _20379_/Q _20443_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _10296_/X sky130_fd_sc_hd__mux2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1610 _09618_/Y vssd1 vssd1 vccd1 vccd1 _11094_/S sky130_fd_sc_hd__buf_6
X_16912_ _19980_/Q _16876_/A _16911_/Y _18795_/A vssd1 vssd1 vccd1 vccd1 _19980_/D
+ sky130_fd_sc_hd__a211o_1
X_12035_ _12035_/A _12035_/B vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__nand2_1
X_19700_ _20451_/CLK _19700_/D vssd1 vssd1 vccd1 vccd1 _19700_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1621 _10322_/S vssd1 vssd1 vccd1 vccd1 _10235_/S sky130_fd_sc_hd__buf_6
XFILLER_104_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17892_ _20663_/Q _17892_/A1 _17916_/S vssd1 vssd1 vccd1 vccd1 _20663_/D sky130_fd_sc_hd__mux2_1
XFILLER_214_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1632 _09615_/Y vssd1 vssd1 vccd1 vccd1 _12059_/C1 sky130_fd_sc_hd__buf_6
Xfanout1643 _12922_/X vssd1 vssd1 vccd1 vccd1 _17494_/B sky130_fd_sc_hd__buf_6
Xfanout1654 _09662_/Y vssd1 vssd1 vccd1 vccd1 _13978_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19631_ _20633_/CLK _19631_/D vssd1 vssd1 vccd1 vccd1 _19631_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1665 _12464_/C vssd1 vssd1 vccd1 vccd1 _13863_/A sky130_fd_sc_hd__buf_12
X_16843_ _20409_/Q _17004_/A2 _17004_/B1 vssd1 vssd1 vccd1 vccd1 _16843_/X sky130_fd_sc_hd__a21o_1
XFILLER_266_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_238_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1676 _09516_/Y vssd1 vssd1 vccd1 vccd1 _11239_/A1 sky130_fd_sc_hd__buf_8
XFILLER_266_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1687 _12711_/A vssd1 vssd1 vccd1 vccd1 _12084_/A sky130_fd_sc_hd__buf_4
Xfanout1698 _12254_/A vssd1 vssd1 vccd1 vccd1 _10692_/A sky130_fd_sc_hd__buf_6
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_266_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19562_ _19574_/CLK _19562_/D vssd1 vssd1 vccd1 vccd1 _19562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16774_ _16869_/A _16774_/B vssd1 vssd1 vccd1 vccd1 _16774_/Y sky130_fd_sc_hd__nand2_1
XFILLER_281_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13986_ _12510_/C _13986_/A2 _14004_/B1 _13985_/X _16143_/A vssd1 vssd1 vccd1 vccd1
+ _19162_/D sky130_fd_sc_hd__o221a_1
XFILLER_253_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18513_ _18891_/A _18513_/B vssd1 vssd1 vccd1 vccd1 _20897_/D sky130_fd_sc_hd__nor2_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15725_ _15882_/A1 _15714_/X _15715_/X _15724_/X vssd1 vssd1 vccd1 vccd1 _15725_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19493_ _20155_/CLK _19493_/D vssd1 vssd1 vccd1 vccd1 _19493_/Q sky130_fd_sc_hd__dfxtp_1
X_12937_ _19255_/Q _12964_/A2 _16945_/B _20003_/Q vssd1 vssd1 vccd1 vccd1 _12944_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_208_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20585_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18444_ _18746_/A _18444_/B vssd1 vssd1 vccd1 vccd1 _20876_/D sky130_fd_sc_hd__and2_1
XFILLER_222_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15656_ _15983_/A _15578_/X _15655_/X vssd1 vssd1 vccd1 vccd1 _15656_/X sky130_fd_sc_hd__a21o_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12868_ _12808_/B _12820_/B _12906_/A vssd1 vssd1 vccd1 vccd1 _12869_/B sky130_fd_sc_hd__o21a_1
XFILLER_222_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _19371_/Q _17891_/A1 _14632_/S vssd1 vssd1 vccd1 vccd1 _19371_/D sky130_fd_sc_hd__mux2_1
XFILLER_222_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ _19686_/Q _20174_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _11819_/X sky130_fd_sc_hd__mux2_1
X_18375_ _18541_/B _18375_/B vssd1 vssd1 vccd1 vccd1 _18375_/Y sky130_fd_sc_hd__nand2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15587_ _15544_/A _15576_/X _15586_/Y _15527_/B vssd1 vssd1 vccd1 vccd1 _15587_/X
+ sky130_fd_sc_hd__o22a_1
X_12799_ _19515_/Q _12811_/A vssd1 vssd1 vccd1 vccd1 _12800_/B sky130_fd_sc_hd__nor2_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17326_ input7/X _15133_/A _17329_/S vssd1 vssd1 vccd1 vccd1 _17326_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14538_ _19308_/Q _17683_/A1 _14562_/S vssd1 vssd1 vccd1 vccd1 _19308_/D sky130_fd_sc_hd__mux2_1
XFILLER_186_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17257_ _17257_/A _17275_/B _17269_/C vssd1 vssd1 vccd1 vccd1 _17257_/X sky130_fd_sc_hd__and3_1
X_14469_ _20230_/Q _19259_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14470_/B sky130_fd_sc_hd__mux2_1
X_16208_ _19631_/Q _17894_/A1 _16230_/S vssd1 vssd1 vccd1 vccd1 _19631_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17188_ _20152_/Q _17922_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20152_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16139_ _19593_/Q _16164_/B _16138_/Y _16165_/C1 vssd1 vssd1 vccd1 vccd1 _19593_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19829_ _20085_/CLK _19829_/D vssd1 vssd1 vccd1 vccd1 _19829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_272_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09513_ _19087_/Q vssd1 vssd1 vccd1 vccd1 _09583_/A sky130_fd_sc_hd__inv_2
XFILLER_271_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_262_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20604_ _20672_/CLK _20604_/D vssd1 vssd1 vccd1 vccd1 _20604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20535_ _20635_/CLK _20535_/D vssd1 vssd1 vccd1 vccd1 _20535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20466_ _20630_/CLK _20466_/D vssd1 vssd1 vccd1 vccd1 _20466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20397_ _20667_/CLK _20397_/D vssd1 vssd1 vccd1 vccd1 _20397_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_133_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ _20410_/Q _20346_/Q _10924_/S vssd1 vssd1 vccd1 vccd1 _10150_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput292 _13834_/X vssd1 vssd1 vccd1 vccd1 addr0[7] sky130_fd_sc_hd__buf_4
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _09829_/A _19474_/Q _19442_/Q _10400_/S vssd1 vssd1 vccd1 vccd1 _10081_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_102_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21018_ _21018_/CLK _21018_/D vssd1 vssd1 vccd1 vccd1 _21018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_263_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _20261_/Q _20258_/Q _20257_/Q _20259_/Q vssd1 vssd1 vccd1 vccd1 _13840_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_47_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_251_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ _12402_/Y _13730_/B _13776_/B1 vssd1 vssd1 vccd1 vccd1 _13774_/A sky130_fd_sc_hd__o21a_2
XFILLER_250_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10983_ _19868_/Q _19769_/Q _10983_/S vssd1 vssd1 vccd1 vccd1 _10983_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15510_ _20926_/Q _15567_/A2 _15509_/X vssd1 vssd1 vccd1 vccd1 _15510_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ _19508_/Q _12758_/B vssd1 vssd1 vccd1 vccd1 _12722_/X sky130_fd_sc_hd__and2_1
X_16490_ _17919_/A _17574_/B _16490_/C vssd1 vssd1 vccd1 vccd1 _16490_/X sky130_fd_sc_hd__and3_4
XFILLER_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15441_ _13155_/A _14878_/B _15440_/X vssd1 vssd1 vccd1 vccd1 _15441_/X sky130_fd_sc_hd__a21bo_1
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12653_ _12653_/A _12653_/B _12653_/C vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__nor3_2
XFILLER_169_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18160_ _18459_/B vssd1 vssd1 vccd1 vccd1 _18160_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _20041_/Q _19916_/Q _11965_/B vssd1 vssd1 vccd1 vccd1 _11604_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15372_ _15372_/A vssd1 vssd1 vccd1 vccd1 _15372_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12584_ _12584_/A _12584_/B _12584_/C vssd1 vssd1 vccd1 vccd1 _12588_/D sky130_fd_sc_hd__or3_1
XFILLER_129_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17111_ _20081_/Q _17111_/A1 _17111_/S vssd1 vssd1 vccd1 vccd1 _20081_/D sky130_fd_sc_hd__mux2_1
X_14323_ _14323_/A _14323_/B _14323_/C vssd1 vssd1 vccd1 vccd1 _14325_/B sky130_fd_sc_hd__and3_1
X_18091_ _20771_/Q _18093_/C _18090_/Y vssd1 vssd1 vccd1 vccd1 _20771_/D sky130_fd_sc_hd__o21a_1
X_11535_ _12157_/A1 _11534_/X _11531_/X _12153_/B1 vssd1 vssd1 vccd1 vccd1 _13742_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_129_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17042_ _20020_/Q _16706_/X _20021_/Q vssd1 vssd1 vccd1 vccd1 _17044_/B sky130_fd_sc_hd__o21ai_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14254_ _14275_/A1 _14253_/X _13294_/Y vssd1 vssd1 vccd1 vccd1 _14255_/C sky130_fd_sc_hd__o21a_1
XFILLER_139_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11466_ _11846_/C _11461_/X _11465_/X _11872_/A vssd1 vssd1 vccd1 vccd1 _11466_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_109_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13205_ _13205_/A _13205_/B vssd1 vssd1 vccd1 vccd1 _13205_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10417_ _12107_/A1 split4/A _10416_/X _12194_/B2 vssd1 vssd1 vccd1 vccd1 _15473_/A
+ sky130_fd_sc_hd__a22o_4
X_11397_ _12277_/A1 _11397_/A2 _11396_/X _11397_/B2 vssd1 vssd1 vccd1 vccd1 _15380_/A
+ sky130_fd_sc_hd__a22o_4
X_14185_ _19221_/Q _14256_/A2 _14183_/X _14184_/X _14185_/C1 vssd1 vssd1 vccd1 vccd1
+ _19221_/D sky130_fd_sc_hd__o221a_1
XFILLER_140_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13136_ _13135_/A _13135_/B _13370_/B vssd1 vssd1 vccd1 vccd1 _13136_/X sky130_fd_sc_hd__a21o_1
XFILLER_225_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10348_ _10260_/S _10347_/X _12342_/A vssd1 vssd1 vccd1 vccd1 _10348_/X sky130_fd_sc_hd__o21a_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _21016_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _18993_/X sky130_fd_sc_hd__or2_1
XFILLER_152_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13067_ _13047_/X _13066_/X _13048_/Y vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__a21boi_4
X_17944_ _20713_/Q _17944_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20713_/D sky130_fd_sc_hd__mux2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _13422_/A vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__clkinv_2
XFILLER_94_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1440 _12412_/B2 vssd1 vssd1 vccd1 vccd1 _09738_/A sky130_fd_sc_hd__buf_12
XFILLER_66_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12018_ _20328_/Q _12025_/S _12017_/X vssd1 vssd1 vccd1 vccd1 _12018_/X sky130_fd_sc_hd__a21o_1
Xfanout1451 _11021_/C vssd1 vssd1 vccd1 vccd1 _11290_/C sky130_fd_sc_hd__buf_6
XFILLER_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17875_ _20648_/Q _17909_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20648_/D sky130_fd_sc_hd__mux2_1
Xfanout1462 _09733_/Y vssd1 vssd1 vccd1 vccd1 _12258_/S sky130_fd_sc_hd__buf_12
XFILLER_226_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1473 _11204_/S vssd1 vssd1 vccd1 vccd1 _11033_/S sky130_fd_sc_hd__buf_12
XFILLER_238_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1484 _12105_/A vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__buf_8
XFILLER_254_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19614_ _20425_/CLK _19614_/D vssd1 vssd1 vccd1 vccd1 _19614_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1495 _12041_/B vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_285_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16826_ _19225_/Q _16862_/A2 _17005_/A2 _19094_/Q _16825_/X vssd1 vssd1 vccd1 vccd1
+ _16826_/X sky130_fd_sc_hd__o221a_1
XFILLER_65_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_235_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16757_ _19218_/Q _16862_/A2 _16713_/X _16754_/Y _16756_/X vssd1 vssd1 vccd1 vccd1
+ _16757_/X sky130_fd_sc_hd__o2111a_1
XFILLER_19_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19545_ _19618_/CLK _19545_/D vssd1 vssd1 vccd1 vccd1 _19545_/Q sky130_fd_sc_hd__dfxtp_1
X_13969_ _14035_/A1 _13969_/A2 _09656_/X _14035_/B1 _19838_/Q vssd1 vssd1 vccd1 vccd1
+ _14059_/C sky130_fd_sc_hd__o32a_1
XFILLER_34_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_281_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15708_ _11882_/Y _15981_/B _15707_/X vssd1 vssd1 vccd1 vccd1 _15708_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19476_ _20703_/CLK _19476_/D vssd1 vssd1 vccd1 vccd1 _19476_/Q sky130_fd_sc_hd__dfxtp_1
X_16688_ _19943_/Q _17900_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19943_/D sky130_fd_sc_hd__mux2_1
XFILLER_221_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_221_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18427_ _20868_/Q _18250_/Y _18449_/S vssd1 vssd1 vccd1 vccd1 _18428_/B sky130_fd_sc_hd__mux2_1
X_15639_ _16046_/A1 _15638_/X _15634_/X vssd1 vssd1 vccd1 vccd1 _15639_/X sky130_fd_sc_hd__o21a_2
XFILLER_221_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18358_ _20834_/Q _18357_/B _18357_/Y _18724_/A vssd1 vssd1 vccd1 vccd1 _20834_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_194_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17309_ _20208_/Q _17321_/A2 _17305_/C _17308_/X _17330_/C1 vssd1 vssd1 vccd1 vccd1
+ _17309_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18289_ _18299_/A1 _14383_/B _18288_/Y vssd1 vssd1 vccd1 vccd1 _18544_/B sky130_fd_sc_hd__o21ai_4
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20320_ _20480_/CLK _20320_/D vssd1 vssd1 vccd1 vccd1 _20320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20251_ _20261_/CLK _20251_/D vssd1 vssd1 vccd1 vccd1 _20251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20182_ _20184_/CLK _20182_/D vssd1 vssd1 vccd1 vccd1 _20182_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_89_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _20417_/Q _20353_/Q _20645_/Q _20609_/Q _12188_/S _11851_/C vssd1 vssd1 vccd1
+ vccd1 _09993_/X sky130_fd_sc_hd__mux4_1
XFILLER_276_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_272_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ _15578_/S _11320_/B vssd1 vssd1 vccd1 vccd1 _11776_/B sky130_fd_sc_hd__nand2_1
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20518_ _20682_/CLK _20518_/D vssd1 vssd1 vccd1 vccd1 _20518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11251_ _19398_/Q _20557_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _11251_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20449_ _20481_/CLK _20449_/D vssd1 vssd1 vccd1 vccd1 _20449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10202_ _09676_/Y _10465_/A _10032_/Y vssd1 vssd1 vccd1 vccd1 _10202_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182_ _12311_/C1 _11165_/X _11181_/X _12401_/A1 vssd1 vssd1 vccd1 vccd1 _11182_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10133_ _20474_/Q _20314_/Q _11257_/S vssd1 vssd1 vccd1 vccd1 _10133_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ _19731_/Q _15990_/B vssd1 vssd1 vccd1 vccd1 _15990_/X sky130_fd_sc_hd__or2_1
XFILLER_0_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14941_ _15314_/B _14980_/B _15314_/C vssd1 vssd1 vccd1 vccd1 _14941_/X sky130_fd_sc_hd__or3_4
X_10064_ _12060_/A1 _20669_/Q _11680_/C1 _09806_/S vssd1 vssd1 vccd1 vccd1 _10064_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17660_ _20446_/Q _17903_/A1 _17671_/S vssd1 vssd1 vccd1 vccd1 _20446_/D sky130_fd_sc_hd__mux2_1
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14872_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16611_ _19870_/Q _17857_/A1 _16620_/S vssd1 vssd1 vccd1 vccd1 _19870_/D sky130_fd_sc_hd__mux2_1
X_13823_ _13826_/A1 _16233_/B _13826_/B1 _20621_/Q vssd1 vssd1 vccd1 vccd1 _13823_/X
+ sky130_fd_sc_hd__a22o_4
X_17591_ _20349_/Q _17902_/A1 _17603_/S vssd1 vssd1 vccd1 vccd1 _20349_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16542_ _19837_/Q _16576_/A2 _16576_/B1 input38/X vssd1 vssd1 vccd1 vccd1 _16543_/B
+ sky130_fd_sc_hd__o22a_1
X_19330_ _20075_/CLK _19330_/D vssd1 vssd1 vccd1 vccd1 _19330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ _13754_/A _13754_/B vssd1 vssd1 vccd1 vccd1 _13755_/B sky130_fd_sc_hd__nor2_8
XFILLER_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10966_ _15150_/C1 _12682_/A _10935_/Y vssd1 vssd1 vccd1 vccd1 _10969_/B sky130_fd_sc_hd__o21bai_4
XFILLER_44_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19261_ _21022_/CLK _19261_/D vssd1 vssd1 vccd1 vccd1 _19261_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _15593_/A _12731_/B vssd1 vssd1 vccd1 vccd1 _12705_/Y sky130_fd_sc_hd__nand2_1
X_16473_ _19782_/Q _17936_/A1 _16485_/S vssd1 vssd1 vccd1 vccd1 _19782_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13685_ _13685_/A _13685_/B vssd1 vssd1 vccd1 vccd1 _13685_/Y sky130_fd_sc_hd__nor2_2
X_10897_ _20337_/Q _09623_/B _10897_/A3 _11170_/B1 vssd1 vssd1 vccd1 vccd1 _10897_/X
+ sky130_fd_sc_hd__o31a_1
X_18212_ _18416_/A _18212_/B vssd1 vssd1 vccd1 vccd1 _20796_/D sky130_fd_sc_hd__and2_1
XFILLER_231_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15424_ _19711_/Q _15423_/X _15454_/S vssd1 vssd1 vccd1 vccd1 _15424_/X sky130_fd_sc_hd__mux2_2
XFILLER_188_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19192_ _19560_/CLK _19192_/D vssd1 vssd1 vccd1 vccd1 _19192_/Q sky130_fd_sc_hd__dfxtp_1
X_12636_ _12633_/Y _12634_/Y _12519_/A _13589_/A1 vssd1 vssd1 vccd1 vccd1 _12636_/Y
+ sky130_fd_sc_hd__o211ai_1
XPHY_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18143_ _12944_/C _19112_/Q _18149_/S vssd1 vssd1 vccd1 vccd1 _18144_/B sky130_fd_sc_hd__mux2_1
XFILLER_200_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15355_ _15159_/Y _15168_/Y _15357_/S vssd1 vssd1 vccd1 vccd1 _15356_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12567_ _14897_/A _13698_/B _15075_/A vssd1 vssd1 vccd1 vccd1 _12567_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14306_ _14306_/A1 _14305_/X _13330_/X vssd1 vssd1 vccd1 vccd1 _14307_/C sky130_fd_sc_hd__o21a_1
X_18074_ _20765_/Q _18077_/C _18080_/A vssd1 vssd1 vccd1 vccd1 _18074_/Y sky130_fd_sc_hd__a21oi_1
X_11518_ _20641_/Q _20605_/Q _12133_/S vssd1 vssd1 vccd1 vccd1 _11518_/X sky130_fd_sc_hd__mux2_1
X_15286_ _10935_/B _15266_/X _15285_/X _10851_/Y vssd1 vssd1 vccd1 vccd1 _15287_/B
+ sky130_fd_sc_hd__a31o_1
X_12498_ _12498_/A _12498_/B vssd1 vssd1 vccd1 vccd1 _12498_/Y sky130_fd_sc_hd__xnor2_1
X_17025_ _20003_/Q input212/X _17026_/S vssd1 vssd1 vccd1 vccd1 _20003_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14237_ _20278_/Q _14237_/A2 _14267_/B1 input218/X vssd1 vssd1 vccd1 vccd1 _14239_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_109_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11449_ _12140_/C1 _11448_/X _11445_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _11449_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14168_ _19499_/Q _14171_/B vssd1 vssd1 vccd1 vccd1 _14170_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_259_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13119_ _13115_/X _13117_/X _13118_/X vssd1 vssd1 vccd1 vccd1 _13119_/X sky130_fd_sc_hd__a21o_1
XFILLER_285_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14099_ _14099_/A _14099_/B _14099_/C vssd1 vssd1 vccd1 vccd1 _14099_/X sky130_fd_sc_hd__or3_1
X_18976_ _19148_/Q _18976_/A2 _18767_/B vssd1 vssd1 vccd1 vccd1 _18976_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_252_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17927_ _20696_/Q _17927_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20696_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1270 _09607_/X vssd1 vssd1 vccd1 vccd1 _09613_/B sky130_fd_sc_hd__buf_6
XFILLER_267_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1281 _11398_/S vssd1 vssd1 vccd1 vccd1 _15589_/S sky130_fd_sc_hd__buf_6
X_17858_ _20631_/Q _17892_/A1 _17882_/S vssd1 vssd1 vccd1 vccd1 _20631_/D sky130_fd_sc_hd__mux2_1
XFILLER_254_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1292 _16062_/B2 vssd1 vssd1 vccd1 vccd1 _15921_/B2 sky130_fd_sc_hd__buf_2
XFILLER_227_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16809_ _19701_/Q _19697_/Q vssd1 vssd1 vccd1 vccd1 _16809_/X sky130_fd_sc_hd__and2_4
XFILLER_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17789_ _20566_/Q _17929_/A1 _17806_/S vssd1 vssd1 vccd1 vccd1 _20566_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19528_ _19603_/CLK _19528_/D vssd1 vssd1 vccd1 vccd1 _19528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19459_ _20468_/CLK _19459_/D vssd1 vssd1 vccd1 vccd1 _19459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20303_ _20463_/CLK _20303_/D vssd1 vssd1 vccd1 vccd1 _20303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20234_ _21026_/CLK _20234_/D vssd1 vssd1 vccd1 vccd1 _20234_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20165_ _20570_/CLK _20165_/D vssd1 vssd1 vccd1 vccd1 _20165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ _20042_/Q _19917_/Q _12121_/S vssd1 vssd1 vccd1 vccd1 _09976_/X sky130_fd_sc_hd__mux2_1
XFILLER_249_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_265_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20096_ _21047_/A _20096_/D vssd1 vssd1 vccd1 vccd1 _20096_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_273_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_604 _20621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_615 _13775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_626 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10820_ _09618_/A _12230_/A1 _19339_/Q _12302_/S vssd1 vssd1 vccd1 vccd1 _10820_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_637 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_648 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ _20998_/CLK _20998_/D vssd1 vssd1 vccd1 vccd1 _20998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_260_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_98_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20760_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10751_ _19372_/Q _20663_/Q _11161_/S vssd1 vssd1 vccd1 vccd1 _10751_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20671_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13470_ _16716_/B _13473_/B vssd1 vssd1 vccd1 vccd1 _16279_/C sky130_fd_sc_hd__nand2_2
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10682_ _12245_/A1 _17893_/A1 _10679_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _13661_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ _20331_/Q _12268_/S _12420_/X vssd1 vssd1 vccd1 vccd1 _12421_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15140_ _20978_/Q _15139_/X _15140_/S vssd1 vssd1 vccd1 vccd1 _15140_/X sky130_fd_sc_hd__mux2_4
X_12352_ _19896_/Q _19797_/Q _12352_/S vssd1 vssd1 vccd1 vccd1 _12352_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11303_ _19865_/Q _19766_/Q _11303_/S vssd1 vssd1 vccd1 vccd1 _11303_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15071_ _12470_/Y _15500_/A0 _15071_/S vssd1 vssd1 vccd1 vccd1 _15071_/X sky130_fd_sc_hd__mux2_1
X_12283_ _12283_/A _12283_/B vssd1 vssd1 vccd1 vccd1 _13182_/A sky130_fd_sc_hd__nor2_8
XFILLER_135_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14022_ _10831_/S _14043_/A2 _14040_/B1 _14021_/X _14104_/C1 vssd1 vssd1 vccd1 vccd1
+ _19174_/D sky130_fd_sc_hd__o221a_1
XFILLER_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11234_ _11234_/A _11234_/B _11233_/X vssd1 vssd1 vccd1 vccd1 _11326_/C sky130_fd_sc_hd__or3b_1
XFILLER_181_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_268_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18830_ _18830_/A _18830_/B vssd1 vssd1 vccd1 vccd1 _18830_/Y sky130_fd_sc_hd__nand2_1
XFILLER_267_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11165_ _09689_/C _11155_/X _11158_/X _11164_/X vssd1 vssd1 vccd1 vccd1 _11165_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10116_ _11228_/A1 _09664_/B _10115_/X _11242_/B1 _19844_/Q vssd1 vssd1 vccd1 vccd1
+ _10116_/X sky130_fd_sc_hd__o32a_1
XFILLER_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xsplit3 split3/A vssd1 vssd1 vccd1 vccd1 split3/X sky130_fd_sc_hd__buf_4
X_11096_ _12400_/A1 _11088_/X _11095_/X _11080_/X vssd1 vssd1 vccd1 vccd1 _11096_/X
+ sky130_fd_sc_hd__o31a_4
X_18761_ _18486_/Y _18756_/B _18760_/X vssd1 vssd1 vccd1 vccd1 _18761_/X sky130_fd_sc_hd__a21o_1
XFILLER_49_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15973_ _15973_/A1 _15972_/X _15960_/X vssd1 vssd1 vccd1 vccd1 _15973_/X sky130_fd_sc_hd__a21o_1
XFILLER_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14924_ _18163_/A _16719_/B vssd1 vssd1 vccd1 vccd1 _18322_/A sky130_fd_sc_hd__and2b_2
X_17712_ _20493_/Q _17852_/A1 _17743_/S vssd1 vssd1 vccd1 vccd1 _20493_/D sky130_fd_sc_hd__mux2_1
X_10047_ _19674_/Q _20162_/Q _10425_/S vssd1 vssd1 vccd1 vccd1 _10047_/X sky130_fd_sc_hd__mux2_1
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18692_ _18692_/A _18692_/B vssd1 vssd1 vccd1 vccd1 _20946_/D sky130_fd_sc_hd__and2_1
XFILLER_49_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17643_ _20429_/Q _17780_/A1 _17657_/S vssd1 vssd1 vccd1 vccd1 _20429_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14855_ _14851_/X _14854_/X _15165_/S vssd1 vssd1 vccd1 vccd1 _14855_/X sky130_fd_sc_hd__mux2_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13806_ _13810_/A1 _13701_/Y _13816_/B1 input221/X vssd1 vssd1 vccd1 vccd1 _13806_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_251_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17574_ _17919_/A _17574_/B _17574_/C vssd1 vssd1 vccd1 vccd1 _17574_/X sky130_fd_sc_hd__and3_4
X_14786_ _19140_/Q _14802_/A2 _14785_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _19517_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_251_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11998_ _12153_/A1 _11997_/X _12153_/B1 vssd1 vssd1 vccd1 vccd1 _11998_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19313_ _20539_/CLK _19313_/D vssd1 vssd1 vccd1 vccd1 _19313_/Q sky130_fd_sc_hd__dfxtp_1
X_16525_ input42/X _16598_/A _18905_/A vssd1 vssd1 vccd1 vccd1 _16525_/X sky130_fd_sc_hd__a21o_1
XFILLER_205_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13737_ _13798_/A1 _13777_/B _13736_/X vssd1 vssd1 vccd1 vccd1 _13738_/B sky130_fd_sc_hd__a21oi_4
X_10949_ _10947_/X _10948_/X _11033_/S vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16456_ _16605_/A _17574_/B _16456_/C vssd1 vssd1 vccd1 vccd1 _16456_/X sky130_fd_sc_hd__and3_4
XFILLER_177_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19244_ _19246_/CLK _19244_/D vssd1 vssd1 vccd1 vccd1 _19244_/Q sky130_fd_sc_hd__dfxtp_4
X_13668_ _13669_/B vssd1 vssd1 vccd1 vccd1 _13668_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15407_ _15049_/X _15064_/X _15407_/S vssd1 vssd1 vccd1 vccd1 _15407_/X sky130_fd_sc_hd__mux2_1
X_19175_ _20665_/CLK _19175_/D vssd1 vssd1 vccd1 vccd1 _19175_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12619_ split8/A _12847_/A2 _12716_/B vssd1 vssd1 vccd1 vccd1 _12744_/B sky130_fd_sc_hd__a21oi_4
X_16387_ _18064_/A _16387_/B _16388_/B vssd1 vssd1 vccd1 vccd1 _19740_/D sky130_fd_sc_hd__nor3_1
X_13599_ _19224_/Q _13587_/B _19225_/Q vssd1 vssd1 vccd1 vccd1 _13599_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18126_ _18126_/A _18126_/B vssd1 vssd1 vccd1 vccd1 _18126_/Y sky130_fd_sc_hd__nor2_1
XFILLER_191_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15338_ _20953_/Q _15568_/A2 _15568_/B1 _20825_/Q _15337_/X vssd1 vssd1 vccd1 vccd1
+ _15338_/X sky130_fd_sc_hd__a221o_4
XFILLER_129_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18057_ _20758_/Q _18055_/B _18056_/Y vssd1 vssd1 vccd1 vccd1 _20758_/D sky130_fd_sc_hd__o21a_1
XFILLER_117_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15269_ _20727_/Q _15445_/A2 _15445_/B1 _20759_/Q vssd1 vssd1 vccd1 vccd1 _15269_/X
+ sky130_fd_sc_hd__a22o_1
X_17008_ _17008_/A1 _17006_/X _17008_/B1 vssd1 vssd1 vccd1 vccd1 _17008_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout507 _17779_/X vssd1 vssd1 vccd1 vccd1 _17794_/S sky130_fd_sc_hd__clkbuf_16
X_09830_ _19820_/Q _10603_/B _09828_/X _12085_/B2 _09829_/X vssd1 vssd1 vccd1 vccd1
+ _09830_/X sky130_fd_sc_hd__o221a_1
Xfanout518 _17706_/S vssd1 vssd1 vccd1 vccd1 _17708_/S sky130_fd_sc_hd__buf_12
XFILLER_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout529 _17574_/X vssd1 vssd1 vccd1 vccd1 _17601_/S sky130_fd_sc_hd__buf_4
XFILLER_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09761_ _09755_/X _09760_/X _12012_/S vssd1 vssd1 vccd1 vccd1 _09761_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18959_ _18550_/X _18964_/B _18957_/X _18958_/Y vssd1 vssd1 vccd1 vccd1 _18960_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_273_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09692_ _19952_/Q _11895_/B vssd1 vssd1 vccd1 vccd1 _09692_/X sky130_fd_sc_hd__or2_1
XFILLER_239_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20921_ _21019_/CLK _20921_/D vssd1 vssd1 vccd1 vccd1 _20921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_255_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20852_ _21016_/CLK _20852_/D vssd1 vssd1 vccd1 vccd1 _20852_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20783_ _20816_/CLK _20783_/D vssd1 vssd1 vccd1 vccd1 _20783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_145_wb_clk_i clkbuf_4_6__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19232_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_278_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20217_ _20261_/CLK _20217_/D vssd1 vssd1 vccd1 vccd1 _20217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20148_ _20180_/CLK _20148_/D vssd1 vssd1 vccd1 vccd1 _20148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_265_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09959_ _19682_/Q _20170_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__mux2_1
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12970_ _19107_/Q _19106_/Q _19104_/Q _19105_/Q vssd1 vssd1 vccd1 vccd1 _12971_/B
+ sky130_fd_sc_hd__or4b_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20079_ _20710_/CLK _20079_/D vssd1 vssd1 vccd1 vccd1 _20079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_218_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _12157_/A1 _17877_/A1 _11920_/X _12153_/B1 vssd1 vssd1 vccd1 vccd1 _11921_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_401 _16811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_412 _18215_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14640_ _19402_/Q _17647_/A1 _14650_/S vssd1 vssd1 vccd1 vccd1 _19402_/D sky130_fd_sc_hd__mux2_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_423 _10379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _19390_/Q _12009_/A2 _11850_/X _11852_/B2 _11851_/X vssd1 vssd1 vccd1 vccd1
+ _11852_/X sky130_fd_sc_hd__o221a_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_434 _13669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_445 _13755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_456 _19105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_467 _19848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10803_ _10799_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10803_/Y sky130_fd_sc_hd__nand2b_2
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _19337_/Q _17923_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19337_/D sky130_fd_sc_hd__mux2_1
XFILLER_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_478 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ _15058_/S _11783_/B vssd1 vssd1 vccd1 vccd1 _14878_/A sky130_fd_sc_hd__or2_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_489 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16310_ _16314_/C _16310_/B vssd1 vssd1 vccd1 vccd1 _19711_/D sky130_fd_sc_hd__nor2_1
XFILLER_199_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13522_ _16241_/A _13911_/A vssd1 vssd1 vccd1 vccd1 _13522_/Y sky130_fd_sc_hd__nor2_2
X_17290_ _17290_/A _17290_/B _17290_/C vssd1 vssd1 vccd1 vccd1 _17290_/X sky130_fd_sc_hd__and3_1
XFILLER_242_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ _09503_/A _10733_/X _10732_/X vssd1 vssd1 vccd1 vccd1 _10734_/X sky130_fd_sc_hd__o21a_1
XFILLER_198_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16241_ _16241_/A _16241_/B vssd1 vssd1 vccd1 vccd1 _19659_/D sky130_fd_sc_hd__nor2_1
XFILLER_158_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13453_ _13453_/A _13453_/B _13453_/C vssd1 vssd1 vccd1 vccd1 _13453_/X sky130_fd_sc_hd__and3_1
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10665_ _12312_/A1 _20500_/Q _12309_/S _10657_/X vssd1 vssd1 vccd1 vccd1 _10665_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ _12517_/B _11726_/S _12403_/Y vssd1 vssd1 vccd1 vccd1 _12436_/A sky130_fd_sc_hd__o21a_1
X_16172_ _19610_/Q _15725_/X _16190_/S vssd1 vssd1 vccd1 vccd1 _16173_/B sky130_fd_sc_hd__mux2_1
X_13384_ _13383_/A _13383_/B _13607_/B vssd1 vssd1 vccd1 vccd1 _13384_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_166_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10596_ _12402_/A1 _17895_/A1 _10595_/X _13657_/A vssd1 vssd1 vccd1 vccd1 _10596_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15123_ _15578_/S _15122_/Y _15548_/B1 vssd1 vssd1 vccd1 vccd1 _15123_/X sky130_fd_sc_hd__a21bo_4
X_12335_ _12333_/X _12334_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _12335_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19931_ _20463_/CLK _19931_/D vssd1 vssd1 vccd1 vccd1 _19931_/Q sky130_fd_sc_hd__dfxtp_1
X_15054_ _14827_/X _14833_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _15054_/X sky130_fd_sc_hd__mux2_1
X_12266_ _12265_/A _12261_/X _12265_/Y _12431_/A1 vssd1 vssd1 vccd1 vccd1 _12275_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14005_ _14035_/A1 _14011_/A2 _10374_/X _14035_/B1 _19850_/Q vssd1 vssd1 vccd1 vccd1
+ _14083_/C sky130_fd_sc_hd__o32a_2
X_11217_ _11375_/S _11212_/X _11216_/X _10260_/S vssd1 vssd1 vccd1 vccd1 _11217_/X
+ sky130_fd_sc_hd__o211a_1
X_19862_ _20014_/CLK _19862_/D vssd1 vssd1 vccd1 vccd1 _19862_/Q sky130_fd_sc_hd__dfxtp_4
X_12197_ _12284_/A _12198_/B vssd1 vssd1 vccd1 vccd1 _12197_/Y sky130_fd_sc_hd__nor2_2
XFILLER_96_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_233_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18813_ _18589_/B _18811_/X _18812_/X vssd1 vssd1 vccd1 vccd1 _18814_/B sky130_fd_sc_hd__a21oi_1
X_11148_ _19592_/Q _11225_/B vssd1 vssd1 vccd1 vccd1 _11148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_268_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19793_ _20580_/CLK _19793_/D vssd1 vssd1 vccd1 vccd1 _19793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_284_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18744_ _18746_/A _18744_/B vssd1 vssd1 vccd1 vccd1 _20972_/D sky130_fd_sc_hd__and2_1
XFILLER_283_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ _11077_/X _11078_/X _12383_/A vssd1 vssd1 vccd1 vccd1 _11079_/X sky130_fd_sc_hd__mux2_1
X_15956_ _12199_/B _12466_/Y _12468_/X _12197_/Y _15365_/A vssd1 vssd1 vccd1 vccd1
+ _15956_/X sky130_fd_sc_hd__o221a_1
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput170 dout1[9] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_hd__clkbuf_2
XFILLER_271_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput181 irq[4] vssd1 vssd1 vccd1 vccd1 _12534_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14907_ _18149_/S _19179_/Q _14906_/X vssd1 vssd1 vccd1 vccd1 _14950_/B sky130_fd_sc_hd__a21o_1
Xinput192 localMemory_wb_adr_i[11] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18675_ _19522_/Q _18683_/B vssd1 vssd1 vccd1 vccd1 _18675_/Y sky130_fd_sc_hd__nand2_1
X_15887_ _15264_/B _15984_/A2 _15887_/S vssd1 vssd1 vccd1 vccd1 _15887_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17626_ _20382_/Q _17903_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20382_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14838_ _14836_/X _14837_/X _15035_/S vssd1 vssd1 vccd1 vccd1 _14838_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17557_ _20317_/Q _17693_/A1 _17569_/S vssd1 vssd1 vccd1 vccd1 _20317_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14769_ _19509_/Q _14773_/B vssd1 vssd1 vccd1 vccd1 _14769_/X sky130_fd_sc_hd__or2_1
XFILLER_205_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16508_ _19815_/Q _17592_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19815_/D sky130_fd_sc_hd__mux2_1
X_17488_ _20279_/Q _17494_/B vssd1 vssd1 vccd1 vccd1 _17488_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19227_ _19505_/CLK _19227_/D vssd1 vssd1 vccd1 vccd1 _19227_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_258_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16439_ _19760_/Q _16442_/C _18835_/A vssd1 vssd1 vccd1 vccd1 _16439_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_176_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19158_ _19577_/CLK _19158_/D vssd1 vssd1 vccd1 vccd1 _19158_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_157_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18109_ _20778_/Q _20777_/Q _18109_/C vssd1 vssd1 vccd1 vccd1 _18111_/B sky130_fd_sc_hd__and3_1
XFILLER_258_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19089_ _20721_/CLK _19089_/D vssd1 vssd1 vccd1 vccd1 _19089_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_219_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20002_ _20004_/CLK _20002_/D vssd1 vssd1 vccd1 vccd1 _20002_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_98_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _20419_/Q _12070_/S _09799_/X _12063_/C1 vssd1 vssd1 vccd1 vccd1 _09813_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09744_ _14668_/B _09744_/B vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__xnor2_1
XFILLER_246_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09675_ _11242_/A1 _14011_/A2 _09672_/C _09673_/X _11229_/S vssd1 vssd1 vccd1 vccd1
+ _09676_/B sky130_fd_sc_hd__o311ai_4
XFILLER_27_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20904_ _21010_/CLK _20904_/D vssd1 vssd1 vccd1 vccd1 _20904_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20835_ _21030_/CLK _20835_/D vssd1 vssd1 vccd1 vccd1 _20835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20766_ _20766_/CLK _20766_/D vssd1 vssd1 vccd1 vccd1 _20766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20697_ _20718_/CLK _20697_/D vssd1 vssd1 vccd1 vccd1 _20697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10450_ _12708_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _10450_/X sky130_fd_sc_hd__or2_1
XFILLER_109_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ _19586_/Q _10380_/X _11229_/S vssd1 vssd1 vccd1 vccd1 _10382_/B sky130_fd_sc_hd__mux2_2
XFILLER_191_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ _12120_/A1 _19490_/Q _19458_/Q _12121_/S _12123_/C1 vssd1 vssd1 vccd1 vccd1
+ _12120_/X sky130_fd_sc_hd__a221o_1
XFILLER_191_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12051_ _12051_/A1 _19488_/Q _19456_/Q _12053_/S _12051_/C1 vssd1 vssd1 vccd1 vccd1
+ _12051_/X sky130_fd_sc_hd__a221o_1
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1803 _16769_/S vssd1 vssd1 vccd1 vccd1 _17009_/S sky130_fd_sc_hd__buf_6
XFILLER_2_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11002_ _19369_/Q _11009_/A2 _11000_/X _11009_/B2 _11001_/X vssd1 vssd1 vccd1 vccd1
+ _11002_/X sky130_fd_sc_hd__o221a_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1814 _19300_/Q vssd1 vssd1 vccd1 vccd1 _14524_/B1 sky130_fd_sc_hd__buf_4
XFILLER_120_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1825 _11670_/S vssd1 vssd1 vccd1 vccd1 _12058_/S sky130_fd_sc_hd__buf_12
XFILLER_278_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1836 _12584_/B vssd1 vssd1 vccd1 vccd1 _11101_/A sky130_fd_sc_hd__buf_12
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1847 _12584_/C vssd1 vssd1 vccd1 vccd1 _12306_/A1 sky130_fd_sc_hd__buf_4
XFILLER_237_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1858 _11118_/A vssd1 vssd1 vccd1 vccd1 _12265_/A sky130_fd_sc_hd__buf_6
Xfanout860 _15337_/A2 vssd1 vssd1 vccd1 vccd1 _15567_/A2 sky130_fd_sc_hd__buf_8
XFILLER_93_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1869 _19166_/Q vssd1 vssd1 vccd1 vccd1 _12015_/A1 sky130_fd_sc_hd__clkbuf_8
X_15810_ _15246_/A _15808_/Y _15809_/Y _13414_/Y _12578_/A vssd1 vssd1 vccd1 vccd1
+ _15810_/X sky130_fd_sc_hd__o32a_1
XFILLER_77_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout871 _15322_/A vssd1 vssd1 vccd1 vccd1 _15937_/A2 sky130_fd_sc_hd__buf_6
XFILLER_120_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16790_ _16790_/A vssd1 vssd1 vccd1 vccd1 _16790_/Y sky130_fd_sc_hd__clkinv_4
Xfanout882 _15999_/C1 vssd1 vssd1 vccd1 vccd1 _15971_/C1 sky130_fd_sc_hd__buf_4
XFILLER_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout893 _18395_/S vssd1 vssd1 vccd1 vccd1 _18449_/S sky130_fd_sc_hd__buf_6
XFILLER_219_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15741_ _15741_/A _15988_/B vssd1 vssd1 vccd1 vccd1 _15741_/X sky130_fd_sc_hd__and2_1
XFILLER_86_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12953_ _20021_/Q _20020_/Q vssd1 vssd1 vccd1 vccd1 _13790_/A sky130_fd_sc_hd__and2b_4
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11904_ _11902_/X _11903_/X _11904_/S vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_261_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20702_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_18460_ _18459_/Y _20882_/Q _18474_/S vssd1 vssd1 vccd1 vccd1 _18460_/X sky130_fd_sc_hd__mux2_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ _16050_/A1 _15671_/X _15659_/X vssd1 vssd1 vccd1 vccd1 _15672_/X sky130_fd_sc_hd__a21o_1
XANTENNA_220 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12884_ _19519_/Q _12884_/B vssd1 vssd1 vccd1 vccd1 _12884_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_242 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14623_ _19387_/Q _17907_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19387_/D sky130_fd_sc_hd__mux2_1
X_17411_ _17402_/Y _17410_/X _17409_/X _17434_/A vssd1 vssd1 vccd1 vccd1 _20252_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _20850_/Q _18160_/Y _18421_/S vssd1 vssd1 vccd1 vccd1 _18392_/B sky130_fd_sc_hd__mux2_1
XANTENNA_253 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11835_ _11988_/S _11834_/X _11833_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _11835_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_264 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_275 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_286 _17236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17342_ _20219_/Q _17364_/A2 _17362_/B1 _20268_/Q _17362_/C1 vssd1 vssd1 vccd1 vccd1
+ _17342_/X sky130_fd_sc_hd__a221o_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_297 input226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _19324_/Q _17874_/A1 _14558_/S vssd1 vssd1 vccd1 vccd1 _19324_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _13611_/A _11766_/B _11773_/A vssd1 vssd1 vccd1 vccd1 _15433_/B sky130_fd_sc_hd__nand3_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13505_/A _13519_/S vssd1 vssd1 vccd1 vccd1 _13505_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17273_ _20196_/Q _17330_/A2 _17279_/C1 vssd1 vssd1 vccd1 vccd1 _17273_/X sky130_fd_sc_hd__a21o_1
X_10717_ _10718_/A _10802_/B vssd1 vssd1 vccd1 vccd1 _10720_/A sky130_fd_sc_hd__and2_4
X_14485_ _17850_/A _17884_/A _09632_/B _16087_/B1 vssd1 vssd1 vccd1 vccd1 _17885_/B
+ sky130_fd_sc_hd__o211a_1
X_11697_ _12102_/A1 _20383_/Q _20447_/Q _11698_/B2 vssd1 vssd1 vccd1 vccd1 _11697_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ _19647_/Q _17876_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19647_/D sky130_fd_sc_hd__mux2_1
X_19012_ _18225_/Y _18982_/B _19016_/B1 _19011_/X vssd1 vssd1 vccd1 vccd1 _21025_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_228_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13436_ _15954_/A _13436_/B _15949_/B _15981_/A vssd1 vssd1 vccd1 vccd1 _13437_/B
+ sky130_fd_sc_hd__or4b_1
X_10648_ _09503_/A _10647_/X _10646_/X vssd1 vssd1 vccd1 vccd1 _10648_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_42_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16155_ _19601_/Q _16178_/S _16154_/Y _16159_/C1 vssd1 vssd1 vccd1 vccd1 _19601_/D
+ sky130_fd_sc_hd__o211a_1
X_13367_ _13025_/Y _13367_/B vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__nand2b_1
X_10579_ _11670_/S _10574_/X _10578_/X _12059_/C1 vssd1 vssd1 vccd1 vccd1 _10579_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15106_ _14813_/X _14823_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15106_/X sky130_fd_sc_hd__mux2_1
X_12318_ _12318_/A1 _12317_/X _12314_/X _11275_/A vssd1 vssd1 vccd1 vccd1 _12318_/X
+ sky130_fd_sc_hd__o211a_2
X_16086_ _11232_/X _16106_/A2 _16085_/X vssd1 vssd1 vccd1 vccd1 _19567_/D sky130_fd_sc_hd__o21a_1
XFILLER_138_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _14110_/B _13365_/B _13296_/Y _13297_/Y vssd1 vssd1 vccd1 vccd1 _13298_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15037_ _15035_/X _15036_/X _15155_/S vssd1 vssd1 vccd1 vccd1 _15037_/X sky130_fd_sc_hd__mux2_1
X_19914_ _20681_/CLK _19914_/D vssd1 vssd1 vccd1 vccd1 _19914_/Q sky130_fd_sc_hd__dfxtp_1
X_12249_ _12337_/A _19331_/Q _12337_/C vssd1 vssd1 vccd1 vccd1 _12249_/X sky130_fd_sc_hd__or3_1
XFILLER_142_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_257_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_284_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19845_ _20014_/CLK _19845_/D vssd1 vssd1 vccd1 vccd1 _19845_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19776_ _21047_/A _19776_/D vssd1 vssd1 vccd1 vccd1 _19776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16988_ _20426_/Q _17004_/A2 _17004_/B1 vssd1 vssd1 vccd1 vccd1 _16988_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18727_ _20964_/Q _18250_/Y _18749_/S vssd1 vssd1 vccd1 vccd1 _18728_/B sky130_fd_sc_hd__mux2_1
XFILLER_243_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15939_ _20973_/Q _15939_/A2 _16016_/S _20845_/Q _15938_/X vssd1 vssd1 vccd1 vccd1
+ _15939_/X sky130_fd_sc_hd__a221o_1
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_264_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18658_ _20938_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18658_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_280_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17609_ _20365_/Q _17780_/A1 _17623_/S vssd1 vssd1 vccd1 vccd1 _20365_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18589_ _19500_/Q _18589_/B vssd1 vssd1 vccd1 vccd1 _18589_/Y sky130_fd_sc_hd__nand2_2
XFILLER_240_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20620_ _20663_/CLK _20620_/D vssd1 vssd1 vccd1 vccd1 _20620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20551_ _20683_/CLK _20551_/D vssd1 vssd1 vccd1 vccd1 _20551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20482_ _20482_/CLK _20482_/D vssd1 vssd1 vccd1 vccd1 _20482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_180_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput430 _19989_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[28] sky130_fd_sc_hd__buf_4
XFILLER_191_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput441 _19970_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[9] sky130_fd_sc_hd__buf_4
Xoutput452 _19505_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[11] sky130_fd_sc_hd__buf_4
XFILLER_105_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput463 _19515_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[21] sky130_fd_sc_hd__buf_4
Xoutput474 _19525_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[31] sky130_fd_sc_hd__buf_4
XFILLER_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput485 _13824_/X vssd1 vssd1 vccd1 vccd1 wmask0[1] sky130_fd_sc_hd__buf_6
XFILLER_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21034_ _21042_/CLK _21034_/D vssd1 vssd1 vccd1 vccd1 _21034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09727_ _12513_/D _11649_/S _09726_/Y vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__o21a_1
XFILLER_262_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09658_ _10373_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _11326_/A sky130_fd_sc_hd__nor2_8
XFILLER_216_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_271_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09589_ _19098_/Q _12967_/B _09610_/A vssd1 vssd1 vccd1 vccd1 _09589_/X sky130_fd_sc_hd__o21a_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _12007_/A1 _20384_/Q _20448_/Q _12013_/S vssd1 vssd1 vccd1 vccd1 _11620_/X
+ sky130_fd_sc_hd__a22o_1
X_20818_ _20818_/CLK _20818_/D vssd1 vssd1 vccd1 vccd1 _20818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _12191_/C1 _11945_/S _11548_/X _11550_/X vssd1 vssd1 vccd1 vccd1 _11551_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_196_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20749_ _20812_/CLK _20749_/D vssd1 vssd1 vccd1 vccd1 _20749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ _19808_/Q _10502_/A2 _10500_/X _11274_/B2 _10501_/X vssd1 vssd1 vccd1 vccd1
+ _10502_/X sky130_fd_sc_hd__o221a_1
XFILLER_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14270_ _14278_/A _14270_/B vssd1 vssd1 vccd1 vccd1 _14271_/C sky130_fd_sc_hd__or2_1
X_11482_ _11846_/C _11481_/X _11478_/X _09839_/A vssd1 vssd1 vccd1 vccd1 _11482_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_160_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21030_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13221_ _13221_/A _13221_/B _13221_/C vssd1 vssd1 vccd1 vccd1 _13221_/X sky130_fd_sc_hd__or3_1
XFILLER_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10433_ _20636_/Q _12043_/B _12072_/A1 vssd1 vssd1 vccd1 vccd1 _10433_/X sky130_fd_sc_hd__a21o_1
XFILLER_152_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13152_ _11774_/B _13570_/B _15374_/S vssd1 vssd1 vccd1 vccd1 _13596_/B sky130_fd_sc_hd__a21o_4
X_10364_ _10365_/A _11414_/B vssd1 vssd1 vccd1 vccd1 _10366_/A sky130_fd_sc_hd__or2_4
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ _12103_/A1 _12102_/X _12828_/A vssd1 vssd1 vccd1 vccd1 _12103_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17960_ _20724_/Q _17962_/C _17963_/B1 vssd1 vssd1 vccd1 vccd1 _17961_/B sky130_fd_sc_hd__o21ai_1
X_13083_ _13258_/A _13258_/C _13258_/B vssd1 vssd1 vccd1 vccd1 _13195_/A sky130_fd_sc_hd__a21boi_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10295_ _20475_/Q _20315_/Q _11255_/S vssd1 vssd1 vccd1 vccd1 _10295_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16911_ _16908_/Y _16910_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16911_/Y sky130_fd_sc_hd__a21oi_4
Xfanout1600 _11833_/C1 vssd1 vssd1 vccd1 vccd1 _09901_/S sky130_fd_sc_hd__buf_6
X_12034_ _12035_/A _12035_/B vssd1 vssd1 vccd1 vccd1 _12034_/Y sky130_fd_sc_hd__nor2_1
Xfanout1611 _11513_/S vssd1 vssd1 vccd1 vccd1 _11902_/S sky130_fd_sc_hd__buf_6
XFILLER_278_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17891_ _20662_/Q _17891_/A1 _17916_/S vssd1 vssd1 vccd1 vccd1 _20662_/D sky130_fd_sc_hd__mux2_1
Xfanout1622 _10152_/S vssd1 vssd1 vccd1 vccd1 _10322_/S sky130_fd_sc_hd__buf_6
XFILLER_239_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1633 _09615_/Y vssd1 vssd1 vccd1 vccd1 _12311_/C1 sky130_fd_sc_hd__buf_12
XFILLER_104_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1644 _18949_/A2 vssd1 vssd1 vccd1 vccd1 _18976_/A2 sky130_fd_sc_hd__buf_6
X_19630_ _20061_/CLK _19630_/D vssd1 vssd1 vccd1 vccd1 _19630_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1655 _09655_/Y vssd1 vssd1 vccd1 vccd1 _13960_/A2 sky130_fd_sc_hd__buf_12
XFILLER_144_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16842_ _16878_/A _16842_/B vssd1 vssd1 vccd1 vccd1 _16842_/Y sky130_fd_sc_hd__nand2_1
XFILLER_265_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1666 _09533_/Y vssd1 vssd1 vccd1 vccd1 _12464_/C sky130_fd_sc_hd__buf_12
XFILLER_265_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1677 _11946_/A1 vssd1 vssd1 vccd1 vccd1 _09986_/A sky130_fd_sc_hd__buf_6
XFILLER_266_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1688 _11191_/A vssd1 vssd1 vccd1 vccd1 _12711_/A sky130_fd_sc_hd__buf_12
Xfanout690 _13805_/B1 vssd1 vssd1 vccd1 vccd1 _13826_/B1 sky130_fd_sc_hd__buf_8
Xfanout1699 _12337_/A vssd1 vssd1 vccd1 vccd1 _12332_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19561_ _19621_/CLK _19561_/D vssd1 vssd1 vccd1 vccd1 _19561_/Q sky130_fd_sc_hd__dfxtp_1
X_13985_ _19194_/Q _14069_/C _14003_/S vssd1 vssd1 vccd1 vccd1 _13985_/X sky130_fd_sc_hd__mux2_1
X_16773_ _19965_/Q _16849_/A _16772_/Y _16451_/A vssd1 vssd1 vccd1 vccd1 _19965_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_168_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18512_ _20897_/Q _18559_/B _18511_/X _18458_/B vssd1 vssd1 vccd1 vccd1 _18513_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12936_ _19260_/Q _12950_/B2 _12930_/X _20008_/Q vssd1 vssd1 vccd1 vccd1 _12945_/A
+ sky130_fd_sc_hd__a22o_4
X_15724_ _19753_/Q _15999_/A2 _15723_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15724_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ _20719_/CLK _19492_/D vssd1 vssd1 vccd1 vccd1 _19492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ _20876_/Q _18290_/Y _18449_/S vssd1 vssd1 vccd1 vccd1 _18444_/B sky130_fd_sc_hd__mux2_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12867_ _12803_/B _12815_/B _12906_/A vssd1 vssd1 vccd1 vccd1 _13389_/B sky130_fd_sc_hd__o21a_2
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15655_ _11496_/Y _16058_/A2 _15264_/B _13420_/A _15890_/A vssd1 vssd1 vccd1 vccd1
+ _15655_/X sky130_fd_sc_hd__a221o_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _19370_/Q _17890_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19370_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11818_ _12120_/A1 _19486_/Q _19454_/Q _11818_/B2 _11892_/C1 vssd1 vssd1 vccd1 vccd1
+ _11818_/X sky130_fd_sc_hd__a221o_1
X_18374_ _20842_/Q _18385_/B _18373_/Y _18734_/A vssd1 vssd1 vccd1 vccd1 _20842_/D
+ sky130_fd_sc_hd__o211a_1
X_15586_ _15582_/Y _15583_/Y _15585_/X vssd1 vssd1 vccd1 vccd1 _15586_/Y sky130_fd_sc_hd__a21oi_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _12750_/Y _13279_/A _12794_/X _12793_/Y vssd1 vssd1 vccd1 vccd1 _13346_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_187_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _19307_/Q _17751_/A1 _14562_/S vssd1 vssd1 vccd1 vccd1 _19307_/D sky130_fd_sc_hd__mux2_1
X_17325_ _20214_/Q _17232_/X _17324_/X _17974_/B1 vssd1 vssd1 vccd1 vccd1 _20214_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11749_ _11791_/A _11791_/B _13421_/A vssd1 vssd1 vccd1 vccd1 _11794_/C sky130_fd_sc_hd__a21o_1
XFILLER_105_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17256_ _20191_/Q _17268_/A2 _17254_/X _17255_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1
+ _20191_/D sky130_fd_sc_hd__o221a_1
X_14468_ _18700_/A _14468_/B vssd1 vssd1 vccd1 vccd1 _19258_/D sky130_fd_sc_hd__and2_1
X_16207_ _19630_/Q _17859_/A1 _16230_/S vssd1 vssd1 vccd1 vccd1 _19630_/D sky130_fd_sc_hd__mux2_1
X_13419_ _13419_/A _13419_/B vssd1 vssd1 vccd1 vccd1 _13427_/A sky130_fd_sc_hd__xor2_4
X_17187_ _20151_/Q _17921_/A1 _17217_/S vssd1 vssd1 vccd1 vccd1 _20151_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14399_ _20294_/Q _14431_/A2 _14431_/B1 input235/X vssd1 vssd1 vccd1 vccd1 _14406_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16138_ _16743_/B _16164_/B vssd1 vssd1 vccd1 vccd1 _16138_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16069_ _19559_/Q _16081_/B _16087_/B1 vssd1 vssd1 vccd1 vccd1 _16069_/X sky130_fd_sc_hd__o21a_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_269_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19828_ _20084_/CLK _19828_/D vssd1 vssd1 vccd1 vccd1 _19828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_257_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_284_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19759_ _19759_/CLK _19759_/D vssd1 vssd1 vccd1 vccd1 _19759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09512_ _19090_/Q vssd1 vssd1 vccd1 vccd1 _09585_/A sky130_fd_sc_hd__inv_2
XFILLER_271_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_262_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20603_ _20635_/CLK _20603_/D vssd1 vssd1 vccd1 vccd1 _20603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20534_ _20675_/CLK _20534_/D vssd1 vssd1 vccd1 vccd1 _20534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20465_ _20465_/CLK _20465_/D vssd1 vssd1 vccd1 vccd1 _20465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20396_ _20687_/CLK _20396_/D vssd1 vssd1 vccd1 vccd1 _20396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput293 _13835_/X vssd1 vssd1 vccd1 vccd1 addr0[8] sky130_fd_sc_hd__buf_4
X_10080_ _19778_/Q _11708_/B _12100_/B1 vssd1 vssd1 vccd1 vccd1 _10080_/X sky130_fd_sc_hd__o21a_1
XFILLER_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21017_ _21017_/CLK _21017_/D vssd1 vssd1 vccd1 vccd1 _21017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13770_ _13780_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13770_/X sky130_fd_sc_hd__and2_1
XFILLER_261_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ _10979_/X _10980_/X _10981_/X _11250_/S _12377_/S vssd1 vssd1 vccd1 vccd1
+ _10982_/X sky130_fd_sc_hd__o221a_1
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12721_ _12719_/X _12720_/Y _12716_/B vssd1 vssd1 vccd1 vccd1 _12721_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ _14837_/S _15438_/Y _15439_/Y _15437_/Y vssd1 vssd1 vccd1 vccd1 _15440_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_230_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12652_ _19175_/Q _12652_/B vssd1 vssd1 vccd1 vccd1 _12653_/C sky130_fd_sc_hd__and2_1
XFILLER_71_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _11980_/S _11602_/X _11601_/X _12144_/A1 vssd1 vssd1 vccd1 vccd1 _11603_/X
+ sky130_fd_sc_hd__a211o_1
X_15371_ _14825_/X _14856_/X _15577_/S vssd1 vssd1 vccd1 vccd1 _15372_/A sky130_fd_sc_hd__mux2_1
XFILLER_212_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12583_ _12978_/A _12583_/B _12583_/C _14809_/A vssd1 vssd1 vccd1 vccd1 _12583_/Y
+ sky130_fd_sc_hd__nor4b_2
XFILLER_230_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14322_ _19514_/Q _14322_/B vssd1 vssd1 vccd1 vccd1 _14323_/C sky130_fd_sc_hd__xnor2_1
XFILLER_90_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17110_ _20080_/Q _17878_/A1 _17111_/S vssd1 vssd1 vccd1 vccd1 _20080_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18090_ _20771_/Q _18093_/C _18094_/A vssd1 vssd1 vccd1 vccd1 _18090_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_196_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11534_ _10561_/A _11532_/X _11533_/X vssd1 vssd1 vccd1 vccd1 _11534_/X sky130_fd_sc_hd__a21o_4
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17041_ _18048_/A _17041_/B vssd1 vssd1 vccd1 vccd1 _20019_/D sky130_fd_sc_hd__nor2_1
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253_ _14262_/A _14249_/B _14252_/X vssd1 vssd1 vccd1 vccd1 _14253_/X sky130_fd_sc_hd__a21bo_1
XFILLER_184_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11465_ _12011_/S _11462_/X _11464_/X _11852_/B2 vssd1 vssd1 vccd1 vccd1 _11465_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13204_ _18683_/B _13196_/X _13197_/Y _13200_/Y _13203_/X vssd1 vssd1 vccd1 vccd1
+ _13205_/B sky130_fd_sc_hd__a32o_1
XFILLER_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10416_ _10395_/X _10403_/X _10409_/X _10415_/X vssd1 vssd1 vccd1 vccd1 _10416_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14184_ _14184_/A _14204_/A _16068_/B vssd1 vssd1 vccd1 vccd1 _14184_/X sky130_fd_sc_hd__or3_1
X_11396_ _11384_/X _11395_/X _11396_/S vssd1 vssd1 vccd1 vccd1 _11396_/X sky130_fd_sc_hd__mux2_4
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13135_ _13135_/A _13135_/B vssd1 vssd1 vccd1 vccd1 _13135_/Y sky130_fd_sc_hd__nor2_1
X_10347_ _10343_/X _10346_/X _10516_/S vssd1 vssd1 vccd1 vccd1 _10347_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18992_ _18175_/Y _18983_/B _19002_/B1 _18991_/X vssd1 vssd1 vccd1 vccd1 _21015_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _20953_/Q _20887_/Q _13563_/A vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__a21o_2
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _20712_/Q _17943_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20712_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10278_ _15613_/S _10278_/B vssd1 vssd1 vccd1 vccd1 _13422_/A sky130_fd_sc_hd__nand2_8
XFILLER_105_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_266_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1430 _09736_/Y vssd1 vssd1 vccd1 vccd1 fanout1430/X sky130_fd_sc_hd__buf_6
X_12017_ _20488_/Q _11708_/B _12103_/A1 vssd1 vssd1 vccd1 vccd1 _12017_/X sky130_fd_sc_hd__a21o_1
XFILLER_78_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1441 _09735_/Y vssd1 vssd1 vccd1 vccd1 _12412_/B2 sky130_fd_sc_hd__buf_12
Xfanout1452 _11021_/C vssd1 vssd1 vccd1 vccd1 _11026_/C sky130_fd_sc_hd__buf_4
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17874_ _20647_/Q _17874_/A1 _17878_/S vssd1 vssd1 vccd1 vccd1 _20647_/D sky130_fd_sc_hd__mux2_1
Xfanout1463 _09733_/Y vssd1 vssd1 vccd1 vccd1 _12415_/S sky130_fd_sc_hd__buf_6
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1474 _12414_/S vssd1 vssd1 vccd1 vccd1 _12345_/S sky130_fd_sc_hd__clkbuf_16
X_19613_ _19620_/CLK _19613_/D vssd1 vssd1 vccd1 vccd1 _19613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16825_ _20407_/Q _17004_/A2 _17004_/B1 vssd1 vssd1 vccd1 vccd1 _16825_/X sky130_fd_sc_hd__a21o_1
Xfanout1485 _12105_/A vssd1 vssd1 vccd1 vccd1 _12191_/C1 sky130_fd_sc_hd__buf_4
XFILLER_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1496 _12043_/B vssd1 vssd1 vccd1 vccd1 _12044_/B sky130_fd_sc_hd__buf_6
XFILLER_253_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19544_ _19609_/CLK _19544_/D vssd1 vssd1 vccd1 vccd1 _19544_/Q sky130_fd_sc_hd__dfxtp_1
X_16756_ _19087_/Q _16996_/B1 _16755_/X vssd1 vssd1 vccd1 vccd1 _16756_/X sky130_fd_sc_hd__o21a_1
X_13968_ _19156_/Q _19050_/S _14043_/B1 _13967_/X _16097_/B1 vssd1 vssd1 vccd1 vccd1
+ _19156_/D sky130_fd_sc_hd__o221a_1
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15707_ _13428_/C _15925_/B _16056_/B1 vssd1 vssd1 vccd1 vccd1 _15707_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_250_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19475_ _20570_/CLK _19475_/D vssd1 vssd1 vccd1 vccd1 _19475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ _12912_/A _12913_/X _12917_/Y _13107_/A vssd1 vssd1 vccd1 vccd1 _12919_/X
+ sky130_fd_sc_hd__a31o_1
X_16687_ _19942_/Q _17097_/A1 _16704_/S vssd1 vssd1 vccd1 vccd1 _19942_/D sky130_fd_sc_hd__mux2_1
X_13899_ _18048_/A _19050_/S vssd1 vssd1 vccd1 vccd1 _14522_/A sky130_fd_sc_hd__or2_4
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18426_ _18728_/A _18426_/B vssd1 vssd1 vccd1 vccd1 _20867_/D sky130_fd_sc_hd__and2_1
XFILLER_221_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15638_ _20962_/Q _15939_/A2 _15996_/B1 _20834_/Q _15637_/X vssd1 vssd1 vccd1 vccd1
+ _15638_/X sky130_fd_sc_hd__a221o_1
XFILLER_222_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18357_ _18514_/B _18357_/B vssd1 vssd1 vccd1 vccd1 _18357_/Y sky130_fd_sc_hd__nand2_1
X_15569_ _20864_/Q _15568_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15569_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17308_ input1/X input267/X _17329_/S vssd1 vssd1 vccd1 vccd1 _17308_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18288_ _19553_/Q _18308_/B vssd1 vssd1 vccd1 vccd1 _18288_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_30_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17239_ _17239_/A _17320_/S _17302_/C vssd1 vssd1 vccd1 vccd1 _17239_/X sky130_fd_sc_hd__and3_1
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20250_ _20261_/CLK _20250_/D vssd1 vssd1 vccd1 vccd1 _20250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20181_ _20181_/CLK _20181_/D vssd1 vssd1 vccd1 vccd1 _20181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09992_ _19386_/Q _12009_/A2 _09990_/X _12183_/C1 _09991_/X vssd1 vssd1 vccd1 vccd1
+ _09992_/X sky130_fd_sc_hd__o221a_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_272_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_272_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_241_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20517_ _20685_/CLK _20517_/D vssd1 vssd1 vccd1 vccd1 _20517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11250_ _11248_/X _11249_/X _11250_/S vssd1 vssd1 vccd1 vccd1 _11250_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20448_ _20480_/CLK _20448_/D vssd1 vssd1 vccd1 vccd1 _20448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10201_ _11326_/B _10201_/B vssd1 vssd1 vccd1 vccd1 _10201_/X sky130_fd_sc_hd__and2_1
XFILLER_162_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11181_ _12513_/C _11173_/X _11180_/X _12400_/A1 vssd1 vssd1 vccd1 vccd1 _11181_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20379_ _20379_/CLK _20379_/D vssd1 vssd1 vccd1 vccd1 _20379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_279_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10132_ _20131_/Q _20099_/Q _12375_/S vssd1 vssd1 vccd1 vccd1 _10132_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14940_ _14945_/A _14983_/A vssd1 vssd1 vccd1 vccd1 _16039_/B sky130_fd_sc_hd__or2_4
X_10063_ _12060_/A1 _20505_/Q _10425_/S _20537_/Q vssd1 vssd1 vccd1 vccd1 _10063_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_282_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ _14869_/X _14870_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__mux2_1
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16610_ _19869_/Q _17647_/A1 _16620_/S vssd1 vssd1 vccd1 vccd1 _19869_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13822_ _13822_/A1 _13780_/B split9/X input239/X vssd1 vssd1 vccd1 vccd1 _13822_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17590_ _20348_/Q _17901_/A1 _17590_/S vssd1 vssd1 vccd1 vccd1 _20348_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16541_ _16551_/A _16541_/B vssd1 vssd1 vccd1 vccd1 _19836_/D sky130_fd_sc_hd__or2_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13753_ _13675_/Y _13741_/B _13741_/Y _13676_/Y _13752_/X vssd1 vssd1 vccd1 vccd1
+ _13754_/B sky130_fd_sc_hd__o221a_4
X_10965_ _12277_/A1 _10894_/X _10964_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _12682_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_250_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ split8/A _12847_/A2 _15526_/A _12703_/X vssd1 vssd1 vccd1 vccd1 _12704_/X
+ sky130_fd_sc_hd__a211o_1
X_19260_ _20621_/CLK _19260_/D vssd1 vssd1 vccd1 vccd1 _19260_/Q sky130_fd_sc_hd__dfxtp_2
X_16472_ _19781_/Q _17935_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19781_/D sky130_fd_sc_hd__mux2_1
XFILLER_189_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13684_ _13684_/A _13684_/B vssd1 vssd1 vccd1 vccd1 _13684_/Y sky130_fd_sc_hd__nand2_4
XFILLER_206_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10896_ _20629_/Q _10897_/A3 _09688_/A vssd1 vssd1 vccd1 vccd1 _10896_/X sky130_fd_sc_hd__a21o_1
XFILLER_231_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18211_ _20796_/Q _18210_/Y _18311_/S vssd1 vssd1 vccd1 vccd1 _18212_/B sky130_fd_sc_hd__mux2_1
XFILLER_93_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15423_ _19743_/Q _15453_/A2 _15415_/X _15606_/A1 _15422_/X vssd1 vssd1 vccd1 vccd1
+ _15423_/X sky130_fd_sc_hd__a221o_1
XFILLER_231_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12635_ _12633_/Y _12634_/Y _12519_/A _13589_/A1 vssd1 vssd1 vccd1 vccd1 _12698_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19191_ _19560_/CLK _19191_/D vssd1 vssd1 vccd1 vccd1 _19191_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18142_ _18149_/S _19113_/Q _14906_/X vssd1 vssd1 vccd1 vccd1 _18144_/A sky130_fd_sc_hd__a21o_1
X_15354_ _15354_/A vssd1 vssd1 vccd1 vccd1 _15354_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12566_ _13653_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _13698_/B sky130_fd_sc_hd__nand2_2
XFILLER_12_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11517_ _12120_/A1 _20509_/Q _12134_/S _11499_/X vssd1 vssd1 vccd1 vccd1 _11517_/X
+ sky130_fd_sc_hd__o211a_1
X_14305_ _14300_/B _14304_/Y _14417_/S vssd1 vssd1 vccd1 vccd1 _14305_/X sky130_fd_sc_hd__mux2_1
X_18073_ _20764_/Q _18071_/B _18072_/Y vssd1 vssd1 vccd1 vccd1 _20764_/D sky130_fd_sc_hd__o21a_1
X_15285_ _15348_/B2 _12647_/X _13539_/B _12578_/A _15284_/X vssd1 vssd1 vccd1 vccd1
+ _15285_/X sky130_fd_sc_hd__o221a_1
X_12497_ _09541_/Y _11312_/X _12738_/B _18765_/A vssd1 vssd1 vccd1 vccd1 _12498_/B
+ sky130_fd_sc_hd__a211o_2
X_17024_ _20002_/Q input211/X _17026_/S vssd1 vssd1 vccd1 vccd1 _20002_/D sky130_fd_sc_hd__mux2_1
X_14236_ _19226_/Q _14256_/A2 _14235_/X _18352_/C1 vssd1 vssd1 vccd1 vccd1 _19226_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_236_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11448_ _11446_/X _11447_/X _12150_/S vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ _20271_/Q _14237_/A2 _14216_/B1 input242/X vssd1 vssd1 vccd1 vccd1 _14171_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ _20309_/Q _11379_/B vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__or2_1
XFILLER_124_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13118_ _20942_/Q _13363_/B _18667_/B vssd1 vssd1 vccd1 vccd1 _13118_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14098_ _19208_/Q _14104_/A2 _14097_/X _16131_/B1 vssd1 vssd1 vccd1 vccd1 _19208_/D
+ sky130_fd_sc_hd__o211a_1
X_18975_ _18975_/A _18975_/B vssd1 vssd1 vccd1 vccd1 _18975_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17926_ _20695_/Q _17926_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20695_/D sky130_fd_sc_hd__mux2_1
X_13049_ _20953_/Q _20887_/Q vssd1 vssd1 vccd1 vccd1 _13049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_267_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_282_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1260 _12730_/A2 vssd1 vssd1 vccd1 vccd1 _12582_/C sky130_fd_sc_hd__clkbuf_8
Xfanout1271 _09594_/X vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__buf_6
XFILLER_78_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17857_ _20630_/Q _17857_/A1 _17882_/S vssd1 vssd1 vccd1 vccd1 _20630_/D sky130_fd_sc_hd__mux2_1
Xfanout1282 _09547_/X vssd1 vssd1 vccd1 vccd1 _11398_/S sky130_fd_sc_hd__buf_6
XFILLER_239_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1293 _12708_/B vssd1 vssd1 vccd1 vccd1 _16062_/B2 sky130_fd_sc_hd__clkbuf_2
XFILLER_227_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16808_ _16804_/Y _16805_/X _16807_/X _17008_/A1 vssd1 vssd1 vccd1 vccd1 _16808_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17788_ _20565_/Q _17788_/A1 _17794_/S vssd1 vssd1 vccd1 vccd1 _20565_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19527_ _19603_/CLK _19527_/D vssd1 vssd1 vccd1 vccd1 _19527_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16739_ _16799_/S _09519_/Y _16726_/X _16738_/Y vssd1 vssd1 vccd1 vccd1 _16739_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_234_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19458_ _20677_/CLK _19458_/D vssd1 vssd1 vccd1 vccd1 _19458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18409_ _20859_/Q _18205_/Y _18419_/S vssd1 vssd1 vccd1 vccd1 _18410_/B sky130_fd_sc_hd__mux2_1
XFILLER_201_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _20574_/CLK _19389_/D vssd1 vssd1 vccd1 vccd1 _19389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20302_ _20694_/CLK _20302_/D vssd1 vssd1 vccd1 vccd1 _20302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20233_ _21024_/CLK _20233_/D vssd1 vssd1 vccd1 vccd1 _20233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_249_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20164_ _20315_/CLK _20164_/D vssd1 vssd1 vccd1 vccd1 _20164_/Q sky130_fd_sc_hd__dfxtp_1
X_09975_ _12134_/S _09974_/X _09973_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _09975_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20095_ _20438_/CLK _20095_/D vssd1 vssd1 vccd1 vccd1 _20095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_264_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_257_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_273_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_242_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_605 _20621_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_616 _13775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_627 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_638 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_649 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20997_ _20998_/CLK _20997_/D vssd1 vssd1 vccd1 vccd1 _20997_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10750_ _20403_/Q _20339_/Q _11161_/S vssd1 vssd1 vccd1 vccd1 _10750_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ _10127_/A _09678_/X _10680_/X vssd1 vssd1 vccd1 vccd1 _10681_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _20491_/Q _11379_/B _12420_/B1 vssd1 vssd1 vccd1 vccd1 _12420_/X sky130_fd_sc_hd__a21o_1
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ _12332_/A _19493_/Q _19461_/Q _12352_/S _11212_/S vssd1 vssd1 vccd1 vccd1
+ _12351_/X sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_67_wb_clk_i clkbuf_leaf_74_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20686_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_194_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ _10262_/A _19462_/Q _19430_/Q _11303_/S vssd1 vssd1 vccd1 vccd1 _11302_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15070_ _15066_/S _15069_/X _15548_/B1 vssd1 vssd1 vccd1 vccd1 _16025_/B sky130_fd_sc_hd__o21ai_4
X_12282_ _12282_/A _12282_/B vssd1 vssd1 vccd1 vccd1 _12283_/B sky130_fd_sc_hd__and2_4
XFILLER_181_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14021_ _19206_/Q _14093_/C _14036_/S vssd1 vssd1 vccd1 vccd1 _14021_/X sky130_fd_sc_hd__mux2_1
X_11233_ _19567_/Q _11232_/X _11240_/S vssd1 vssd1 vccd1 vccd1 _11233_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ _12241_/S _11159_/X _11160_/X _11163_/X _11275_/A vssd1 vssd1 vccd1 vccd1
+ _11164_/X sky130_fd_sc_hd__o311a_2
XFILLER_96_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10115_ input111/X input146/X _11241_/S vssd1 vssd1 vccd1 vccd1 _10115_/X sky130_fd_sc_hd__mux2_8
XFILLER_122_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18760_ _20978_/Q _18760_/B vssd1 vssd1 vccd1 vccd1 _18760_/X sky130_fd_sc_hd__and2_4
XFILLER_95_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xsplit4 split4/A vssd1 vssd1 vccd1 vccd1 split4/X sky130_fd_sc_hd__buf_2
X_11095_ _12398_/C1 _11094_/X _11091_/X _12399_/C1 vssd1 vssd1 vccd1 vccd1 _11095_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ _16000_/A1 _15961_/X _15962_/X _15971_/X vssd1 vssd1 vccd1 vccd1 _15972_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17711_ _17745_/A _17851_/B _17711_/C vssd1 vssd1 vccd1 vccd1 _17711_/X sky130_fd_sc_hd__and3_4
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ _14980_/B _14973_/B vssd1 vssd1 vccd1 vccd1 _14945_/A sky130_fd_sc_hd__or2_4
X_10046_ _20130_/Q _20098_/Q _10425_/S vssd1 vssd1 vccd1 vccd1 _10046_/X sky130_fd_sc_hd__mux2_1
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18691_ _20946_/Q _18160_/Y _18707_/S vssd1 vssd1 vccd1 vccd1 _18692_/B sky130_fd_sc_hd__mux2_1
XFILLER_282_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17642_ _17745_/A _17676_/B _17642_/C vssd1 vssd1 vccd1 vccd1 _17642_/X sky130_fd_sc_hd__and3_4
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14854_ _14852_/X _14853_/X _15058_/S vssd1 vssd1 vccd1 vccd1 _14854_/X sky130_fd_sc_hd__mux2_1
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13805_ _13810_/A1 _13696_/Y _13805_/B1 input220/X vssd1 vssd1 vccd1 vccd1 _13805_/X
+ sky130_fd_sc_hd__a22o_1
X_17573_ _17884_/A _17812_/A vssd1 vssd1 vccd1 vccd1 _17574_/C sky130_fd_sc_hd__nor2_1
X_14785_ _19517_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14785_/X sky130_fd_sc_hd__or2_1
X_11997_ _12152_/A1 _11989_/X _11996_/X _11982_/X vssd1 vssd1 vccd1 vccd1 _11997_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_223_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19312_ _20657_/CLK _19312_/D vssd1 vssd1 vccd1 vccd1 _19312_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16524_ _16594_/B _16594_/C _19830_/Q vssd1 vssd1 vccd1 vccd1 _16524_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10948_ _20465_/Q _20305_/Q _11035_/S vssd1 vssd1 vccd1 vccd1 _10948_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13736_ _13659_/A _13698_/X _13735_/Y _13714_/S vssd1 vssd1 vccd1 vccd1 _13736_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_204_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19243_ _19520_/CLK _19243_/D vssd1 vssd1 vccd1 vccd1 _19243_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16455_ _16604_/B _17812_/A vssd1 vssd1 vccd1 vccd1 _16456_/C sky130_fd_sc_hd__nor2_1
X_10879_ _12275_/A _10879_/B vssd1 vssd1 vccd1 vccd1 _10879_/Y sky130_fd_sc_hd__nor2_1
X_13667_ _13718_/A _13665_/Y _13666_/Y _13655_/A vssd1 vssd1 vccd1 vccd1 _13669_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_220_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _15066_/S _15290_/X _15548_/B1 vssd1 vssd1 vccd1 vccd1 _15406_/Y sky130_fd_sc_hd__o21ai_1
X_19174_ _20426_/CLK _19174_/D vssd1 vssd1 vccd1 vccd1 _19174_/Q sky130_fd_sc_hd__dfxtp_1
X_12618_ _12483_/Y _12617_/Y _16009_/A _12486_/B vssd1 vssd1 vccd1 vccd1 _12618_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16386_ _19739_/Q _19740_/Q _16386_/C vssd1 vssd1 vccd1 vccd1 _16388_/B sky130_fd_sc_hd__and3_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13598_ _20924_/Q _13598_/A2 _18604_/B vssd1 vssd1 vccd1 vccd1 _13598_/Y sky130_fd_sc_hd__a21oi_1
X_18125_ _20784_/Q _18125_/B vssd1 vssd1 vccd1 vccd1 _18126_/B sky130_fd_sc_hd__and2_1
X_15337_ _20921_/Q _15337_/A2 _15336_/X vssd1 vssd1 vccd1 vccd1 _15337_/X sky130_fd_sc_hd__o21a_1
X_12549_ _20869_/Q _12549_/B _12549_/C vssd1 vssd1 vccd1 vccd1 _12553_/D sky130_fd_sc_hd__and3_1
XFILLER_129_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18056_ _18056_/A _18061_/C vssd1 vssd1 vccd1 vccd1 _18056_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_1 _19656_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15268_ _19707_/Q _15475_/A2 _15475_/B1 _19739_/Q vssd1 vssd1 vccd1 vccd1 _15268_/X
+ sky130_fd_sc_hd__a22o_1
X_17007_ _12952_/X _16717_/X _17006_/X vssd1 vssd1 vccd1 vccd1 _17461_/B sky130_fd_sc_hd__a21oi_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14219_ _14219_/A _14219_/B vssd1 vssd1 vccd1 vccd1 _14221_/A sky130_fd_sc_hd__nand2_1
X_15199_ _17281_/A _15482_/A2 _15191_/X _15198_/X vssd1 vssd1 vccd1 vccd1 _15199_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout508 _17745_/X vssd1 vssd1 vccd1 vccd1 _17774_/S sky130_fd_sc_hd__buf_12
Xfanout519 _17676_/X vssd1 vssd1 vccd1 vccd1 _17706_/S sky130_fd_sc_hd__buf_12
XFILLER_112_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09760_ _09758_/X _09759_/X _11933_/S vssd1 vssd1 vccd1 vccd1 _09760_/X sky130_fd_sc_hd__mux2_1
X_18958_ _21008_/Q _18964_/B vssd1 vssd1 vccd1 vccd1 _18958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17909_ _20680_/Q _17909_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20680_/D sky130_fd_sc_hd__mux2_1
XFILLER_255_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09691_ _20548_/Q _11915_/S vssd1 vssd1 vccd1 vccd1 _09691_/X sky130_fd_sc_hd__or2_1
XFILLER_66_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18889_ _20998_/Q _18978_/B vssd1 vssd1 vccd1 vccd1 _18889_/Y sky130_fd_sc_hd__nand2_1
XFILLER_187_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1090 _17951_/A1 vssd1 vssd1 vccd1 vccd1 _17917_/A1 sky130_fd_sc_hd__buf_6
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_266_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20920_ _21013_/CLK _20920_/D vssd1 vssd1 vccd1 vccd1 _20920_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20851_ _20861_/CLK _20851_/D vssd1 vssd1 vccd1 vccd1 _20851_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20782_ _20816_/CLK _20782_/D vssd1 vssd1 vccd1 vccd1 _20782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20216_ _20759_/CLK _20216_/D vssd1 vssd1 vccd1 vccd1 _20216_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_235_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20147_ _20179_/CLK _20147_/D vssd1 vssd1 vccd1 vccd1 _20147_/Q sky130_fd_sc_hd__dfxtp_1
X_09958_ _12120_/A1 _19482_/Q _19450_/Q _11889_/S _11892_/C1 vssd1 vssd1 vccd1 vccd1
+ _09958_/X sky130_fd_sc_hd__a221o_1
XFILLER_77_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_249_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_185_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20425_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20078_ _20649_/CLK _20078_/D vssd1 vssd1 vccd1 vccd1 _20078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_114_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21020_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _11981_/C1 _09888_/X _09885_/X _12137_/C1 vssd1 vssd1 vccd1 vccd1 _09889_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_257_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _11905_/X _11919_/X _12153_/A1 vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__a21o_2
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_402 _16811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_413 _18215_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ _11851_/A _20681_/Q _11851_/C vssd1 vssd1 vccd1 vccd1 _11851_/X sky130_fd_sc_hd__or3_1
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_424 _10462_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_435 _13697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_214_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10802_ _10718_/A _10802_/B vssd1 vssd1 vccd1 vccd1 _10802_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_446 _13755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14570_ _19336_/Q _17922_/A1 _14598_/S vssd1 vssd1 vccd1 vccd1 _19336_/D sky130_fd_sc_hd__mux2_1
XANTENNA_457 _19107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_468 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11782_ _15058_/S _11783_/B vssd1 vssd1 vccd1 vccd1 _13694_/A sky130_fd_sc_hd__nand2_8
XANTENNA_479 _19998_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10733_ _19404_/Q _20563_/Q _11074_/S vssd1 vssd1 vccd1 vccd1 _10733_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13521_ _18763_/A1 _19219_/Q _13520_/X vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__a21oi_4
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16240_ _16240_/A1 _16239_/X _19695_/D vssd1 vssd1 vccd1 vccd1 _19658_/D sky130_fd_sc_hd__o21a_2
X_13452_ split6/X _13448_/Y _13451_/X vssd1 vssd1 vccd1 vccd1 _13452_/Y sky130_fd_sc_hd__a21oi_1
X_10664_ _09502_/A _10655_/X _10662_/X _10663_/Y _12385_/C1 vssd1 vssd1 vccd1 vccd1
+ _10664_/X sky130_fd_sc_hd__a221o_2
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12403_ _12403_/A1 _12402_/Y _12403_/B1 vssd1 vssd1 vccd1 vccd1 _12403_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16171_ _16171_/A _16171_/B vssd1 vssd1 vccd1 vccd1 _19609_/D sky130_fd_sc_hd__and2_1
X_13383_ _13383_/A _13383_/B vssd1 vssd1 vccd1 vccd1 _13383_/X sky130_fd_sc_hd__or2_2
X_10595_ _12074_/B1 _10594_/X _12075_/C1 vssd1 vssd1 vccd1 vccd1 _10595_/X sky130_fd_sc_hd__o21a_4
X_12334_ _19654_/Q _19960_/Q _19298_/Q _20085_/Q _12334_/S0 _12411_/C vssd1 vssd1
+ vccd1 vccd1 _12334_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15122_ _15407_/S _15121_/Y _14885_/X vssd1 vssd1 vccd1 vccd1 _15122_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_181_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19930_ _20670_/CLK _19930_/D vssd1 vssd1 vccd1 vccd1 _19930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15053_ _15053_/A vssd1 vssd1 vccd1 vccd1 _15053_/Y sky130_fd_sc_hd__inv_2
X_12265_ _12265_/A _12265_/B vssd1 vssd1 vccd1 vccd1 _12265_/Y sky130_fd_sc_hd__nand2_1
X_14004_ _19168_/Q _14004_/A2 _14004_/B1 _14003_/X _16159_/C1 vssd1 vssd1 vccd1 vccd1
+ _19168_/D sky130_fd_sc_hd__o221a_1
X_11216_ _11213_/X _11214_/X _11215_/X _09731_/A _12430_/S vssd1 vssd1 vccd1 vccd1
+ _11216_/X sky130_fd_sc_hd__a221o_1
XFILLER_269_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19861_ _20862_/CLK _19861_/D vssd1 vssd1 vccd1 vccd1 _19861_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12196_ _12198_/B vssd1 vssd1 vccd1 vccd1 _12284_/B sky130_fd_sc_hd__inv_2
X_18812_ _18486_/Y _20987_/Q _18819_/B vssd1 vssd1 vccd1 vccd1 _18812_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11147_ _11236_/A _11236_/B _10558_/B _10549_/Y vssd1 vssd1 vccd1 vccd1 _11147_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_256_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19792_ _20583_/CLK _19792_/D vssd1 vssd1 vccd1 vccd1 _19792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18743_ _20972_/Q _18290_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18744_/B sky130_fd_sc_hd__mux2_1
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11078_ _12306_/A1 _11066_/X _11067_/X vssd1 vssd1 vccd1 vccd1 _11078_/X sky130_fd_sc_hd__o21a_1
X_15955_ _15955_/A _15981_/B vssd1 vssd1 vccd1 vccd1 _15955_/Y sky130_fd_sc_hd__nand2_1
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput160 dout1[58] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__clkbuf_2
XFILLER_248_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput171 irq[0] vssd1 vssd1 vccd1 vccd1 _12543_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_37_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_264_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14906_ _18149_/S _14906_/B vssd1 vssd1 vccd1 vccd1 _14906_/X sky130_fd_sc_hd__and2b_1
X_10029_ _11234_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10029_/Y sky130_fd_sc_hd__nor2_1
Xinput182 irq[5] vssd1 vssd1 vccd1 vccd1 _12536_/C sky130_fd_sc_hd__clkbuf_2
Xinput193 localMemory_wb_adr_i[12] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_hd__clkbuf_2
X_18674_ _20942_/Q _18682_/B vssd1 vssd1 vccd1 vccd1 _18674_/Y sky130_fd_sc_hd__nand2_1
XFILLER_270_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15886_ _15975_/B2 _13439_/C _15885_/X vssd1 vssd1 vccd1 vccd1 _15893_/A sky130_fd_sc_hd__a21o_1
XFILLER_252_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _20381_/Q _17693_/A1 _17637_/S vssd1 vssd1 vccd1 vccd1 _20381_/D sky130_fd_sc_hd__mux2_1
X_14837_ _11223_/B _12443_/B _14837_/S vssd1 vssd1 vccd1 vccd1 _14837_/X sky130_fd_sc_hd__mux2_1
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17556_ _20316_/Q _17935_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20316_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14768_ _19131_/Q _14774_/A2 _14767_/X _14772_/C1 vssd1 vssd1 vccd1 vccd1 _19508_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_251_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16507_ _19814_/Q _17202_/A1 _16519_/S vssd1 vssd1 vccd1 vccd1 _19814_/D sky130_fd_sc_hd__mux2_1
XFILLER_60_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13719_ _13655_/A _13680_/Y _13718_/Y _13714_/S vssd1 vssd1 vccd1 vccd1 _13719_/X
+ sky130_fd_sc_hd__o211a_1
X_17487_ _17487_/A1 _17486_/Y _16451_/A vssd1 vssd1 vccd1 vccd1 _20278_/D sky130_fd_sc_hd__a21oi_1
XFILLER_20_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14699_ _19458_/Q _17112_/A1 _14699_/S vssd1 vssd1 vccd1 vccd1 _19458_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19226_ _19228_/CLK _19226_/D vssd1 vssd1 vccd1 vccd1 _19226_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16438_ _18863_/A _16438_/B _16442_/C vssd1 vssd1 vccd1 vccd1 _19759_/D sky130_fd_sc_hd__nor3_1
XFILLER_158_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19157_ _19560_/CLK _19157_/D vssd1 vssd1 vccd1 vccd1 _19157_/Q sky130_fd_sc_hd__dfxtp_4
X_16369_ _19733_/Q _16370_/C _19734_/Q vssd1 vssd1 vccd1 vccd1 _16371_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18108_ _20777_/Q _18109_/C _20778_/Q vssd1 vssd1 vccd1 vccd1 _18110_/B sky130_fd_sc_hd__a21oi_1
XFILLER_258_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19088_ _19701_/CLK _19088_/D vssd1 vssd1 vccd1 vccd1 _19088_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_219_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18039_ _20752_/Q _18039_/B vssd1 vssd1 vccd1 vccd1 _18045_/C sky130_fd_sc_hd__and2_4
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20001_ _20004_/CLK _20001_/D vssd1 vssd1 vccd1 vccd1 _20001_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09812_ _11995_/S _09811_/X _09810_/X _11684_/A1 vssd1 vssd1 vccd1 vccd1 _09812_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_98_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ _17538_/C _12342_/A _11305_/B _16454_/A vssd1 vssd1 vccd1 vccd1 _09743_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09674_ _19582_/Q _11061_/A vssd1 vssd1 vccd1 vccd1 _09676_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_255_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20903_ _21010_/CLK _20903_/D vssd1 vssd1 vccd1 vccd1 _20903_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20834_ _21027_/CLK _20834_/D vssd1 vssd1 vccd1 vccd1 _20834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_270_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20765_ _20795_/CLK _20765_/D vssd1 vssd1 vccd1 vccd1 _20765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_210_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20696_ _20719_/CLK _20696_/D vssd1 vssd1 vccd1 vccd1 _20696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10380_ _11242_/A1 _14038_/A2 _10379_/X _11228_/B1 _19858_/Q vssd1 vssd1 vccd1 vccd1
+ _10380_/X sky130_fd_sc_hd__o32a_1
XFILLER_124_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12050_ _19891_/Q _19792_/Q _12053_/S vssd1 vssd1 vccd1 vccd1 _12050_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11001_ _11008_/A1 _20660_/Q _11008_/A3 _10322_/S vssd1 vssd1 vccd1 vccd1 _11001_/X
+ sky130_fd_sc_hd__o31a_1
Xfanout1804 _19700_/Q vssd1 vssd1 vccd1 vccd1 _16769_/S sky130_fd_sc_hd__buf_4
Xfanout1815 _19181_/Q vssd1 vssd1 vccd1 vccd1 _12708_/A sky130_fd_sc_hd__buf_8
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1826 _11345_/S vssd1 vssd1 vccd1 vccd1 _12383_/A sky130_fd_sc_hd__buf_6
XFILLER_132_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1837 _19172_/Q vssd1 vssd1 vccd1 vccd1 _12584_/B sky130_fd_sc_hd__buf_8
XFILLER_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1848 _12584_/C vssd1 vssd1 vccd1 vccd1 _11259_/S sky130_fd_sc_hd__buf_12
Xfanout850 _18157_/Y vssd1 vssd1 vccd1 vccd1 _18296_/S sky130_fd_sc_hd__buf_8
Xfanout861 _14964_/X vssd1 vssd1 vccd1 vccd1 _15337_/A2 sky130_fd_sc_hd__buf_6
Xfanout1859 _10866_/A vssd1 vssd1 vccd1 vccd1 _11118_/A sky130_fd_sc_hd__buf_6
Xfanout872 _15322_/A vssd1 vssd1 vccd1 vccd1 _14971_/A sky130_fd_sc_hd__buf_8
Xfanout883 _16048_/C1 vssd1 vssd1 vccd1 vccd1 _15999_/C1 sky130_fd_sc_hd__clkbuf_4
XFILLER_58_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout894 _18419_/S vssd1 vssd1 vccd1 vccd1 _18421_/S sky130_fd_sc_hd__buf_6
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ _15734_/X _15735_/Y _15739_/X vssd1 vssd1 vccd1 vccd1 _15740_/Y sky130_fd_sc_hd__o21ai_1
X_12952_ _18134_/A _16714_/C _16714_/B vssd1 vssd1 vccd1 vccd1 _12952_/X sky130_fd_sc_hd__or3b_4
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _11903_/A1 _11889_/X _11890_/X vssd1 vssd1 vccd1 vccd1 _11903_/X sky130_fd_sc_hd__o21a_1
XFILLER_234_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15671_ _16000_/A1 _15660_/X _15661_/X _15670_/X vssd1 vssd1 vccd1 vccd1 _15671_/X
+ sky130_fd_sc_hd__a22o_4
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_210 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12911_/A _12883_/B vssd1 vssd1 vccd1 vccd1 _13209_/A sky130_fd_sc_hd__xnor2_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17410_ _20259_/Q _20251_/Q _17442_/A vssd1 vssd1 vccd1 vccd1 _17410_/X sky130_fd_sc_hd__mux2_1
XANTENNA_243 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _19386_/Q _17906_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19386_/D sky130_fd_sc_hd__mux2_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _18390_/A _18981_/C _18755_/B vssd1 vssd1 vccd1 vccd1 _18395_/S sky130_fd_sc_hd__nor3_4
XANTENNA_254 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11834_ _19822_/Q _19326_/Q _11987_/S vssd1 vssd1 vccd1 vccd1 _11834_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_276 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _20219_/Q _17371_/A2 _17340_/X _18702_/A vssd1 vssd1 vccd1 vccd1 _20219_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_287 input216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14553_ _19323_/Q _17835_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19323_/D sky130_fd_sc_hd__mux2_1
XANTENNA_298 input227/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ _11764_/B _15433_/A _13459_/A vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_82_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _19606_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13504_ _20948_/Q _20882_/Q _13060_/C _13060_/D vssd1 vssd1 vccd1 vccd1 _13504_/X
+ sky130_fd_sc_hd__a22o_1
X_10716_ _15150_/C1 _15331_/A _10685_/Y vssd1 vssd1 vccd1 vccd1 _10802_/B sky130_fd_sc_hd__o21ba_4
X_17272_ _17272_/A _17275_/B _17290_/C vssd1 vssd1 vccd1 vccd1 _17272_/X sky130_fd_sc_hd__and3_1
XFILLER_158_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14484_ _18746_/A _14484_/B vssd1 vssd1 vccd1 vccd1 _19266_/D sky130_fd_sc_hd__and2_1
X_11696_ _20479_/Q _11718_/S _11708_/B _11694_/X _11695_/X vssd1 vssd1 vccd1 vccd1
+ _11696_/X sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20579_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19011_ _21025_/Q _19015_/B vssd1 vssd1 vccd1 vccd1 _19011_/X sky130_fd_sc_hd__or2_1
XFILLER_174_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16223_ _19646_/Q _17107_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19646_/D sky130_fd_sc_hd__mux2_1
X_10647_ _19872_/Q _19773_/Q _12381_/S vssd1 vssd1 vccd1 vccd1 _10647_/X sky130_fd_sc_hd__mux2_1
X_13435_ _16066_/B _15898_/A _13439_/C _15843_/A vssd1 vssd1 vccd1 vccd1 _13436_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16154_ _16824_/B _16178_/S vssd1 vssd1 vccd1 vccd1 _16154_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13366_ _13334_/A _13365_/Y _13364_/X _13366_/C1 vssd1 vssd1 vccd1 vccd1 _13366_/X
+ sky130_fd_sc_hd__a211o_1
X_10578_ _11514_/A1 _20698_/Q _11676_/S _10576_/X _10577_/X vssd1 vssd1 vccd1 vccd1
+ _10578_/X sky130_fd_sc_hd__a311o_1
XFILLER_115_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105_ _15067_/X _15104_/X _15254_/S vssd1 vssd1 vccd1 vccd1 _15105_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12317_ _12315_/X _12316_/X _12317_/S vssd1 vssd1 vccd1 vccd1 _12317_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16085_ _19567_/Q _16067_/X _16143_/A vssd1 vssd1 vccd1 vccd1 _16085_/X sky130_fd_sc_hd__o21a_1
XFILLER_182_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13297_ _20933_/Q _13350_/B _18671_/B vssd1 vssd1 vccd1 vccd1 _13297_/Y sky130_fd_sc_hd__a21oi_1
X_12248_ _12337_/A _19926_/Q _12248_/B1 _20051_/Q vssd1 vssd1 vccd1 vccd1 _12248_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_244_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15036_ _14857_/X _14862_/A _15062_/S vssd1 vssd1 vccd1 vccd1 _15036_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19913_ _20573_/CLK _19913_/D vssd1 vssd1 vccd1 vccd1 _19913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_268_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_257_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19844_ _20751_/CLK _19844_/D vssd1 vssd1 vccd1 vccd1 _19844_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_268_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12179_ _12189_/A _12178_/X _12177_/X _11851_/C vssd1 vssd1 vccd1 vccd1 _12179_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_257_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19775_ _20706_/CLK _19775_/D vssd1 vssd1 vccd1 vccd1 _19775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_256_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16987_ _19244_/Q _16996_/A2 _17005_/A2 _19113_/Q _16945_/X vssd1 vssd1 vccd1 vccd1
+ _16987_/X sky130_fd_sc_hd__o221a_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18726_ _18726_/A _18726_/B vssd1 vssd1 vccd1 vccd1 _20963_/D sky130_fd_sc_hd__and2_1
XFILLER_97_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15938_ _20941_/Q _16044_/A2 _15937_/X vssd1 vssd1 vccd1 vccd1 _15938_/X sky130_fd_sc_hd__o21a_1
XFILLER_265_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_264_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18657_ _18960_/A _18657_/B vssd1 vssd1 vccd1 vccd1 _20937_/D sky130_fd_sc_hd__nor2_1
X_15869_ _19551_/Q _15980_/A2 _15867_/X _15868_/X _17432_/A vssd1 vssd1 vccd1 vccd1
+ _19551_/D sky130_fd_sc_hd__o221a_1
XFILLER_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17608_ _17745_/A _17676_/B _17608_/C vssd1 vssd1 vccd1 vccd1 _17608_/X sky130_fd_sc_hd__and3_4
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18588_ _20920_/Q _18619_/B vssd1 vssd1 vccd1 vccd1 _18588_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_252_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17539_ _17812_/A _17675_/B vssd1 vssd1 vccd1 vccd1 _17540_/C sky130_fd_sc_hd__nor2_1
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20550_ _20682_/CLK _20550_/D vssd1 vssd1 vccd1 vccd1 _20550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19209_ _20665_/CLK _19209_/D vssd1 vssd1 vccd1 vccd1 _19209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_192_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20481_ _20481_/CLK _20481_/D vssd1 vssd1 vccd1 vccd1 _20481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput420 _19980_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[19] sky130_fd_sc_hd__buf_4
XFILLER_218_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput431 _19990_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[29] sky130_fd_sc_hd__buf_4
Xoutput442 _19994_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_stall_o sky130_fd_sc_hd__buf_4
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput453 _19506_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[12] sky130_fd_sc_hd__buf_4
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput464 _19516_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[22] sky130_fd_sc_hd__buf_4
Xoutput475 _19497_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[3] sky130_fd_sc_hd__buf_4
XFILLER_232_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput486 _13825_/X vssd1 vssd1 vccd1 vccd1 wmask0[2] sky130_fd_sc_hd__buf_6
X_21033_ _21042_/CLK _21033_/D vssd1 vssd1 vccd1 vccd1 _21033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_275_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_259_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09726_ _11922_/A1 _13734_/A _12158_/B1 vssd1 vssd1 vccd1 vccd1 _09726_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_228_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09657_ _11228_/A1 _13969_/A2 _09656_/X _11242_/B1 _19838_/Q vssd1 vssd1 vccd1 vccd1
+ _09657_/X sky130_fd_sc_hd__o32a_1
XFILLER_242_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09588_ _19087_/Q _19086_/Q _09588_/C _09592_/B vssd1 vssd1 vccd1 vccd1 _09588_/X
+ sky130_fd_sc_hd__and4_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20817_ _21022_/CLK _20817_/D vssd1 vssd1 vccd1 vccd1 _20817_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11550_ _12191_/C1 _12006_/S _11549_/X _10409_/A vssd1 vssd1 vccd1 vccd1 _11550_/X
+ sky130_fd_sc_hd__a31o_1
X_20748_ _20812_/CLK _20748_/D vssd1 vssd1 vccd1 vccd1 _20748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10501_ _11266_/A1 _19312_/Q _11270_/A2 _10322_/S vssd1 vssd1 vccd1 vccd1 _10501_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_211_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11481_ _11479_/X _11480_/X _12189_/A vssd1 vssd1 vccd1 vccd1 _11481_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20679_ _20679_/CLK _20679_/D vssd1 vssd1 vccd1 vccd1 _20679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13220_ _13220_/A vssd1 vssd1 vccd1 vccd1 _13220_/Y sky130_fd_sc_hd__clkinv_2
X_10432_ _11281_/A _20600_/Q _11268_/C vssd1 vssd1 vccd1 vccd1 _10432_/X sky130_fd_sc_hd__and3_1
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13151_ _10719_/Y _13150_/A _13150_/B _10720_/A vssd1 vssd1 vccd1 vccd1 _13570_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10363_ _19508_/Q _15561_/A _11726_/S vssd1 vssd1 vccd1 vccd1 _11414_/B sky130_fd_sc_hd__mux2_4
XFILLER_152_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12102_ _12102_/A1 _20391_/Q _20455_/Q _12097_/S vssd1 vssd1 vccd1 vccd1 _12102_/X
+ sky130_fd_sc_hd__a22o_1
X_13082_ _13021_/Y _13395_/A _13394_/B vssd1 vssd1 vccd1 vccd1 _13258_/C sky130_fd_sc_hd__o21ai_4
X_10294_ _19541_/Q _09596_/B _10280_/X _10293_/Y vssd1 vssd1 vccd1 vccd1 _10294_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_151_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16910_ _16885_/A _16909_/X _16740_/B2 vssd1 vssd1 vccd1 vccd1 _16910_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _12035_/B vssd1 vssd1 vccd1 vccd1 _12033_/Y sky130_fd_sc_hd__inv_2
Xfanout1601 _09618_/Y vssd1 vssd1 vccd1 vccd1 _11833_/C1 sky130_fd_sc_hd__buf_4
XFILLER_78_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17890_ _20661_/Q _17890_/A1 _17917_/S vssd1 vssd1 vccd1 vccd1 _20661_/D sky130_fd_sc_hd__mux2_1
Xfanout1612 _11513_/S vssd1 vssd1 vccd1 vccd1 _11980_/S sky130_fd_sc_hd__buf_6
XFILLER_78_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1623 fanout1630/X vssd1 vssd1 vccd1 vccd1 _10152_/S sky130_fd_sc_hd__buf_6
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1634 _09615_/Y vssd1 vssd1 vccd1 vccd1 _12385_/C1 sky130_fd_sc_hd__buf_4
X_16841_ _19972_/Q _16876_/A _16840_/Y _16896_/C1 vssd1 vssd1 vccd1 vccd1 _19972_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1645 _18949_/A2 vssd1 vssd1 vccd1 vccd1 _12533_/B sky130_fd_sc_hd__buf_6
XFILLER_265_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1656 _09655_/Y vssd1 vssd1 vccd1 vccd1 _13969_/A2 sky130_fd_sc_hd__buf_4
XFILLER_38_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_266_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1667 _14112_/B vssd1 vssd1 vccd1 vccd1 _09734_/B sky130_fd_sc_hd__buf_12
Xfanout680 _14004_/A2 vssd1 vssd1 vccd1 vccd1 _16605_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_144_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1678 _12008_/A vssd1 vssd1 vccd1 vccd1 _11946_/A1 sky130_fd_sc_hd__buf_6
X_19560_ _19560_/CLK _19560_/D vssd1 vssd1 vccd1 vccd1 _19560_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1689 _11026_/A vssd1 vssd1 vccd1 vccd1 _11290_/A sky130_fd_sc_hd__buf_4
Xfanout691 split9/A vssd1 vssd1 vccd1 vccd1 _13805_/B1 sky130_fd_sc_hd__buf_6
XFILLER_219_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16772_ _16768_/Y _16771_/X _17011_/B1 vssd1 vssd1 vccd1 vccd1 _16772_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_265_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13984_ _14002_/A1 _09664_/B _10025_/X _14002_/B1 _19843_/Q vssd1 vssd1 vccd1 vccd1
+ _14069_/C sky130_fd_sc_hd__o32a_1
XFILLER_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18511_ _18628_/B _18511_/B vssd1 vssd1 vccd1 vccd1 _18511_/X sky130_fd_sc_hd__or2_1
X_15723_ _20805_/Q _15941_/A2 _15716_/X _15882_/A1 _15722_/X vssd1 vssd1 vccd1 vccd1
+ _15723_/X sky130_fd_sc_hd__a221o_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19491_ _20468_/CLK _19491_/D vssd1 vssd1 vccd1 vccd1 _19491_/Q sky130_fd_sc_hd__dfxtp_1
X_12935_ _19262_/Q _12950_/B2 _16716_/A _20010_/Q vssd1 vssd1 vccd1 vccd1 _14899_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_46_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18442_ _18748_/A _18442_/B vssd1 vssd1 vccd1 vccd1 _20875_/D sky130_fd_sc_hd__and2_1
XFILLER_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15654_ _16053_/A _15654_/B vssd1 vssd1 vccd1 vccd1 _15654_/Y sky130_fd_sc_hd__nor2_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12866_ _12866_/A _12866_/B vssd1 vssd1 vccd1 vccd1 _13362_/B sky130_fd_sc_hd__nor2_2
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14605_ _19369_/Q _17889_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19369_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11817_ _19889_/Q _19790_/Q _11891_/B vssd1 vssd1 vccd1 vccd1 _11817_/X sky130_fd_sc_hd__mux2_1
X_18373_ _18538_/B _18385_/B vssd1 vssd1 vccd1 vccd1 _18373_/Y sky130_fd_sc_hd__nand2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _14815_/S _15654_/B _15584_/Y _15365_/A vssd1 vssd1 vccd1 vccd1 _15585_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _13448_/A _12771_/C _12771_/D _12795_/X _12796_/X vssd1 vssd1 vccd1 vccd1
+ _13279_/A sky130_fd_sc_hd__a41o_2
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _20213_/Q _17356_/A2 _17302_/C _17323_/X _17324_/C1 vssd1 vssd1 vccd1 vccd1
+ _17324_/X sky130_fd_sc_hd__a221o_1
X_14536_ _19306_/Q _17750_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19306_/D sky130_fd_sc_hd__mux2_1
XFILLER_42_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11748_ _13413_/A _11748_/B vssd1 vssd1 vccd1 vccd1 _11748_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17255_ _20190_/Q _17235_/Y _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17255_/X sky130_fd_sc_hd__a21o_1
XFILLER_187_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14467_ _20229_/Q _19258_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14468_/B sky130_fd_sc_hd__mux2_1
XFILLER_175_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ _19816_/Q _19320_/Q _11994_/S vssd1 vssd1 vccd1 vccd1 _11679_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16206_ _19629_/Q _17683_/A1 _16230_/S vssd1 vssd1 vccd1 vccd1 _19629_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13418_ _13418_/A _13418_/B vssd1 vssd1 vccd1 vccd1 _13428_/C sky130_fd_sc_hd__xor2_4
XFILLER_128_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17186_ _20150_/Q _17780_/A1 _17215_/S vssd1 vssd1 vccd1 vccd1 _20150_/D sky130_fd_sc_hd__mux2_1
XFILLER_190_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14398_ _19242_/Q _14398_/A2 _14397_/X _14794_/C1 vssd1 vssd1 vccd1 vccd1 _19242_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_217_wb_clk_i clkbuf_leaf_4_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20481_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _19592_/Q _16196_/S _16136_/Y _16165_/C1 vssd1 vssd1 vccd1 vccd1 _19592_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13349_ _19230_/Q _13403_/B _19231_/Q vssd1 vssd1 vccd1 vccd1 _13349_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_255_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ _16068_/A _16068_/B _16068_/C vssd1 vssd1 vccd1 vccd1 _16068_/Y sky130_fd_sc_hd__nand3_4
XFILLER_64_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15019_ _15019_/A _15019_/B _15019_/C vssd1 vssd1 vccd1 vccd1 _15134_/B sky130_fd_sc_hd__nand3_2
XFILLER_151_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19827_ _20662_/CLK _19827_/D vssd1 vssd1 vccd1 vccd1 _19827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_256_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_257_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19758_ _20742_/CLK _19758_/D vssd1 vssd1 vccd1 vccd1 _19758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ _19091_/Q vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__inv_2
X_18709_ _20955_/Q _18205_/Y _18719_/S vssd1 vssd1 vccd1 vccd1 _18710_/B sky130_fd_sc_hd__mux2_1
XFILLER_253_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19689_ _20716_/CLK _19689_/D vssd1 vssd1 vccd1 vccd1 _19689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20602_ _20638_/CLK _20602_/D vssd1 vssd1 vccd1 vccd1 _20602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20533_ _20633_/CLK _20533_/D vssd1 vssd1 vccd1 vccd1 _20533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20464_ _20565_/CLK _20464_/D vssd1 vssd1 vccd1 vccd1 _20464_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20395_ _20468_/CLK _20395_/D vssd1 vssd1 vccd1 vccd1 _20395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_279_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput294 _13781_/X vssd1 vssd1 vccd1 vccd1 addr1[0] sky130_fd_sc_hd__buf_4
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21016_ _21016_/CLK _21016_/D vssd1 vssd1 vccd1 vccd1 _21016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_256_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09709_ _11981_/C1 _09708_/X _09705_/X _12137_/C1 vssd1 vssd1 vccd1 vccd1 _09709_/X
+ sky130_fd_sc_hd__a211o_2
X_10981_ _20368_/Q _20432_/Q _10986_/B vssd1 vssd1 vccd1 vccd1 _10981_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12720_ _15561_/A _12731_/B vssd1 vssd1 vccd1 vccd1 _12720_/Y sky130_fd_sc_hd__nand2_1
XFILLER_215_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ _19499_/Q _12758_/B vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__and2_1
XFILLER_130_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11602_ _19817_/Q _19321_/Q _11965_/B vssd1 vssd1 vccd1 vccd1 _11602_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15370_ _11788_/B _15127_/B _15369_/X _12579_/D vssd1 vssd1 vccd1 vccd1 _15378_/A
+ sky130_fd_sc_hd__o211a_1
X_12582_ _14112_/B _16066_/A _12582_/C _15095_/B vssd1 vssd1 vccd1 vccd1 _12583_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_196_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14321_ _19514_/Q _14322_/B vssd1 vssd1 vccd1 vccd1 _14333_/A sky130_fd_sc_hd__nand2_1
XFILLER_90_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ _19543_/Q _12365_/A2 _09607_/X _19607_/Q vssd1 vssd1 vccd1 vccd1 _11533_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_278_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17040_ _20018_/Q _13466_/A _17040_/S vssd1 vssd1 vccd1 vccd1 _20018_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11464_ _12186_/S _11464_/B vssd1 vssd1 vccd1 vccd1 _11464_/X sky130_fd_sc_hd__or2_1
X_14252_ _14262_/A _14252_/B _14260_/B vssd1 vssd1 vccd1 vccd1 _14252_/X sky130_fd_sc_hd__or3b_1
XFILLER_99_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13203_ _13002_/A _12664_/C _13199_/Y _13202_/X _13366_/C1 vssd1 vssd1 vccd1 vccd1
+ _13203_/X sky130_fd_sc_hd__a311o_2
X_10415_ _12088_/S _10414_/X _12105_/A vssd1 vssd1 vccd1 vccd1 _10415_/X sky130_fd_sc_hd__o21a_1
X_11395_ _11389_/X _11394_/X _12415_/S vssd1 vssd1 vccd1 vccd1 _11395_/X sky130_fd_sc_hd__mux2_1
X_14183_ _14202_/S _14177_/B _14182_/Y _18763_/A1 vssd1 vssd1 vccd1 vccd1 _14183_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10346_ _10344_/X _10345_/X _12426_/S vssd1 vssd1 vccd1 vccd1 _10346_/X sky130_fd_sc_hd__mux2_1
X_13134_ _13007_/Y _13134_/B vssd1 vssd1 vccd1 vccd1 _13135_/B sky130_fd_sc_hd__nand2b_1
X_18991_ _21015_/Q _19013_/B vssd1 vssd1 vccd1 vccd1 _18991_/X sky130_fd_sc_hd__or2_1
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13065_ _13051_/X _13064_/X _13049_/Y _13050_/X vssd1 vssd1 vccd1 vccd1 _13563_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _20711_/Q _17942_/A1 _17946_/S vssd1 vssd1 vccd1 vccd1 _20711_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10277_ _10277_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _10278_/B sky130_fd_sc_hd__or2_4
XFILLER_124_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1420 _12272_/B2 vssd1 vssd1 vccd1 vccd1 _11116_/S sky130_fd_sc_hd__buf_6
X_12016_ _09752_/A _20392_/Q _20456_/Q _12013_/S _12016_/C1 vssd1 vssd1 vccd1 vccd1
+ _12016_/X sky130_fd_sc_hd__a221o_1
Xfanout1431 _12190_/C1 vssd1 vssd1 vccd1 vccd1 _11563_/S sky130_fd_sc_hd__buf_6
X_17873_ _20646_/Q _17907_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20646_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1442 _10611_/B vssd1 vssd1 vccd1 vccd1 _12003_/C sky130_fd_sc_hd__buf_6
Xfanout1453 _11191_/C vssd1 vssd1 vccd1 vccd1 _11021_/C sky130_fd_sc_hd__buf_6
Xfanout1464 _09744_/B vssd1 vssd1 vccd1 vccd1 _10409_/A sky130_fd_sc_hd__clkbuf_16
Xfanout1475 _12414_/S vssd1 vssd1 vccd1 vccd1 _12340_/S sky130_fd_sc_hd__buf_8
X_16824_ _16878_/A _16824_/B vssd1 vssd1 vccd1 vccd1 _16824_/Y sky130_fd_sc_hd__nand2_1
X_19612_ _20263_/CLK _19612_/D vssd1 vssd1 vccd1 vccd1 _19612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1486 _09729_/Y vssd1 vssd1 vccd1 vccd1 _12105_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_281_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1497 _12041_/B vssd1 vssd1 vccd1 vccd1 _12043_/B sky130_fd_sc_hd__buf_6
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19543_ _19607_/CLK _19543_/D vssd1 vssd1 vccd1 vccd1 _19543_/Q sky130_fd_sc_hd__dfxtp_1
X_16755_ _20400_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16755_/X sky130_fd_sc_hd__a21o_1
X_13967_ _19188_/Q _14057_/C _13967_/S vssd1 vssd1 vccd1 vccd1 _13967_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15706_ _19545_/Q _16007_/A _15705_/X _16189_/A vssd1 vssd1 vccd1 vccd1 _19545_/D
+ sky130_fd_sc_hd__o211a_1
X_12918_ _12912_/A _12913_/X _12917_/Y vssd1 vssd1 vccd1 vccd1 _12918_/Y sky130_fd_sc_hd__a21oi_1
X_19474_ _20451_/CLK _19474_/D vssd1 vssd1 vccd1 vccd1 _19474_/Q sky130_fd_sc_hd__dfxtp_1
X_16686_ _19941_/Q _17096_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19941_/D sky130_fd_sc_hd__mux2_1
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13898_ _19115_/Q _14527_/A2 _13897_/X _16193_/A vssd1 vssd1 vccd1 vccd1 _19115_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_181_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_261_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18425_ _20867_/Q _18245_/Y _18449_/S vssd1 vssd1 vccd1 vccd1 _18426_/B sky130_fd_sc_hd__mux2_1
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15637_ _20930_/Q _15995_/A2 _15636_/X vssd1 vssd1 vccd1 vccd1 _15637_/X sky130_fd_sc_hd__o21a_1
X_12849_ _19511_/Q _12857_/B vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__or2_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18356_ _20833_/Q _18357_/B _18355_/Y _18724_/A vssd1 vssd1 vccd1 vccd1 _20833_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _20960_/Q _15568_/A2 _15568_/B1 _20832_/Q _15567_/X vssd1 vssd1 vccd1 vccd1
+ _15568_/X sky130_fd_sc_hd__a221o_4
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17307_ _20208_/Q _17328_/A2 _17305_/X _17306_/X _17974_/B1 vssd1 vssd1 vccd1 vccd1
+ _20208_/D sky130_fd_sc_hd__o221a_1
XFILLER_148_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14519_ _19297_/Q _17707_/A1 _14519_/S vssd1 vssd1 vccd1 vccd1 _19297_/D sky130_fd_sc_hd__mux2_1
X_18287_ _18746_/A _18287_/B vssd1 vssd1 vccd1 vccd1 _20811_/D sky130_fd_sc_hd__and2_1
X_15499_ _15612_/S _15164_/X _15610_/B1 vssd1 vssd1 vccd1 vccd1 _15499_/X sky130_fd_sc_hd__a21bo_1
XFILLER_174_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17238_ _20185_/Q _17268_/A2 _17237_/X _17241_/C1 vssd1 vssd1 vccd1 vccd1 _20185_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17169_ _20135_/Q _17869_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20135_/D sky130_fd_sc_hd__mux2_1
XFILLER_155_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20180_ _20180_/CLK _20180_/D vssd1 vssd1 vccd1 vccd1 _20180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09991_ _11851_/A _20677_/Q _11851_/C vssd1 vssd1 vccd1 vccd1 _09991_/X sky130_fd_sc_hd__or3_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_253_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_139_wb_clk_i _19214_/CLK vssd1 vssd1 vccd1 vccd1 _19701_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20516_ _20717_/CLK _20516_/D vssd1 vssd1 vccd1 vccd1 _20516_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_181_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20447_ _20715_/CLK _20447_/D vssd1 vssd1 vccd1 vccd1 _20447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10200_ _11326_/A _11234_/B _09680_/X vssd1 vssd1 vccd1 vccd1 _10201_/B sky130_fd_sc_hd__a21o_1
XFILLER_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11180_ _11101_/A _11178_/X _11179_/X _11176_/X _12302_/S vssd1 vssd1 vccd1 vccd1
+ _11180_/X sky130_fd_sc_hd__a311o_1
X_20378_ _20570_/CLK _20378_/D vssd1 vssd1 vccd1 vccd1 _20378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10131_ _19675_/Q _20163_/Q _12375_/S vssd1 vssd1 vccd1 vccd1 _10131_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10062_ _20409_/Q _10502_/A2 _10059_/X _10060_/X _10061_/X vssd1 vssd1 vccd1 vccd1
+ _10062_/X sky130_fd_sc_hd__o221a_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_276_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14870_ _11054_/B _12284_/B _14870_/S vssd1 vssd1 vccd1 vccd1 _14870_/X sky130_fd_sc_hd__mux2_1
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13821_ _13822_/A1 _13775_/B split9/X input238/X vssd1 vssd1 vccd1 vccd1 _13821_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_251_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16540_ _19836_/Q _16578_/A2 _16578_/B1 input37/X vssd1 vssd1 vccd1 vccd1 _16541_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13752_ _13777_/A _13752_/B vssd1 vssd1 vccd1 vccd1 _13752_/X sky130_fd_sc_hd__or2_1
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10964_ _10954_/X _10963_/Y _11201_/A _10946_/X vssd1 vssd1 vccd1 vccd1 _10964_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_250_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12703_ _12855_/B _12703_/B vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__or2_1
X_16471_ _19780_/Q _17657_/A1 _16471_/S vssd1 vssd1 vccd1 vccd1 _19780_/D sky130_fd_sc_hd__mux2_1
XFILLER_245_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13683_ _13775_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__and2_1
XFILLER_70_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10895_ _11268_/A _20593_/Q _11261_/C vssd1 vssd1 vccd1 vccd1 _10895_/X sky130_fd_sc_hd__and3_1
X_18210_ _18496_/B vssd1 vssd1 vccd1 vccd1 _18210_/Y sky130_fd_sc_hd__clkinv_4
X_15422_ _17266_/A _15421_/X _15452_/S vssd1 vssd1 vccd1 vccd1 _15422_/X sky130_fd_sc_hd__mux2_1
XPHY_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19190_ _20670_/CLK _19190_/D vssd1 vssd1 vccd1 vccd1 _19190_/Q sky130_fd_sc_hd__dfxtp_1
X_12634_ _12634_/A _12744_/B vssd1 vssd1 vccd1 vccd1 _12634_/Y sky130_fd_sc_hd__nor2_2
XPHY_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18141_ _18389_/A vssd1 vssd1 vccd1 vccd1 _18319_/A sky130_fd_sc_hd__inv_2
XFILLER_86_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15353_ _14888_/X _15352_/X _15611_/S vssd1 vssd1 vccd1 vccd1 _15354_/A sky130_fd_sc_hd__mux2_2
X_12565_ _13657_/A _12565_/B vssd1 vssd1 vccd1 vccd1 _13684_/B sky130_fd_sc_hd__nor2_8
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ _14304_/A _14304_/B vssd1 vssd1 vccd1 vccd1 _14304_/Y sky130_fd_sc_hd__xnor2_1
X_18072_ _18080_/A _18077_/C vssd1 vssd1 vccd1 vccd1 _18072_/Y sky130_fd_sc_hd__nor2_1
X_11516_ _11981_/C1 _11515_/X _11512_/X _12137_/C1 vssd1 vssd1 vccd1 vccd1 _11516_/X
+ sky130_fd_sc_hd__a211o_1
X_15284_ _15283_/B _15282_/X _15283_/Y _15673_/B1 _15246_/A vssd1 vssd1 vccd1 vccd1
+ _15284_/X sky130_fd_sc_hd__a221o_1
X_12496_ _12496_/A _12496_/B vssd1 vssd1 vccd1 vccd1 _12498_/A sky130_fd_sc_hd__xnor2_2
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17023_ _20001_/Q input210/X _17026_/S vssd1 vssd1 vccd1 vccd1 _20001_/D sky130_fd_sc_hd__mux2_1
X_14235_ _14255_/A _16068_/B _14235_/C vssd1 vssd1 vccd1 vccd1 _14235_/X sky130_fd_sc_hd__or3_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ _19284_/Q _20071_/Q _12146_/S vssd1 vssd1 vccd1 vccd1 _11447_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11378_ _11376_/X _11377_/X _11378_/S vssd1 vssd1 vccd1 vccd1 _11378_/X sky130_fd_sc_hd__mux2_1
X_14166_ _19219_/Q _14256_/A2 _14165_/X _18698_/A vssd1 vssd1 vccd1 vccd1 _19219_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_252_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10329_ _12402_/A1 _17866_/A1 _10328_/X vssd1 vssd1 vccd1 vccd1 _13693_/A sky130_fd_sc_hd__o21ai_4
XFILLER_140_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13117_ _12909_/X _13107_/Y _13116_/Y _13323_/C vssd1 vssd1 vccd1 vccd1 _13117_/X
+ sky130_fd_sc_hd__a31o_1
X_14097_ _14099_/A _14099_/B _14097_/C vssd1 vssd1 vccd1 vccd1 _14097_/X sky130_fd_sc_hd__or3_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18974_ _19115_/Q _18974_/A2 _18974_/B1 _13181_/B vssd1 vssd1 vccd1 vccd1 _18975_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_267_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17925_ _20694_/Q _17925_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20694_/D sky130_fd_sc_hd__mux2_1
X_13048_ _20954_/Q _20888_/Q vssd1 vssd1 vccd1 vccd1 _13048_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1250 _17381_/A2 vssd1 vssd1 vccd1 vccd1 _17401_/A2 sky130_fd_sc_hd__buf_4
XFILLER_38_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1261 _12730_/A2 vssd1 vssd1 vccd1 vccd1 _12657_/A2 sky130_fd_sc_hd__buf_2
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17856_ _20629_/Q _17890_/A1 _17883_/S vssd1 vssd1 vccd1 vccd1 _20629_/D sky130_fd_sc_hd__mux2_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1272 _15303_/A vssd1 vssd1 vccd1 vccd1 _15975_/B2 sky130_fd_sc_hd__buf_4
XFILLER_227_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1283 _09547_/X vssd1 vssd1 vccd1 vccd1 _11189_/B sky130_fd_sc_hd__buf_4
XFILLER_281_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1294 _12708_/B vssd1 vssd1 vccd1 vccd1 _15703_/B2 sky130_fd_sc_hd__buf_8
X_16807_ _19223_/Q _16996_/A2 _17005_/A2 _19092_/Q _16806_/X vssd1 vssd1 vccd1 vccd1
+ _16807_/X sky130_fd_sc_hd__o221a_1
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_282_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17787_ _20564_/Q _17927_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20564_/D sky130_fd_sc_hd__mux2_1
X_14999_ _15314_/B _15314_/C _15314_/D vssd1 vssd1 vccd1 vccd1 _14999_/X sky130_fd_sc_hd__or3_1
XFILLER_254_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19526_ _19697_/CLK _19526_/D vssd1 vssd1 vccd1 vccd1 _19526_/Q sky130_fd_sc_hd__dfxtp_1
X_16738_ _16799_/S input69/X vssd1 vssd1 vccd1 vccd1 _16738_/Y sky130_fd_sc_hd__nand2_1
XFILLER_235_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_222_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19457_ _20580_/CLK _19457_/D vssd1 vssd1 vccd1 vccd1 _19457_/Q sky130_fd_sc_hd__dfxtp_1
X_16669_ _19926_/Q _17915_/A1 _16671_/S vssd1 vssd1 vccd1 vccd1 _19926_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18408_ _18708_/A _18408_/B vssd1 vssd1 vccd1 vccd1 _20858_/D sky130_fd_sc_hd__and2_1
X_19388_ _20679_/CLK _19388_/D vssd1 vssd1 vccd1 vccd1 _19388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18339_ _18487_/B _18349_/B vssd1 vssd1 vccd1 vccd1 _18339_/Y sky130_fd_sc_hd__nand2_1
XFILLER_277_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20301_ _21047_/A _20301_/D vssd1 vssd1 vccd1 vccd1 _20301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20232_ _20990_/CLK _20232_/D vssd1 vssd1 vccd1 vccd1 _20232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20163_ _20180_/CLK _20163_/D vssd1 vssd1 vccd1 vccd1 _20163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _19818_/Q _19322_/Q _12121_/S vssd1 vssd1 vccd1 vccd1 _09974_/X sky130_fd_sc_hd__mux2_1
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20094_ _20720_/CLK _20094_/D vssd1 vssd1 vccd1 vccd1 _20094_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_272_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_260_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_606 _20624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_617 _13775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_628 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ _21025_/CLK _20996_/D vssd1 vssd1 vccd1 vccd1 _20996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_639 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10680_ _19534_/Q _12365_/A2 _11225_/B _19598_/Q vssd1 vssd1 vccd1 vccd1 _10680_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12350_ _10866_/A _12348_/Y _12349_/Y vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__a21o_1
XFILLER_275_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11301_ _11297_/X _11300_/X _12514_/C vssd1 vssd1 vccd1 vccd1 _11301_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12281_ _12283_/A vssd1 vssd1 vccd1 vccd1 _12281_/Y sky130_fd_sc_hd__inv_2
X_14020_ _14035_/A1 _14038_/A2 _11227_/X _14035_/B1 _19855_/Q vssd1 vssd1 vccd1 vccd1
+ _14093_/C sky130_fd_sc_hd__o32a_1
X_11232_ _11239_/A1 _13978_/A2 _11231_/X _11239_/B1 _19839_/Q vssd1 vssd1 vccd1 vccd1
+ _11232_/X sky130_fd_sc_hd__o32a_1
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11163_ _12398_/C1 _11161_/X _11162_/X _12317_/S vssd1 vssd1 vccd1 vccd1 _11163_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20315_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10114_ _19540_/Q _09596_/A _11225_/B _19604_/Q _11246_/A1 vssd1 vssd1 vccd1 vccd1
+ _10114_/X sky130_fd_sc_hd__a221o_1
XFILLER_150_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_267_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11094_ _11092_/X _11093_/X _11094_/S vssd1 vssd1 vccd1 vccd1 _11094_/X sky130_fd_sc_hd__mux2_1
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15971_ _19762_/Q _15999_/A2 _15970_/X _15971_/C1 vssd1 vssd1 vccd1 vccd1 _15971_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_121_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17710_ _17918_/A _17850_/B vssd1 vssd1 vccd1 vccd1 _17711_/C sky130_fd_sc_hd__nor2_1
XFILLER_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14922_ _14917_/A _19177_/Q _14921_/X vssd1 vssd1 vccd1 vccd1 _14973_/B sky130_fd_sc_hd__a21o_4
X_10045_ _19539_/Q _09596_/B _10019_/X _10044_/Y vssd1 vssd1 vccd1 vccd1 _10045_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18690_ _18690_/A _18755_/B vssd1 vssd1 vccd1 vccd1 _18690_/Y sky130_fd_sc_hd__nor2_8
XFILLER_121_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_248_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _17918_/A _17675_/B vssd1 vssd1 vccd1 vccd1 _17642_/C sky130_fd_sc_hd__nor2_1
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_263_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14853_ _11411_/B _11733_/B _14853_/S vssd1 vssd1 vccd1 vccd1 _14853_/X sky130_fd_sc_hd__mux2_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _13822_/A1 _13691_/Y _13790_/X input219/X vssd1 vssd1 vccd1 vccd1 _13804_/X
+ sky130_fd_sc_hd__a22o_1
X_17572_ _20332_/Q _17708_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20332_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_263_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14784_ _19139_/Q _14802_/A2 _14783_/X _17434_/A vssd1 vssd1 vccd1 vccd1 _19516_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11996_ _12151_/A1 _11995_/X _11992_/X _12151_/C1 vssd1 vssd1 vccd1 vccd1 _11996_/X
+ sky130_fd_sc_hd__o211a_1
X_19311_ _20438_/CLK _19311_/D vssd1 vssd1 vccd1 vccd1 _19311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16523_ _19864_/Q _19863_/Q vssd1 vssd1 vccd1 vccd1 _16594_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13735_ _13735_/A _13735_/B vssd1 vssd1 vccd1 vccd1 _13735_/Y sky130_fd_sc_hd__nand2_1
X_10947_ _20369_/Q _20433_/Q _11035_/S vssd1 vssd1 vccd1 vccd1 _10947_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_232_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19242_ _19523_/CLK _19242_/D vssd1 vssd1 vccd1 vccd1 _19242_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_220_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16454_ _16454_/A _16454_/B vssd1 vssd1 vccd1 vccd1 _17812_/A sky130_fd_sc_hd__nand2_4
XFILLER_231_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13666_ _13718_/A _13666_/B vssd1 vssd1 vccd1 vccd1 _13666_/Y sky130_fd_sc_hd__nor2_1
X_10878_ _11309_/A1 _10877_/X _10874_/X _12504_/A vssd1 vssd1 vccd1 vccd1 _10879_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_220_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15405_ _11773_/X _15127_/B _15404_/X vssd1 vssd1 vccd1 vccd1 _15405_/Y sky130_fd_sc_hd__o21ai_1
X_19173_ _20426_/CLK _19173_/D vssd1 vssd1 vccd1 vccd1 _19173_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12914_/B _12617_/B vssd1 vssd1 vccd1 vccd1 _12617_/Y sky130_fd_sc_hd__nand2_2
X_16385_ _19739_/Q _16386_/C _19740_/Q vssd1 vssd1 vccd1 vccd1 _16387_/B sky130_fd_sc_hd__a21oi_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _19661_/D _13595_/Y _13596_/X _13624_/B2 vssd1 vssd1 vccd1 vccd1 _13597_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18124_ _20783_/Q _18120_/B _18123_/Y vssd1 vssd1 vccd1 vccd1 _20783_/D sky130_fd_sc_hd__o21a_1
X_15336_ _20889_/Q _14971_/A _15323_/B _15335_/X _15478_/C1 vssd1 vssd1 vccd1 vccd1
+ _15336_/X sky130_fd_sc_hd__a221o_1
XFILLER_185_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12548_ _20868_/Q _12548_/B _12548_/C vssd1 vssd1 vccd1 vccd1 _12552_/D sky130_fd_sc_hd__and3_1
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18055_ _20758_/Q _18055_/B vssd1 vssd1 vccd1 vccd1 _18061_/C sky130_fd_sc_hd__and2_2
X_15267_ _15267_/A _15528_/B vssd1 vssd1 vccd1 vccd1 _15283_/B sky130_fd_sc_hd__nand2_1
XANTENNA_2 _19656_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12479_/A _12582_/C vssd1 vssd1 vccd1 vccd1 _12479_/X sky130_fd_sc_hd__and2_2
XFILLER_172_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17006_ _17006_/A1 _16049_/X _17003_/X _17005_/X vssd1 vssd1 vccd1 vccd1 _17006_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14218_ _19504_/Q _14218_/B vssd1 vssd1 vccd1 vccd1 _14219_/B sky130_fd_sc_hd__or2_1
X_15198_ _20789_/Q _16047_/A2 _15196_/X _15197_/X vssd1 vssd1 vccd1 vccd1 _15198_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14149_ _14161_/A _14160_/A vssd1 vssd1 vccd1 vccd1 _14151_/A sky130_fd_sc_hd__or2_1
Xfanout509 _17745_/X vssd1 vssd1 vccd1 vccd1 _17772_/S sky130_fd_sc_hd__buf_4
XFILLER_112_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18957_ _18675_/Y _18970_/A2 _18955_/Y _18956_/Y vssd1 vssd1 vccd1 vccd1 _18957_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17908_ _20679_/Q _17908_/A1 _17912_/S vssd1 vssd1 vccd1 vccd1 _20679_/D sky130_fd_sc_hd__mux2_1
X_09690_ _20356_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _09690_/X sky130_fd_sc_hd__or2_1
XFILLER_255_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18888_ _18636_/Y _18977_/A2 _18886_/Y _18887_/Y vssd1 vssd1 vccd1 vccd1 _18888_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1080 _12577_/X vssd1 vssd1 vccd1 vccd1 _15520_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_266_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1091 _12293_/X vssd1 vssd1 vccd1 vccd1 _17951_/A1 sky130_fd_sc_hd__buf_8
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17839_ _20614_/Q _17877_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20614_/D sky130_fd_sc_hd__mux2_1
XFILLER_66_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_255_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_254_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_254_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20850_ _20856_/CLK _20850_/D vssd1 vssd1 vccd1 vccd1 _20850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_270_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19509_ _20930_/CLK _19509_/D vssd1 vssd1 vccd1 vccd1 _19509_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20781_ _21043_/CLK _20781_/D vssd1 vssd1 vccd1 vccd1 _20781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_250_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20215_ _20763_/CLK _20215_/D vssd1 vssd1 vccd1 vccd1 _20215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_277_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20146_ _20641_/CLK _20146_/D vssd1 vssd1 vccd1 vccd1 _20146_/Q sky130_fd_sc_hd__dfxtp_1
X_09957_ _19885_/Q _19786_/Q _11979_/S vssd1 vssd1 vccd1 vccd1 _09957_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20077_ _20077_/CLK _20077_/D vssd1 vssd1 vccd1 vccd1 _20077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09886_/X _09887_/X _11904_/S vssd1 vssd1 vccd1 vccd1 _09888_/X sky130_fd_sc_hd__mux2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_258_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_246_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_261_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_403 _16911_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _11851_/A _20517_/Q _12165_/S _20549_/Q vssd1 vssd1 vccd1 vccd1 _11850_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_414 _18220_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_425 _10813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_154_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19970_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_272_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_436 _13716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ _13541_/A vssd1 vssd1 vccd1 vccd1 _10801_/Y sky130_fd_sc_hd__inv_2
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_447 _13755_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_458 _19107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11781_ _13482_/A _11781_/B vssd1 vssd1 vccd1 vccd1 _11786_/C sky130_fd_sc_hd__xnor2_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20979_ _21015_/CLK _20979_/D vssd1 vssd1 vccd1 vccd1 _20979_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_469 _19997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13520_ _18462_/A _13519_/X _13516_/X _18152_/B vssd1 vssd1 vccd1 vccd1 _13520_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_242_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10732_ _12371_/A1 _19340_/Q _20695_/Q _11074_/S _12371_/C1 vssd1 vssd1 vccd1 vccd1
+ _10732_/X sky130_fd_sc_hd__a221o_1
XFILLER_198_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13451_ _20925_/Q _13602_/A1 _13575_/C _13450_/Y _18612_/B vssd1 vssd1 vccd1 vccd1
+ _13451_/X sky130_fd_sc_hd__a221o_1
X_10663_ _12383_/A _10648_/Y _09502_/A vssd1 vssd1 vccd1 vccd1 _10663_/Y sky130_fd_sc_hd__a21oi_1
X_12402_ _12402_/A1 _17916_/A1 _12401_/X vssd1 vssd1 vccd1 vccd1 _12402_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16170_ _19609_/Q _15698_/X _16170_/S vssd1 vssd1 vccd1 vccd1 _16171_/B sky130_fd_sc_hd__mux2_1
X_10594_ _12073_/C1 _10586_/X _10593_/X _10570_/X _10579_/X vssd1 vssd1 vccd1 vccd1
+ _10594_/X sky130_fd_sc_hd__o32a_1
X_13382_ _13035_/Y _13382_/B vssd1 vssd1 vccd1 vccd1 _13383_/B sky130_fd_sc_hd__nand2b_1
XFILLER_182_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15121_ _15121_/A vssd1 vssd1 vccd1 vccd1 _15121_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12333_ _19829_/Q _12412_/A2 _12331_/X _09738_/A _12332_/X vssd1 vssd1 vccd1 vccd1
+ _12333_/X sky130_fd_sc_hd__o221a_1
XFILLER_127_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15052_ _14886_/X _15051_/X _15155_/S vssd1 vssd1 vccd1 vccd1 _15053_/A sky130_fd_sc_hd__mux2_1
X_12264_ _12420_/B1 _12262_/X _12263_/X vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__o21ai_1
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14003_ _19200_/Q _14081_/C _14003_/S vssd1 vssd1 vccd1 vccd1 _14003_/X sky130_fd_sc_hd__mux2_1
X_11215_ _11391_/A _20366_/Q _20430_/Q _12346_/S vssd1 vssd1 vccd1 vccd1 _11215_/X
+ sky130_fd_sc_hd__a22o_1
X_19860_ _20017_/CLK _19860_/D vssd1 vssd1 vccd1 vccd1 _19860_/Q sky130_fd_sc_hd__dfxtp_4
X_12195_ _19522_/Q _15960_/A _15895_/S vssd1 vssd1 vccd1 vccd1 _12198_/B sky130_fd_sc_hd__mux2_8
XFILLER_269_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18811_ _19501_/Q _18810_/X _18811_/S vssd1 vssd1 vccd1 vccd1 _18811_/X sky130_fd_sc_hd__mux2_1
X_11146_ _10385_/A _11145_/X _09613_/A vssd1 vssd1 vccd1 vccd1 _11146_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19791_ _20077_/CLK _19791_/D vssd1 vssd1 vccd1 vccd1 _19791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_284_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_283_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11077_ _11064_/X _11065_/X _12391_/S vssd1 vssd1 vccd1 vccd1 _11077_/X sky130_fd_sc_hd__mux2_1
XFILLER_249_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18742_ _18748_/A _18742_/B vssd1 vssd1 vccd1 vccd1 _20971_/D sky130_fd_sc_hd__and2_1
X_15954_ _15954_/A _15982_/C vssd1 vssd1 vccd1 vccd1 _15954_/Y sky130_fd_sc_hd__nand2_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput150 dout1[49] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__clkbuf_2
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput161 dout1[59] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__clkbuf_2
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905_ _12944_/C _19178_/Q _18149_/S vssd1 vssd1 vccd1 vccd1 _14950_/A sky130_fd_sc_hd__mux2_1
X_10028_ _10373_/A _11234_/B _10027_/X vssd1 vssd1 vccd1 vccd1 _10028_/X sky130_fd_sc_hd__or3b_2
Xinput172 irq[10] vssd1 vssd1 vccd1 vccd1 _12546_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_264_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18673_ _18980_/A _18673_/B vssd1 vssd1 vccd1 vccd1 _20941_/D sky130_fd_sc_hd__nor2_1
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput183 irq[6] vssd1 vssd1 vccd1 vccd1 _12545_/C sky130_fd_sc_hd__clkbuf_2
X_15885_ _16024_/A1 _15883_/X _15884_/Y _15976_/B2 vssd1 vssd1 vccd1 vccd1 _15885_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_236_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput194 localMemory_wb_adr_i[13] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_hd__clkbuf_2
XFILLER_264_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17624_ _20380_/Q _17935_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20380_/D sky130_fd_sc_hd__mux2_1
X_14836_ _11783_/B _14882_/A _14836_/S vssd1 vssd1 vccd1 vccd1 _14836_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ _20315_/Q _17691_/A1 _17570_/S vssd1 vssd1 vccd1 vccd1 _20315_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14767_ _19508_/Q _14773_/B vssd1 vssd1 vccd1 vccd1 _14767_/X sky130_fd_sc_hd__or2_1
X_11979_ _20392_/Q _20456_/Q _11979_/S vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16506_ _19813_/Q _17099_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19813_/D sky130_fd_sc_hd__mux2_1
XFILLER_205_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13718_ _13718_/A _13718_/B vssd1 vssd1 vccd1 vccd1 _13718_/Y sky130_fd_sc_hd__nand2_1
X_17486_ _20278_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17486_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14698_ _19457_/Q _17947_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19457_/D sky130_fd_sc_hd__mux2_1
XFILLER_108_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16437_ _19759_/Q _16437_/B vssd1 vssd1 vccd1 vccd1 _16442_/C sky130_fd_sc_hd__and2_2
X_19225_ _19505_/CLK _19225_/D vssd1 vssd1 vccd1 vccd1 _19225_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_258_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13649_ _13663_/A _13663_/B _13718_/B vssd1 vssd1 vccd1 vccd1 _13649_/X sky130_fd_sc_hd__and3_4
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19156_ _21044_/CLK _19156_/D vssd1 vssd1 vccd1 vccd1 _19156_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_176_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16368_ _19733_/Q _16370_/C _16367_/Y vssd1 vssd1 vccd1 vccd1 _19733_/D sky130_fd_sc_hd__o21a_1
X_18107_ _20777_/Q _18109_/C _18106_/Y vssd1 vssd1 vccd1 vccd1 _20777_/D sky130_fd_sc_hd__o21a_1
X_15319_ _17257_/A _14938_/Y _14979_/B _14980_/X _15318_/X vssd1 vssd1 vccd1 vccd1
+ _15319_/X sky130_fd_sc_hd__o311a_1
X_19087_ _19701_/CLK _19087_/D vssd1 vssd1 vccd1 vccd1 _19087_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16299_ _19707_/Q _16300_/C _16298_/Y vssd1 vssd1 vccd1 vccd1 _19707_/D sky130_fd_sc_hd__o21a_1
XFILLER_274_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18038_ _20751_/Q _18034_/B _18037_/Y vssd1 vssd1 vccd1 vccd1 _20751_/D sky130_fd_sc_hd__o21a_1
XFILLER_145_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_259_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20000_ _20624_/CLK _20000_/D vssd1 vssd1 vccd1 vccd1 _20000_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_141_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09811_ _20647_/Q _20611_/Q _12070_/S vssd1 vssd1 vccd1 vccd1 _09811_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19989_ _19992_/CLK _19989_/D vssd1 vssd1 vccd1 vccd1 _19989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_274_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ _12504_/A _13863_/A _17709_/C vssd1 vssd1 vccd1 vccd1 _09747_/C sky130_fd_sc_hd__and3_1
XFILLER_228_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09673_ _19854_/Q _19660_/Q _20019_/Q vssd1 vssd1 vccd1 vccd1 _09673_/X sky130_fd_sc_hd__or3b_4
XFILLER_67_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20902_ _21000_/CLK _20902_/D vssd1 vssd1 vccd1 vccd1 _20902_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20833_ _20962_/CLK _20833_/D vssd1 vssd1 vccd1 vccd1 _20833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_270_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20764_ _20795_/CLK _20764_/D vssd1 vssd1 vccd1 vccd1 _20764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_211_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20695_ _20718_/CLK _20695_/D vssd1 vssd1 vccd1 vccd1 _20695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11000_ _11273_/A1 _20496_/Q _10303_/S _20528_/Q vssd1 vssd1 vccd1 vccd1 _11000_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_278_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1816 _19181_/Q vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__buf_4
XFILLER_131_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_266_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1827 _10831_/S vssd1 vssd1 vccd1 vccd1 _11345_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout840 _18491_/B2 vssd1 vssd1 vccd1 vccd1 _18509_/B2 sky130_fd_sc_hd__buf_6
Xfanout1838 _11977_/A1 vssd1 vssd1 vccd1 vccd1 _11903_/A1 sky130_fd_sc_hd__buf_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1849 _19171_/Q vssd1 vssd1 vccd1 vccd1 _12584_/C sky130_fd_sc_hd__buf_12
Xfanout851 _18157_/Y vssd1 vssd1 vccd1 vccd1 _18316_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20129_ _20711_/CLK _20129_/D vssd1 vssd1 vccd1 vccd1 _20129_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout862 _15937_/C1 vssd1 vssd1 vccd1 vccd1 _16043_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout873 _14954_/X vssd1 vssd1 vccd1 vccd1 _15322_/A sky130_fd_sc_hd__buf_8
XFILLER_284_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout884 _14939_/Y vssd1 vssd1 vccd1 vccd1 _16048_/C1 sky130_fd_sc_hd__buf_6
XFILLER_19_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout895 _18395_/S vssd1 vssd1 vccd1 vccd1 _18419_/S sky130_fd_sc_hd__buf_4
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _18134_/A _16714_/C _16714_/B vssd1 vssd1 vccd1 vccd1 _16945_/C sky130_fd_sc_hd__nor3b_4
XFILLER_86_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_280_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_274_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_219_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _11887_/X _11888_/X _11902_/S vssd1 vssd1 vccd1 vccd1 _11902_/X sky130_fd_sc_hd__mux2_1
X_15670_ _19751_/Q _15942_/A2 _15669_/X _15999_/C1 vssd1 vssd1 vccd1 vccd1 _15670_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _16062_/B2 _12881_/X _12758_/B _19521_/Q vssd1 vssd1 vccd1 vccd1 _12883_/B
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA_200 _20424_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_273_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_211 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14621_ _19385_/Q _17871_/A1 _14630_/S vssd1 vssd1 vccd1 vccd1 _19385_/D sky130_fd_sc_hd__mux2_1
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11833_ _19647_/Q _11987_/S _11810_/X _11833_/C1 vssd1 vssd1 vccd1 vccd1 _11833_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_266 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_277 _20003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17340_ _20218_/Q _17364_/A2 _17370_/B1 _20267_/Q _17370_/C1 vssd1 vssd1 vccd1 vccd1
+ _17340_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14552_ _19322_/Q _17872_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19322_/D sky130_fd_sc_hd__mux2_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _13459_/A _11764_/B _15433_/A vssd1 vssd1 vccd1 vccd1 _11764_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_288 input219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_299 input227/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13503_ _13589_/A1 _13501_/X _13502_/Y _13500_/X vssd1 vssd1 vccd1 vccd1 _13507_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _20196_/Q _17280_/A2 _17270_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1 _20196_/D
+ sky130_fd_sc_hd__o211a_1
X_10715_ _12277_/A1 _17893_/A1 _10714_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _15331_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_42_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14483_ _20237_/Q _19266_/Q _14483_/S vssd1 vssd1 vccd1 vccd1 _14484_/B sky130_fd_sc_hd__mux2_1
X_11695_ _20319_/Q _11718_/S _12097_/S _10629_/A vssd1 vssd1 vccd1 vccd1 _11695_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_202_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19010_ _18220_/Y _18982_/B _19016_/B1 _19009_/X vssd1 vssd1 vccd1 vccd1 _21024_/D
+ sky130_fd_sc_hd__o211a_1
X_16222_ _19645_/Q _17874_/A1 _16227_/S vssd1 vssd1 vccd1 vccd1 _19645_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13434_ _13434_/A _13434_/B vssd1 vssd1 vccd1 vccd1 _15843_/A sky130_fd_sc_hd__xnor2_4
X_10646_ _12396_/A1 _19469_/Q _19437_/Q _12381_/S _12371_/C1 vssd1 vssd1 vccd1 vccd1
+ _10646_/X sky130_fd_sc_hd__a221o_1
XFILLER_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16153_ _19600_/Q _16178_/S _16152_/Y _16159_/C1 vssd1 vssd1 vccd1 vccd1 _19600_/D
+ sky130_fd_sc_hd__o211a_1
Xrebuffer5 _11408_/X vssd1 vssd1 vccd1 vccd1 _11409_/B sky130_fd_sc_hd__buf_2
XFILLER_6_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13365_ _19235_/Q _13365_/B vssd1 vssd1 vccd1 vccd1 _13365_/Y sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_51_wb_clk_i clkbuf_leaf_59_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _20468_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10577_ _11514_/A1 _12752_/A _19343_/Q _12059_/A1 vssd1 vssd1 vccd1 vccd1 _10577_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_177_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ _14828_/X _14835_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15104_/X sky130_fd_sc_hd__mux2_1
X_12316_ _19397_/Q _20688_/Q _12316_/S vssd1 vssd1 vccd1 vccd1 _12316_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16084_ _09657_/X _16126_/A2 _16083_/X vssd1 vssd1 vccd1 vccd1 _19566_/D sky130_fd_sc_hd__o21a_1
XFILLER_138_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ _19234_/Q _13296_/B vssd1 vssd1 vccd1 vccd1 _13296_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19912_ _20692_/CLK _19912_/D vssd1 vssd1 vccd1 vccd1 _19912_/Q sky130_fd_sc_hd__dfxtp_1
X_15035_ _14845_/X _14858_/X _15035_/S vssd1 vssd1 vccd1 vccd1 _15035_/X sky130_fd_sc_hd__mux2_2
X_12247_ _12517_/C _15922_/B2 _12246_/X vssd1 vssd1 vccd1 vccd1 _12282_/A sky130_fd_sc_hd__a21oi_4
XFILLER_244_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19843_ _20751_/CLK _19843_/D vssd1 vssd1 vccd1 vccd1 _19843_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _19295_/Q _20082_/Q _12188_/S vssd1 vssd1 vccd1 vccd1 _12178_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_268_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11129_ _11126_/X _11127_/X _11128_/X _12357_/A1 _11118_/A vssd1 vssd1 vccd1 vccd1
+ _11129_/X sky130_fd_sc_hd__a221o_1
X_19774_ _20718_/CLK _19774_/D vssd1 vssd1 vccd1 vccd1 _19774_/Q sky130_fd_sc_hd__dfxtp_1
X_16986_ _19989_/Q _17012_/A2 _16985_/Y _17998_/A vssd1 vssd1 vccd1 vccd1 _19989_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18725_ _20963_/Q _18245_/Y _18749_/S vssd1 vssd1 vccd1 vccd1 _18726_/B sky130_fd_sc_hd__mux2_1
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15937_ _20909_/Q _15937_/A2 _16043_/B1 _15936_/X _15937_/C1 vssd1 vssd1 vccd1 vccd1
+ _15937_/X sky130_fd_sc_hd__a221o_1
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_265_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_252_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15868_ _12058_/S _15978_/A2 _15980_/A2 vssd1 vssd1 vccd1 vccd1 _15868_/X sky130_fd_sc_hd__a21bo_1
X_18656_ _18535_/X _18684_/A2 _18654_/Y _18655_/Y vssd1 vssd1 vccd1 vccd1 _18657_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17607_ _17744_/A _17675_/B vssd1 vssd1 vccd1 vccd1 _17608_/C sky130_fd_sc_hd__nor2_1
X_14819_ _11799_/B _11404_/B _14822_/S vssd1 vssd1 vccd1 vccd1 _14819_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18587_ _18814_/A _18587_/B vssd1 vssd1 vccd1 vccd1 _20919_/D sky130_fd_sc_hd__nor2_1
X_15799_ _20872_/Q _16018_/A2 fanout818/X vssd1 vssd1 vccd1 vccd1 _15799_/X sky130_fd_sc_hd__o21ba_1
XFILLER_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_251_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17538_ _19095_/Q _19093_/Q _17538_/C vssd1 vssd1 vccd1 vccd1 _17675_/B sky130_fd_sc_hd__or3_2
XFILLER_189_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17469_ _17495_/A1 _17468_/Y _18795_/A vssd1 vssd1 vccd1 vccd1 _20269_/D sky130_fd_sc_hd__a21oi_1
XFILLER_60_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19208_ _19590_/CLK _19208_/D vssd1 vssd1 vccd1 vccd1 _19208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20480_ _20480_/CLK _20480_/D vssd1 vssd1 vccd1 vccd1 _20480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19139_ _20300_/CLK _19139_/D vssd1 vssd1 vccd1 vccd1 _19139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_285_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_218_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput410 _19961_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[0] sky130_fd_sc_hd__buf_4
Xoutput421 _19962_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[1] sky130_fd_sc_hd__buf_4
XFILLER_145_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput432 _19963_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[2] sky130_fd_sc_hd__buf_4
XFILLER_218_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput443 _18949_/B1 vssd1 vssd1 vccd1 vccd1 probe_env[0] sky130_fd_sc_hd__buf_4
XFILLER_271_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput454 _19507_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[13] sky130_fd_sc_hd__buf_4
Xoutput465 _19517_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[23] sky130_fd_sc_hd__buf_4
X_21032_ _21041_/CLK _21032_/D vssd1 vssd1 vccd1 vccd1 _21032_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput476 _19498_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[4] sky130_fd_sc_hd__buf_4
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput487 _13826_/X vssd1 vssd1 vccd1 vccd1 wmask0[3] sky130_fd_sc_hd__buf_6
XFILLER_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09725_ _12157_/A1 _17909_/A1 _12153_/B1 _09724_/X vssd1 vssd1 vccd1 vccd1 _13734_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09656_ input168/X input139/X _11241_/S vssd1 vssd1 vccd1 vccd1 _09656_/X sky130_fd_sc_hd__mux2_8
XFILLER_28_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_271_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09587_ _14112_/A _19088_/Q _19089_/Q _19090_/Q vssd1 vssd1 vccd1 vccd1 _09592_/B
+ sky130_fd_sc_hd__and4bb_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20816_ _20816_/CLK _20816_/D vssd1 vssd1 vccd1 vccd1 _20816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20747_ _20812_/CLK _20747_/D vssd1 vssd1 vccd1 vccd1 _20747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_184_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ _11266_/A1 _19907_/Q _10324_/S _20032_/Q vssd1 vssd1 vccd1 vccd1 _10500_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11480_ _20542_/Q _20510_/Q _12165_/S vssd1 vssd1 vccd1 vccd1 _11480_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20678_ _20678_/CLK _20678_/D vssd1 vssd1 vccd1 vccd1 _20678_/Q sky130_fd_sc_hd__dfxtp_1
X_10431_ _10421_/X _10424_/X _10427_/X _10430_/X _12058_/S _12059_/A1 vssd1 vssd1
+ vccd1 vccd1 _10431_/X sky130_fd_sc_hd__mux4_2
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13150_ _13150_/A _13150_/B vssd1 vssd1 vccd1 vccd1 _13567_/B sky130_fd_sc_hd__nand2_2
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ _12433_/A1 _17866_/A1 _10361_/X _12433_/B2 vssd1 vssd1 vccd1 vccd1 _15561_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12101_ _20327_/Q _11708_/B _12100_/X vssd1 vssd1 vccd1 vccd1 _12101_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10293_ _10385_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10293_/Y sky130_fd_sc_hd__nand2_1
X_13081_ _13270_/A _13270_/C _13270_/B vssd1 vssd1 vccd1 vccd1 _13395_/A sky130_fd_sc_hd__a21boi_4
XFILLER_151_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ _19521_/Q _12031_/Y _15949_/A vssd1 vssd1 vccd1 vccd1 _12035_/B sky130_fd_sc_hd__mux2_8
XFILLER_278_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1602 _11995_/S vssd1 vssd1 vccd1 vccd1 _12071_/S sky130_fd_sc_hd__buf_6
Xfanout1613 fanout1630/X vssd1 vssd1 vccd1 vccd1 _11513_/S sky130_fd_sc_hd__buf_6
XFILLER_132_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1624 _12376_/S vssd1 vssd1 vccd1 vccd1 _12391_/S sky130_fd_sc_hd__buf_6
XFILLER_239_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1635 _09614_/X vssd1 vssd1 vccd1 vccd1 _12152_/A1 sky130_fd_sc_hd__buf_8
X_16840_ _16876_/A _16840_/B vssd1 vssd1 vccd1 vccd1 _16840_/Y sky130_fd_sc_hd__nor2_1
Xfanout1646 _12532_/X vssd1 vssd1 vccd1 vccd1 _18949_/A2 sky130_fd_sc_hd__buf_8
Xfanout1657 _11228_/B1 vssd1 vssd1 vccd1 vccd1 _11242_/B1 sky130_fd_sc_hd__buf_4
Xfanout670 _13943_/S vssd1 vssd1 vccd1 vccd1 _13941_/B sky130_fd_sc_hd__buf_6
Xfanout1668 _09532_/X vssd1 vssd1 vccd1 vccd1 _14112_/B sky130_fd_sc_hd__buf_12
Xfanout681 _13986_/A2 vssd1 vssd1 vccd1 vccd1 _14004_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout1679 _12007_/A1 vssd1 vssd1 vccd1 vccd1 _09752_/A sky130_fd_sc_hd__buf_6
X_16771_ _16726_/X _16770_/Y _16886_/B2 vssd1 vssd1 vccd1 vccd1 _16771_/X sky130_fd_sc_hd__a21o_2
Xfanout692 split9/A vssd1 vssd1 vccd1 vccd1 _13816_/B1 sky130_fd_sc_hd__buf_4
X_13983_ _19161_/Q _13986_/A2 _14004_/B1 _13982_/X _14070_/C1 vssd1 vssd1 vccd1 vccd1
+ _19161_/D sky130_fd_sc_hd__o221a_1
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_265_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15722_ _16017_/C1 _15721_/X _15717_/X vssd1 vssd1 vccd1 vccd1 _15722_/X sky130_fd_sc_hd__o21a_1
X_18510_ _18856_/A _18510_/B vssd1 vssd1 vccd1 vccd1 _20896_/D sky130_fd_sc_hd__nor2_1
XFILLER_218_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12934_ _16720_/A vssd1 vssd1 vccd1 vccd1 _12946_/B sky130_fd_sc_hd__inv_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19490_ _20677_/CLK _19490_/D vssd1 vssd1 vccd1 vccd1 _19490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18441_ _20875_/Q _18285_/Y _18453_/S vssd1 vssd1 vccd1 vccd1 _18442_/B sky130_fd_sc_hd__mux2_1
X_15653_ _13427_/B _15982_/C _16056_/B1 vssd1 vssd1 vccd1 vccd1 _15653_/X sky130_fd_sc_hd__a21o_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12865_ _13248_/A _13321_/B _12864_/Y vssd1 vssd1 vccd1 vccd1 _12866_/B sky130_fd_sc_hd__o21ai_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _19368_/Q _17888_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19368_/D sky130_fd_sc_hd__mux2_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18372_ _20841_/Q _18375_/B _18371_/Y _18748_/A vssd1 vssd1 vccd1 vccd1 _20841_/D
+ sky130_fd_sc_hd__o211a_1
X_11816_ _20389_/Q _20453_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _11816_/X sky130_fd_sc_hd__mux2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15468_/A _15578_/X _15581_/X vssd1 vssd1 vccd1 vccd1 _15584_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12517_/B split6/X _12771_/B _12767_/X _12759_/X vssd1 vssd1 vccd1 vccd1
+ _12796_/X sky130_fd_sc_hd__a41o_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ input6/X _15081_/A _17329_/S vssd1 vssd1 vccd1 vccd1 _17323_/X sky130_fd_sc_hd__mux2_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14535_ _19305_/Q _17855_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19305_/D sky130_fd_sc_hd__mux2_1
XFILLER_159_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _09859_/X _15789_/A vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__and2b_2
XFILLER_159_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17254_ _17254_/A _17275_/B _17269_/C vssd1 vssd1 vccd1 vccd1 _17254_/X sky130_fd_sc_hd__and3_1
XFILLER_186_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14466_ _18700_/A _14466_/B vssd1 vssd1 vccd1 vccd1 _19257_/D sky130_fd_sc_hd__and2_1
X_11678_ _19641_/Q _11682_/S _11655_/X _11995_/S vssd1 vssd1 vccd1 vccd1 _11678_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16205_ _19628_/Q _17751_/A1 _16230_/S vssd1 vssd1 vccd1 vccd1 _19628_/D sky130_fd_sc_hd__mux2_1
XFILLER_30_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13417_ _13417_/A vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__clkinv_2
XFILLER_174_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17185_ _17745_/A _17676_/B _17185_/C vssd1 vssd1 vccd1 vccd1 _17185_/X sky130_fd_sc_hd__and3_2
X_10629_ _10629_/A _10629_/B vssd1 vssd1 vccd1 vccd1 _10629_/X sky130_fd_sc_hd__or2_1
XFILLER_190_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14397_ _14397_/A _14397_/B _14397_/C vssd1 vssd1 vccd1 vccd1 _14397_/X sky130_fd_sc_hd__or3_1
XFILLER_128_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16136_ _16732_/B _16196_/S vssd1 vssd1 vccd1 vccd1 _16136_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13348_ _12664_/C _13347_/Y _13334_/A vssd1 vssd1 vccd1 vccd1 _13352_/A sky130_fd_sc_hd__a21o_1
XFILLER_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16067_ _14524_/A1 _16133_/A _16068_/A _16068_/C vssd1 vssd1 vccd1 vccd1 _16067_/X
+ sky130_fd_sc_hd__and4bb_4
X_13279_ _13279_/A _13279_/B vssd1 vssd1 vccd1 vccd1 _13309_/B sky130_fd_sc_hd__or2_1
XFILLER_142_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15018_ _15314_/D _15018_/B vssd1 vssd1 vccd1 vccd1 _15018_/X sky130_fd_sc_hd__and2b_1
XFILLER_69_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_271_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_257_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19826_ _20075_/CLK _19826_/D vssd1 vssd1 vccd1 vccd1 _19826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_284_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19757_ _20742_/CLK _19757_/D vssd1 vssd1 vccd1 vccd1 _19757_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_284_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16969_ _16966_/Y _16968_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16969_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_77_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09510_ _19093_/Q vssd1 vssd1 vccd1 vccd1 _16243_/B sky130_fd_sc_hd__inv_2
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18708_ _18708_/A _18708_/B vssd1 vssd1 vccd1 vccd1 _20954_/D sky130_fd_sc_hd__and2_1
XFILLER_237_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19688_ _20579_/CLK _19688_/D vssd1 vssd1 vccd1 vccd1 _19688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18639_ _20933_/Q _18686_/B vssd1 vssd1 vccd1 vccd1 _18639_/Y sky130_fd_sc_hd__nand2_1
XFILLER_213_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20601_ _20668_/CLK _20601_/D vssd1 vssd1 vccd1 vccd1 _20601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20532_ _20664_/CLK _20532_/D vssd1 vssd1 vccd1 vccd1 _20532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20463_ _20463_/CLK _20463_/D vssd1 vssd1 vccd1 vccd1 _20463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20394_ _20491_/CLK _20394_/D vssd1 vssd1 vccd1 vccd1 _20394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput295 _13782_/X vssd1 vssd1 vccd1 vccd1 addr1[1] sky130_fd_sc_hd__buf_4
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21015_ _21015_/CLK _21015_/D vssd1 vssd1 vccd1 vccd1 _21015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09708_ _09706_/X _09707_/X _11904_/S vssd1 vssd1 vccd1 vccd1 _09708_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10980_ _20464_/Q _12213_/B _10235_/S vssd1 vssd1 vccd1 vccd1 _10980_/X sky130_fd_sc_hd__a21o_1
XFILLER_215_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _11235_/A _10020_/B _09610_/C vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__a21bo_1
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12650_ _12648_/X _12649_/Y _12752_/B vssd1 vssd1 vccd1 vccd1 _12653_/A sky130_fd_sc_hd__a21oi_2
XFILLER_215_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11601_ _19642_/Q _11965_/B _11586_/X _11528_/S vssd1 vssd1 vccd1 vccd1 _11601_/X
+ sky130_fd_sc_hd__o211a_1
X_12581_ _12581_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12583_/B sky130_fd_sc_hd__or2_2
XFILLER_157_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14320_ _20286_/Q _14330_/A2 _14330_/B1 input227/X vssd1 vssd1 vccd1 vccd1 _14322_/B
+ sky130_fd_sc_hd__a22o_4
X_11532_ _12039_/A1 _11243_/X split7/X vssd1 vssd1 vccd1 vccd1 _11532_/X sky130_fd_sc_hd__a21o_4
XFILLER_278_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14251_ _14250_/A _14250_/B _14250_/C vssd1 vssd1 vccd1 vccd1 _14260_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_278_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11463_ _19882_/Q _19783_/Q _12185_/S vssd1 vssd1 vccd1 vccd1 _11464_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13202_ _13231_/B _13201_/Y _13334_/A vssd1 vssd1 vccd1 vccd1 _13202_/X sky130_fd_sc_hd__o21a_1
XFILLER_183_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10414_ _10412_/X _10413_/X _12082_/S vssd1 vssd1 vccd1 vccd1 _10414_/X sky130_fd_sc_hd__mux2_1
X_14182_ _14202_/S _14182_/B vssd1 vssd1 vccd1 vccd1 _14182_/Y sky130_fd_sc_hd__nand2_1
XFILLER_152_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11394_ _11392_/X _11393_/X _12340_/S vssd1 vssd1 vccd1 vccd1 _11394_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13133_ _13128_/X _13131_/X _13132_/Y vssd1 vssd1 vccd1 vccd1 _13133_/Y sky130_fd_sc_hd__o21ai_1
X_10345_ _20132_/Q _20100_/Q _10345_/S vssd1 vssd1 vccd1 vccd1 _10345_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18990_ _18170_/Y _18983_/B _19002_/B1 _18989_/X vssd1 vssd1 vccd1 vccd1 _21014_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _13064_/A _13064_/B _13064_/C _13064_/D vssd1 vssd1 vccd1 vccd1 _13064_/X
+ sky130_fd_sc_hd__and4_2
X_17941_ _20710_/Q _17941_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20710_/D sky130_fd_sc_hd__mux2_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_239_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10276_ _15613_/S vssd1 vssd1 vccd1 vccd1 _10276_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_279_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1410 _10174_/S vssd1 vssd1 vccd1 vccd1 _11035_/S sky130_fd_sc_hd__buf_6
X_12015_ _12015_/A1 _12013_/X _12014_/X vssd1 vssd1 vccd1 vccd1 _12015_/Y sky130_fd_sc_hd__o21ai_1
Xfanout1421 fanout1422/X vssd1 vssd1 vccd1 vccd1 _12272_/B2 sky130_fd_sc_hd__buf_6
X_17872_ _20645_/Q _17872_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20645_/D sky130_fd_sc_hd__mux2_1
Xfanout1432 _12190_/C1 vssd1 vssd1 vccd1 vccd1 _11641_/S sky130_fd_sc_hd__buf_6
XFILLER_266_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1443 _09986_/C vssd1 vssd1 vccd1 vccd1 _12008_/C sky130_fd_sc_hd__clkbuf_4
Xfanout1454 _09734_/Y vssd1 vssd1 vccd1 vccd1 _11191_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19611_ _20263_/CLK _19611_/D vssd1 vssd1 vccd1 vccd1 _19611_/Q sky130_fd_sc_hd__dfxtp_1
X_16823_ _19970_/Q _16707_/X _16822_/Y _18821_/A vssd1 vssd1 vccd1 vccd1 _19970_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1465 _11204_/S vssd1 vssd1 vccd1 vccd1 _12006_/S sky130_fd_sc_hd__buf_8
XFILLER_93_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1476 _11204_/S vssd1 vssd1 vccd1 vccd1 _12414_/S sky130_fd_sc_hd__buf_12
Xfanout1487 _11396_/S vssd1 vssd1 vccd1 vccd1 _12275_/A sky130_fd_sc_hd__buf_12
XFILLER_65_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1498 _11169_/B vssd1 vssd1 vccd1 vccd1 _09688_/B sky130_fd_sc_hd__buf_6
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19542_ _19607_/CLK _19542_/D vssd1 vssd1 vccd1 vccd1 _19542_/Q sky130_fd_sc_hd__dfxtp_4
X_13966_ _14002_/A1 _13969_/A2 _10724_/X _14002_/B1 _19837_/Q vssd1 vssd1 vccd1 vccd1
+ _14057_/C sky130_fd_sc_hd__o32a_1
X_16754_ _16869_/A _16754_/B vssd1 vssd1 vccd1 vccd1 _16754_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_234_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12917_ _12917_/A _12917_/B vssd1 vssd1 vccd1 vccd1 _12917_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_74_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15705_ _15705_/A _15705_/B _16007_/A vssd1 vssd1 vccd1 vccd1 _15705_/X sky130_fd_sc_hd__or3b_1
X_19473_ _20711_/CLK _19473_/D vssd1 vssd1 vccd1 vccd1 _19473_/Q sky130_fd_sc_hd__dfxtp_1
X_16685_ _19940_/Q _17095_/A1 _16701_/S vssd1 vssd1 vccd1 vccd1 _19940_/D sky130_fd_sc_hd__mux2_1
X_13897_ _13897_/A _14112_/B _14527_/A2 vssd1 vssd1 vccd1 vccd1 _13897_/X sky130_fd_sc_hd__or3b_1
XFILLER_234_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ _18724_/A _18424_/B vssd1 vssd1 vccd1 vccd1 _20866_/D sky130_fd_sc_hd__and2_1
XFILLER_221_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12848_ _12843_/X _12847_/X _15703_/B2 vssd1 vssd1 vccd1 vccd1 _12852_/A sky130_fd_sc_hd__a21o_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15636_ _20898_/Q _15937_/A2 _15994_/B1 _15635_/X _15937_/C1 vssd1 vssd1 vccd1 vccd1
+ _15636_/X sky130_fd_sc_hd__a221o_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18355_ _18511_/B _18357_/B vssd1 vssd1 vccd1 vccd1 _18355_/Y sky130_fd_sc_hd__nand2_1
X_15567_ _20928_/Q _15567_/A2 _15566_/X vssd1 vssd1 vccd1 vccd1 _15567_/X sky130_fd_sc_hd__o21a_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _11367_/A _13589_/A1 _12776_/Y _12777_/X vssd1 vssd1 vccd1 vccd1 _12790_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_148_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17306_ _20207_/Q _17321_/A2 _17324_/C1 vssd1 vssd1 vccd1 vccd1 _17306_/X sky130_fd_sc_hd__a21o_1
X_14518_ _19296_/Q _17915_/A1 _14520_/S vssd1 vssd1 vccd1 vccd1 _19296_/D sky130_fd_sc_hd__mux2_1
XFILLER_203_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_230_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18286_ _20811_/Q _18285_/Y _18296_/S vssd1 vssd1 vccd1 vccd1 _18287_/B sky130_fd_sc_hd__mux2_1
X_15498_ _15612_/S _15181_/X _15497_/X vssd1 vssd1 vccd1 vccd1 _15498_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_266_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17237_ _17236_/A _17321_/A2 _17302_/C _20259_/Q _17291_/B1 vssd1 vssd1 vccd1 vccd1
+ _17237_/X sky130_fd_sc_hd__a221o_1
X_14449_ _20220_/Q _19249_/Q _14477_/S vssd1 vssd1 vccd1 vccd1 _14450_/B sky130_fd_sc_hd__mux2_1
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17168_ _20134_/Q _17202_/A1 _17180_/S vssd1 vssd1 vccd1 vccd1 _20134_/D sky130_fd_sc_hd__mux2_1
XFILLER_115_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16119_ _19584_/Q _16127_/A2 _16127_/B1 vssd1 vssd1 vccd1 vccd1 _16119_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17099_ _20069_/Q _17099_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20069_/D sky130_fd_sc_hd__mux2_1
XFILLER_170_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ _12008_/A _20513_/Q _12185_/S _20545_/Q vssd1 vssd1 vccd1 vccd1 _09990_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19809_ _20539_/CLK _19809_/D vssd1 vssd1 vccd1 vccd1 _19809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_285_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_244_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_253_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20515_ _20679_/CLK _20515_/D vssd1 vssd1 vccd1 vccd1 _20515_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_179_wb_clk_i clkbuf_4_4__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20291_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20446_ _20446_/CLK _20446_/D vssd1 vssd1 vccd1 vccd1 _20446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_108_wb_clk_i clkbuf_4_15__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20796_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_238_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_279_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20377_ _20451_/CLK _20377_/D vssd1 vssd1 vccd1 vccd1 _20377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10130_ _11258_/A1 _19347_/Q _20702_/Q _10217_/S _11338_/A1 vssd1 vssd1 vccd1 vccd1
+ _10130_/X sky130_fd_sc_hd__a221o_1
XFILLER_161_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10061_ _20345_/Q _11680_/C1 _12044_/B _12071_/S vssd1 vssd1 vccd1 vccd1 _10061_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13820_ _13822_/A1 _13770_/B split9/X input236/X vssd1 vssd1 vccd1 vccd1 _13820_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_217_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ _12075_/Y _13730_/B _13776_/B1 vssd1 vssd1 vccd1 vccd1 _13754_/A sky130_fd_sc_hd__o21a_2
XFILLER_250_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10963_ _12275_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10963_/Y sky130_fd_sc_hd__nor2_1
XFILLER_216_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12702_ _19509_/Q _12718_/A vssd1 vssd1 vccd1 vccd1 _12703_/B sky130_fd_sc_hd__nor2_1
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16470_ _19779_/Q _17933_/A1 _16488_/S vssd1 vssd1 vccd1 vccd1 _19779_/D sky130_fd_sc_hd__mux2_1
XFILLER_245_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13682_ _13718_/A _13680_/Y _13681_/Y _13655_/A vssd1 vssd1 vccd1 vccd1 _13683_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_243_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10894_ _10127_/A _10889_/Y _10893_/X _10887_/X vssd1 vssd1 vccd1 vccd1 _10894_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15421_ _17299_/A _15482_/A2 _15016_/A _20795_/Q _15420_/X vssd1 vssd1 vccd1 vccd1
+ _15421_/X sky130_fd_sc_hd__a221o_1
XFILLER_232_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12633_ _12631_/X _12632_/Y _12752_/B vssd1 vssd1 vccd1 vccd1 _12633_/Y sky130_fd_sc_hd__a21oi_2
XPHY_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18140_ _12944_/A _19110_/Q _18148_/S vssd1 vssd1 vccd1 vccd1 _18389_/A sky130_fd_sc_hd__mux2_2
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15352_ _15155_/X _15161_/A _15357_/S vssd1 vssd1 vccd1 vccd1 _15352_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12564_ _13658_/A _13740_/B vssd1 vssd1 vccd1 vccd1 _13714_/S sky130_fd_sc_hd__or2_4
XFILLER_129_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14303_ _14303_/A _14303_/B vssd1 vssd1 vccd1 vccd1 _14304_/B sky130_fd_sc_hd__nor2_1
X_18071_ _20764_/Q _18071_/B vssd1 vssd1 vccd1 vccd1 _18077_/C sky130_fd_sc_hd__and2_2
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11515_ _11513_/X _11514_/X _12135_/A vssd1 vssd1 vccd1 vccd1 _11515_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15283_ _15283_/A _15283_/B vssd1 vssd1 vccd1 vccd1 _15283_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12495_ _12496_/A _12496_/B vssd1 vssd1 vccd1 vccd1 _12495_/Y sky130_fd_sc_hd__nand2_1
XFILLER_200_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17022_ _20000_/Q input209/X _17026_/S vssd1 vssd1 vccd1 vccd1 _20000_/D sky130_fd_sc_hd__mux2_1
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14234_ _14244_/A1 _14233_/X _13457_/X vssd1 vssd1 vccd1 vccd1 _14235_/C sky130_fd_sc_hd__o21ba_1
XFILLER_172_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11446_ _20039_/Q _19914_/Q _12139_/S vssd1 vssd1 vccd1 vccd1 _11446_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14165_ _14255_/A _14204_/B _14165_/C vssd1 vssd1 vccd1 vccd1 _14165_/X sky130_fd_sc_hd__or3_1
XFILLER_166_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11377_ _19873_/Q _19774_/Q _11377_/S vssd1 vssd1 vccd1 vccd1 _11377_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ _13116_/A _13116_/B _13116_/C vssd1 vssd1 vccd1 vccd1 _13116_/Y sky130_fd_sc_hd__nand3_1
X_10328_ _11012_/A _10327_/X _13675_/A vssd1 vssd1 vccd1 vccd1 _10328_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14096_ _19207_/Q _14108_/A2 _14095_/X _16127_/B1 vssd1 vssd1 vccd1 vccd1 _19207_/D
+ sky130_fd_sc_hd__o211a_1
X_18973_ _18973_/A _18973_/B vssd1 vssd1 vccd1 vccd1 _21010_/D sky130_fd_sc_hd__nor2_1
XFILLER_113_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17924_ _20693_/Q _17924_/A1 _17934_/S vssd1 vssd1 vccd1 vccd1 _20693_/D sky130_fd_sc_hd__mux2_1
X_13047_ _20954_/Q _20888_/Q vssd1 vssd1 vccd1 vccd1 _13047_/X sky130_fd_sc_hd__or2_2
X_10259_ _11375_/S _10254_/X _10258_/X vssd1 vssd1 vccd1 vccd1 _10259_/X sky130_fd_sc_hd__o21a_1
XFILLER_140_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_252_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1240 _09596_/X vssd1 vssd1 vccd1 vccd1 _12365_/A2 sky130_fd_sc_hd__buf_8
XFILLER_61_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1251 _17335_/X vssd1 vssd1 vccd1 vccd1 _17381_/A2 sky130_fd_sc_hd__buf_6
X_17855_ _20628_/Q _17855_/A1 _17883_/S vssd1 vssd1 vccd1 vccd1 _20628_/D sky130_fd_sc_hd__mux2_1
XFILLER_38_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1262 _12477_/X vssd1 vssd1 vccd1 vccd1 _12730_/A2 sky130_fd_sc_hd__buf_4
XFILLER_266_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1273 _15303_/A vssd1 vssd1 vccd1 vccd1 _16052_/B2 sky130_fd_sc_hd__clkbuf_4
XFILLER_267_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1284 _09547_/X vssd1 vssd1 vccd1 vccd1 _10935_/B sky130_fd_sc_hd__buf_4
X_16806_ _20405_/Q _16870_/A2 _16870_/B1 vssd1 vssd1 vccd1 vccd1 _16806_/X sky130_fd_sc_hd__a21o_2
Xfanout1295 _12752_/B vssd1 vssd1 vccd1 vccd1 _12716_/B sky130_fd_sc_hd__buf_6
XFILLER_281_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17786_ _20563_/Q _17926_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20563_/D sky130_fd_sc_hd__mux2_1
X_14998_ _20946_/Q _14972_/B _14997_/X _20818_/Q _15322_/B vssd1 vssd1 vccd1 vccd1
+ _14998_/X sky130_fd_sc_hd__a221o_1
XFILLER_226_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_281_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19525_ _20300_/CLK _19525_/D vssd1 vssd1 vccd1 vccd1 _19525_/Q sky130_fd_sc_hd__dfxtp_4
X_16737_ _16735_/X _16736_/X _12930_/B vssd1 vssd1 vccd1 vccd1 _16737_/X sky130_fd_sc_hd__a21bo_1
X_13949_ _19182_/Q _14045_/C _14003_/S vssd1 vssd1 vccd1 vccd1 _13949_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19456_ _20583_/CLK _19456_/D vssd1 vssd1 vccd1 vccd1 _19456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16668_ _19925_/Q _17112_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19925_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18407_ _20858_/Q _18200_/Y _18419_/S vssd1 vssd1 vccd1 vccd1 _18408_/B sky130_fd_sc_hd__mux2_1
XFILLER_222_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15619_ _15616_/X _15618_/X _15703_/B2 vssd1 vssd1 vccd1 vccd1 _15619_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_222_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19387_ _20678_/CLK _19387_/D vssd1 vssd1 vccd1 vccd1 _19387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_250_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16599_ _16596_/X _16598_/X _16567_/A vssd1 vssd1 vccd1 vccd1 _16599_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_277_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18338_ _20824_/Q _18343_/B _18337_/Y _18692_/A vssd1 vssd1 vccd1 vccd1 _20824_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_194_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19956_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_187_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18269_ _18299_/A1 _14342_/B _18268_/Y vssd1 vssd1 vccd1 vccd1 _18532_/B sky130_fd_sc_hd__o21ai_4
XFILLER_147_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20300_ _20300_/CLK _20300_/D vssd1 vssd1 vccd1 vccd1 _20300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_201_wb_clk_i _19552_/CLK vssd1 vssd1 vccd1 vccd1 _20646_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20231_ _20621_/CLK _20231_/D vssd1 vssd1 vccd1 vccd1 _20231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20162_ _20711_/CLK _20162_/D vssd1 vssd1 vccd1 vccd1 _20162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_277_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09973_ _19643_/Q _12124_/S _09950_/X _11833_/C1 vssd1 vssd1 vccd1 vccd1 _09973_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20093_ _20719_/CLK _20093_/D vssd1 vssd1 vccd1 vccd1 _20093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_245_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_607 _20624_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_618 _13775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_629 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20995_ _21027_/CLK _20995_/D vssd1 vssd1 vccd1 vccd1 _20995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_253_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_213_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11300_ _09507_/A _11298_/X _11299_/X vssd1 vssd1 vccd1 vccd1 _11300_/X sky130_fd_sc_hd__o21a_1
XFILLER_267_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ _12282_/A _12282_/B vssd1 vssd1 vccd1 vccd1 _12283_/A sky130_fd_sc_hd__nor2_4
XFILLER_119_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11231_ input169/X input141/X _11241_/S vssd1 vssd1 vccd1 vccd1 _11231_/X sky130_fd_sc_hd__mux2_8
X_20429_ _21047_/A _20429_/D vssd1 vssd1 vccd1 vccd1 _20429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11162_ _11268_/A _20626_/Q _20590_/Q _12295_/B _12318_/A1 vssd1 vssd1 vccd1 vccd1
+ _11162_/X sky130_fd_sc_hd__o221a_1
XFILLER_162_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _10113_/A _15500_/S vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__nand2_4
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11093_ _19269_/Q _20056_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _11093_/X sky130_fd_sc_hd__mux2_1
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ _20814_/Q _15998_/A2 _15963_/X _16000_/A1 _15969_/X vssd1 vssd1 vccd1 vccd1
+ _15970_/X sky130_fd_sc_hd__a221o_1
XFILLER_267_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xsplit6 split6/A vssd1 vssd1 vccd1 vccd1 split6/X sky130_fd_sc_hd__clkbuf_4
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14921_ _18148_/S _14921_/B vssd1 vssd1 vccd1 vccd1 _14921_/X sky130_fd_sc_hd__and2b_1
X_10044_ _10385_/A _10044_/B vssd1 vssd1 vccd1 vccd1 _10044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_76_wb_clk_i clkbuf_4_9__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20638_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17640_ _20396_/Q _17708_/A1 _17640_/S vssd1 vssd1 vccd1 vccd1 _20396_/D sky130_fd_sc_hd__mux2_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14852_ _11412_/B _11737_/B _14853_/S vssd1 vssd1 vccd1 vccd1 _14852_/X sky130_fd_sc_hd__mux2_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13803_ _13822_/A1 _13687_/B _13790_/X input218/X vssd1 vssd1 vccd1 vccd1 _13803_/X
+ sky130_fd_sc_hd__a22o_1
X_17571_ _20331_/Q _17707_/A1 _17572_/S vssd1 vssd1 vccd1 vccd1 _20331_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14783_ _19516_/Q _14801_/B vssd1 vssd1 vccd1 vccd1 _14783_/X sky130_fd_sc_hd__or2_1
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11995_ _11993_/X _11994_/X _11995_/S vssd1 vssd1 vccd1 vccd1 _11995_/X sky130_fd_sc_hd__mux2_1
XFILLER_189_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19310_ _20658_/CLK _19310_/D vssd1 vssd1 vccd1 vccd1 _19310_/Q sky130_fd_sc_hd__dfxtp_1
X_16522_ _19829_/Q _17674_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19829_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13734_ _13734_/A _13742_/B vssd1 vssd1 vccd1 vccd1 _13777_/B sky130_fd_sc_hd__or2_4
X_10946_ _10940_/X _10945_/X _12258_/S vssd1 vssd1 vccd1 vccd1 _10946_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19241_ _19520_/CLK _19241_/D vssd1 vssd1 vccd1 vccd1 _19241_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16453_ _19765_/Q _16451_/C _16452_/Y vssd1 vssd1 vccd1 vccd1 _19765_/D sky130_fd_sc_hd__o21a_1
X_13665_ _13665_/A vssd1 vssd1 vccd1 vccd1 _13665_/Y sky130_fd_sc_hd__inv_2
X_10877_ _09731_/A _10876_/X _10875_/X vssd1 vssd1 vccd1 vccd1 _10877_/X sky130_fd_sc_hd__o21a_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ _19524_/Q _12624_/A vssd1 vssd1 vccd1 vccd1 _12617_/B sky130_fd_sc_hd__or2_1
X_15404_ _13596_/X _15494_/B _12579_/D vssd1 vssd1 vccd1 vccd1 _15404_/X sky130_fd_sc_hd__o21a_1
X_16384_ _19739_/Q _16386_/C _16383_/Y vssd1 vssd1 vccd1 vccd1 _19739_/D sky130_fd_sc_hd__o21a_1
X_19172_ _20428_/CLK _19172_/D vssd1 vssd1 vccd1 vccd1 _19172_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13596_/A _13596_/B vssd1 vssd1 vccd1 vccd1 _13596_/X sky130_fd_sc_hd__xor2_4
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18123_ _18126_/A _18125_/B vssd1 vssd1 vccd1 vccd1 _18123_/Y sky130_fd_sc_hd__nor2_1
XFILLER_200_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15335_ _21019_/Q _20987_/Q _15508_/S vssd1 vssd1 vccd1 vccd1 _15335_/X sky130_fd_sc_hd__mux2_1
X_12547_ _20881_/Q _12548_/B _12547_/C vssd1 vssd1 vccd1 vccd1 _12553_/C sky130_fd_sc_hd__and3_1
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18054_ _18054_/A _18054_/B _18055_/B vssd1 vssd1 vccd1 vccd1 _20757_/D sky130_fd_sc_hd__nor3_1
XFILLER_177_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15266_ _15258_/X _15264_/Y _15265_/X _15326_/A vssd1 vssd1 vccd1 vccd1 _15266_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_129_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12478_ _12582_/C vssd1 vssd1 vccd1 vccd1 _12478_/Y sky130_fd_sc_hd__inv_2
XANTENNA_3 _19658_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17005_ _19115_/Q _17005_/A2 _16945_/X _17004_/X vssd1 vssd1 vccd1 vccd1 _17005_/X
+ sky130_fd_sc_hd__o211a_1
X_14217_ _19504_/Q _14218_/B vssd1 vssd1 vccd1 vccd1 _14219_/A sky130_fd_sc_hd__nand2_1
X_11429_ _19679_/Q _20167_/Q _12133_/S vssd1 vssd1 vccd1 vccd1 _11429_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15197_ _15021_/A _14957_/B _15021_/C _15021_/X input4/X vssd1 vssd1 vccd1 vccd1
+ _15197_/X sky130_fd_sc_hd__a32o_1
XFILLER_141_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14148_ _19497_/Q _14148_/B vssd1 vssd1 vccd1 vccd1 _14160_/A sky130_fd_sc_hd__and2_1
XFILLER_259_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_258_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14079_ _14099_/A _14099_/B _14079_/C vssd1 vssd1 vccd1 vccd1 _14079_/X sky130_fd_sc_hd__or3_1
X_18956_ _19145_/Q _18976_/A2 _18767_/B vssd1 vssd1 vccd1 vccd1 _18956_/Y sky130_fd_sc_hd__a21oi_1
X_17907_ _20678_/Q _17907_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20678_/D sky130_fd_sc_hd__mux2_1
XFILLER_227_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18887_ _19135_/Q _18976_/A2 _18767_/B vssd1 vssd1 vccd1 vccd1 _18887_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1070 _12433_/A1 vssd1 vssd1 vccd1 vccd1 _12277_/A1 sky130_fd_sc_hd__buf_8
Xfanout1081 _15326_/A vssd1 vssd1 vccd1 vccd1 _15890_/B sky130_fd_sc_hd__clkbuf_8
Xfanout1092 _17706_/A1 vssd1 vssd1 vccd1 vccd1 _17915_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17838_ _20613_/Q _17910_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20613_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_282_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17769_ _20548_/Q _17909_/A1 _17774_/S vssd1 vssd1 vccd1 vccd1 _20548_/D sky130_fd_sc_hd__mux2_1
XFILLER_270_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_212_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19508_ _20930_/CLK _19508_/D vssd1 vssd1 vccd1 vccd1 _19508_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20780_ _21043_/CLK _20780_/D vssd1 vssd1 vccd1 vccd1 _20780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19439_ _20666_/CLK _19439_/D vssd1 vssd1 vccd1 vccd1 _19439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20214_ _20766_/CLK _20214_/D vssd1 vssd1 vccd1 vccd1 _20214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09956_ _20385_/Q _20449_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _09956_/X sky130_fd_sc_hd__mux2_1
X_20145_ _20716_/CLK _20145_/D vssd1 vssd1 vccd1 vccd1 _20145_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _11903_/A1 _09880_/X _09881_/X vssd1 vssd1 vccd1 vccd1 _09887_/X sky130_fd_sc_hd__o21a_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20076_ _20479_/CLK _20076_/D vssd1 vssd1 vccd1 vccd1 _20076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_264_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_253_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_404 _16919_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_415 _18220_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_426 _11260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10800_ _10798_/X _13150_/A vssd1 vssd1 vccd1 vccd1 _13541_/A sky130_fd_sc_hd__and2b_4
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_437 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _13495_/A _11780_/B vssd1 vssd1 vccd1 vccd1 _11786_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_448 _13770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_459 _19109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20978_ _21015_/CLK _20978_/D vssd1 vssd1 vccd1 vccd1 _20978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_281_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10731_ _09503_/A _10730_/X _10729_/X vssd1 vssd1 vccd1 vccd1 _10731_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_241_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_194_wb_clk_i _20408_/CLK vssd1 vssd1 vccd1 vccd1 _20698_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_198_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13450_ _13450_/A _13450_/B vssd1 vssd1 vccd1 vccd1 _13450_/Y sky130_fd_sc_hd__nor2_1
X_10662_ _12383_/A _10662_/B vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__or2_1
XFILLER_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _12401_/A1 _12400_/X _12401_/B1 vssd1 vssd1 vccd1 vccd1 _12401_/X sky130_fd_sc_hd__o21a_1
XFILLER_185_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_123_wb_clk_i clkbuf_4_13__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _19978_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13381_ _12982_/B _13376_/X _13377_/Y _13380_/X vssd1 vssd1 vccd1 vccd1 _13381_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_210_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10593_ _11680_/C1 _10589_/X _10592_/X _12072_/C1 vssd1 vssd1 vccd1 vccd1 _10593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15120_ _14883_/Y _15053_/Y _15254_/S vssd1 vssd1 vccd1 vccd1 _15121_/A sky130_fd_sc_hd__mux2_1
X_12332_ _12332_/A _19333_/Q _12406_/C vssd1 vssd1 vccd1 vccd1 _12332_/X sky130_fd_sc_hd__or3_1
XFILLER_182_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _14834_/X _14837_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _15051_/X sky130_fd_sc_hd__mux2_1
X_12263_ _12427_/A1 _19363_/Q _20718_/Q _12428_/S _12270_/B1 vssd1 vssd1 vccd1 vccd1
+ _12263_/X sky130_fd_sc_hd__a221o_1
XFILLER_182_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14002_ _14002_/A1 _09670_/Y _10462_/X _14002_/B1 _19849_/Q vssd1 vssd1 vccd1 vccd1
+ _14081_/C sky130_fd_sc_hd__o32a_1
X_11214_ _20462_/Q _12346_/S _11212_/S vssd1 vssd1 vccd1 vccd1 _11214_/X sky130_fd_sc_hd__o21a_1
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12194_ _12194_/A1 _17948_/A1 _12193_/X _12194_/B2 vssd1 vssd1 vccd1 vccd1 _15960_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18810_ _19124_/Q _18809_/X _18968_/A vssd1 vssd1 vccd1 vccd1 _18810_/X sky130_fd_sc_hd__mux2_1
X_11145_ _11235_/A _10549_/A _11144_/X vssd1 vssd1 vccd1 vccd1 _11145_/X sky130_fd_sc_hd__a21o_1
X_19790_ _20713_/CLK _19790_/D vssd1 vssd1 vccd1 vccd1 _19790_/Q sky130_fd_sc_hd__dfxtp_1
X_18741_ _20971_/Q _18285_/Y _18753_/S vssd1 vssd1 vccd1 vccd1 _18742_/B sky130_fd_sc_hd__mux2_1
XFILLER_283_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11076_ _11069_/X _11071_/X _11075_/X _12383_/A _12311_/A1 vssd1 vssd1 vccd1 vccd1
+ _11076_/X sky130_fd_sc_hd__o221a_1
X_15953_ _19554_/Q _15814_/A _15952_/Y _16187_/A vssd1 vssd1 vccd1 vccd1 _19554_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput140 dout1[3] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput151 dout1[4] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__clkbuf_2
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10027_ _19571_/Q _10026_/X _11240_/S vssd1 vssd1 vccd1 vccd1 _10027_/X sky130_fd_sc_hd__mux2_1
Xinput162 dout1[5] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_hd__clkbuf_2
X_14904_ _18198_/B _18152_/B _16133_/C _16869_/A vssd1 vssd1 vccd1 vccd1 _14904_/X
+ sky130_fd_sc_hd__a31o_4
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput173 irq[11] vssd1 vssd1 vccd1 vccd1 _12539_/C sky130_fd_sc_hd__clkbuf_2
X_18672_ _18547_/X _18684_/A2 _18670_/Y _18671_/Y vssd1 vssd1 vccd1 vccd1 _18673_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput184 irq[7] vssd1 vssd1 vccd1 vccd1 _12535_/C sky130_fd_sc_hd__clkbuf_2
X_15884_ _16051_/A1 _15870_/X _16051_/B1 vssd1 vssd1 vccd1 vccd1 _15884_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 localMemory_wb_adr_i[14] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _20379_/Q _17657_/A1 _17623_/S vssd1 vssd1 vccd1 vccd1 _20379_/D sky130_fd_sc_hd__mux2_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _14833_/X _14834_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _14835_/X sky130_fd_sc_hd__mux2_1
XFILLER_264_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17554_ _20314_/Q _17933_/A1 _17570_/S vssd1 vssd1 vccd1 vccd1 _20314_/D sky130_fd_sc_hd__mux2_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11978_ _20488_/Q _20328_/Q _11978_/S vssd1 vssd1 vccd1 vccd1 _11978_/X sky130_fd_sc_hd__mux2_1
X_14766_ _19130_/Q _14774_/A2 _14765_/X _14776_/C1 vssd1 vssd1 vccd1 vccd1 _19507_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_205_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16505_ _19812_/Q _17934_/A1 _16522_/S vssd1 vssd1 vccd1 vccd1 _19812_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10929_ _12402_/A1 _17890_/A1 _10928_/X _13675_/A vssd1 vssd1 vccd1 vccd1 _13650_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13717_ _13717_/A _13742_/B vssd1 vssd1 vccd1 vccd1 _13757_/B sky130_fd_sc_hd__or2_2
X_17485_ _17487_/A1 _17484_/Y _18126_/A vssd1 vssd1 vccd1 vccd1 _20277_/D sky130_fd_sc_hd__a21oi_1
X_14697_ _19456_/Q _17806_/A1 _14699_/S vssd1 vssd1 vccd1 vccd1 _19456_/D sky130_fd_sc_hd__mux2_1
XFILLER_205_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19224_ _19505_/CLK _19224_/D vssd1 vssd1 vccd1 vccd1 _19224_/Q sky130_fd_sc_hd__dfxtp_4
X_16436_ _19759_/Q _16437_/B vssd1 vssd1 vccd1 vccd1 _16438_/B sky130_fd_sc_hd__nor2_1
XFILLER_177_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13648_ _13653_/A _13648_/B vssd1 vssd1 vccd1 vccd1 _13718_/B sky130_fd_sc_hd__and2_4
XFILLER_176_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _21044_/CLK _19155_/D vssd1 vssd1 vccd1 vccd1 _19155_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_9_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16367_ _19733_/Q _16370_/C _18126_/A vssd1 vssd1 vccd1 vccd1 _16367_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_201_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13579_ _13577_/Y _13578_/X _20954_/Q _13564_/B vssd1 vssd1 vccd1 vccd1 _13579_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18106_ _20777_/Q _18109_/C _18104_/A vssd1 vssd1 vccd1 vccd1 _18106_/Y sky130_fd_sc_hd__a21oi_1
X_15318_ _17290_/A _15308_/B _14978_/B _14979_/Y _15317_/X vssd1 vssd1 vccd1 vccd1
+ _15318_/X sky130_fd_sc_hd__a311o_1
XFILLER_258_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16298_ _18064_/A _16298_/B vssd1 vssd1 vccd1 vccd1 _16298_/Y sky130_fd_sc_hd__nor2_1
X_19086_ _20410_/CLK _19086_/D vssd1 vssd1 vccd1 vccd1 _19086_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_172_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_274_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18037_ _18795_/A _18039_/B vssd1 vssd1 vccd1 vccd1 _18037_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15249_ _10935_/Y _15248_/X _14810_/X vssd1 vssd1 vccd1 vccd1 _15249_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_67_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09810_ _12051_/A1 _20515_/Q _12056_/S _09800_/X vssd1 vssd1 vccd1 vccd1 _09810_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_259_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19988_ _19992_/CLK _19988_/D vssd1 vssd1 vccd1 vccd1 _19988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09741_ _17709_/C _11191_/C vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__nor2_1
X_18939_ _18966_/A _18939_/B vssd1 vssd1 vccd1 vccd1 _21005_/D sky130_fd_sc_hd__nor2_1
XFILLER_268_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09672_ _09672_/A _09672_/B _09672_/C vssd1 vssd1 vccd1 vccd1 _09672_/X sky130_fd_sc_hd__or3_1
XFILLER_227_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_283_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_254_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20901_ _21011_/CLK _20901_/D vssd1 vssd1 vccd1 vccd1 _20901_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_270_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_270_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20832_ _21024_/CLK _20832_/D vssd1 vssd1 vccd1 vccd1 _20832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20763_ _20763_/CLK _20763_/D vssd1 vssd1 vccd1 vccd1 _20763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_251_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20694_ _20694_/CLK _20694_/D vssd1 vssd1 vccd1 vccd1 _20694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1806 _10284_/A vssd1 vssd1 vccd1 vccd1 _11234_/A sky130_fd_sc_hd__buf_6
Xfanout1817 _12512_/B vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__buf_8
XFILLER_81_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_278_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1828 _12513_/C vssd1 vssd1 vccd1 vccd1 _10831_/S sky130_fd_sc_hd__buf_12
Xfanout830 _13637_/A vssd1 vssd1 vccd1 vccd1 _13740_/A sky130_fd_sc_hd__buf_4
Xfanout841 _18457_/Y vssd1 vssd1 vccd1 vccd1 _18491_/B2 sky130_fd_sc_hd__buf_6
Xfanout1839 _11514_/A1 vssd1 vssd1 vccd1 vccd1 _11977_/A1 sky130_fd_sc_hd__buf_6
Xfanout852 _18311_/S vssd1 vssd1 vccd1 vccd1 _18236_/S sky130_fd_sc_hd__buf_6
X_20128_ _20703_/CLK _20128_/D vssd1 vssd1 vccd1 vccd1 _20128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_265_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09939_ _09939_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _09941_/B sky130_fd_sc_hd__nand2_2
XFILLER_265_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout863 _15323_/A vssd1 vssd1 vccd1 vccd1 _15937_/C1 sky130_fd_sc_hd__buf_6
XFILLER_120_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout874 _15942_/A2 vssd1 vssd1 vccd1 vccd1 _15999_/A2 sky130_fd_sc_hd__buf_4
Xfanout885 _15067_/S vssd1 vssd1 vccd1 vccd1 _15167_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_218_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12950_ _16716_/A _12948_/X _12949_/X _12950_/B2 vssd1 vssd1 vccd1 vccd1 _16714_/C
+ sky130_fd_sc_hd__a22o_4
Xfanout896 _16974_/A1 vssd1 vssd1 vccd1 vccd1 _16932_/A1 sky130_fd_sc_hd__buf_6
X_20059_ _20085_/CLK _20059_/D vssd1 vssd1 vccd1 vccd1 _20059_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_274_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _11892_/X _11894_/X _11900_/X _11904_/S _12137_/A1 vssd1 vssd1 vccd1 vccd1
+ _11901_/X sky130_fd_sc_hd__o221a_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _15931_/A _15527_/A _12484_/X _12880_/X vssd1 vssd1 vccd1 vccd1 _12881_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_212 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 _20005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _12143_/S _11831_/X _11830_/X _12144_/A1 vssd1 vssd1 vccd1 vccd1 _11832_/X
+ sky130_fd_sc_hd__a211o_1
X_14620_ _19384_/Q _17904_/A1 _14628_/S vssd1 vssd1 vccd1 vccd1 _19384_/D sky130_fd_sc_hd__mux2_1
XANTENNA_234 _19999_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 _20001_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_267 _20002_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ _19321_/Q _17905_/A1 _14560_/S vssd1 vssd1 vccd1 vccd1 _19321_/D sky130_fd_sc_hd__mux2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_278 _20004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11766_/B _11773_/A _13611_/A vssd1 vssd1 vccd1 vccd1 _15433_/A sky130_fd_sc_hd__a21o_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 input220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10704_/X _10713_/Y _11201_/A _10696_/X vssd1 vssd1 vccd1 vccd1 _10714_/X
+ sky130_fd_sc_hd__o2bb2a_4
X_13502_ _13501_/A _13501_/B _13501_/C vssd1 vssd1 vccd1 vccd1 _13502_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _20195_/Q _17330_/A2 _17279_/C1 _17269_/X vssd1 vssd1 vccd1 vccd1 _17270_/X
+ sky130_fd_sc_hd__a211o_1
X_14482_ _14482_/A _14482_/B vssd1 vssd1 vccd1 vccd1 _19265_/D sky130_fd_sc_hd__and2_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _19680_/Q _12097_/S _11693_/X _09834_/C vssd1 vssd1 vccd1 vccd1 _11694_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16221_ _19644_/Q _17907_/A1 _16228_/S vssd1 vssd1 vccd1 vccd1 _19644_/D sky130_fd_sc_hd__mux2_1
X_13433_ _13433_/A _13433_/B vssd1 vssd1 vccd1 vccd1 _13439_/C sky130_fd_sc_hd__xnor2_4
X_10645_ _10645_/A _11405_/A vssd1 vssd1 vccd1 vccd1 _10645_/X sky130_fd_sc_hd__or2_1
XFILLER_167_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16152_ _16815_/B _16178_/S vssd1 vssd1 vccd1 vccd1 _16152_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13364_ _13249_/Y _13362_/X _13350_/A _12664_/C vssd1 vssd1 vccd1 vccd1 _13364_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10576_ _19407_/Q _11676_/S _10575_/X _11423_/C1 vssd1 vssd1 vccd1 vccd1 _10576_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12315_ _20428_/Q _20364_/Q _12316_/S vssd1 vssd1 vccd1 vccd1 _12315_/X sky130_fd_sc_hd__mux2_1
X_15103_ _15103_/A1 _15492_/A _15102_/Y _16159_/C1 vssd1 vssd1 vccd1 vccd1 _19528_/D
+ sky130_fd_sc_hd__o211a_1
X_16083_ _19566_/Q _16079_/B _16107_/B1 vssd1 vssd1 vccd1 vccd1 _16083_/X sky130_fd_sc_hd__o21a_1
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13295_ _14275_/A1 _19228_/Q _18352_/C1 _13294_/Y vssd1 vssd1 vccd1 vccd1 _13388_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_177_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _19527_/Q _15492_/A _15031_/X _15033_/Y _16179_/A vssd1 vssd1 vccd1 vccd1
+ _19527_/D sky130_fd_sc_hd__o221a_1
XFILLER_154_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19911_ _20539_/CLK _19911_/D vssd1 vssd1 vccd1 vccd1 _19911_/Q sky130_fd_sc_hd__dfxtp_1
X_12246_ _12403_/A1 _12245_/Y _12403_/B1 vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__o21a_2
Xclkbuf_leaf_91_wb_clk_i clkbuf_leaf_99_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _19589_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19842_ _20014_/CLK _19842_/D vssd1 vssd1 vccd1 vccd1 _19842_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_69_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_269_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12177_ _11851_/A _20050_/Q _12011_/S _12160_/X vssd1 vssd1 vccd1 vccd1 _12177_/X
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_20_wb_clk_i _20408_/CLK vssd1 vssd1 vccd1 vccd1 _20438_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11128_ _12347_/A1 _20120_/Q _20088_/Q _11126_/B vssd1 vssd1 vccd1 vccd1 _11128_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_268_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19773_ _20468_/CLK _19773_/D vssd1 vssd1 vccd1 vccd1 _19773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16985_ _16982_/Y _16984_/Y _16985_/B1 vssd1 vssd1 vccd1 vccd1 _16985_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_283_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18724_ _18724_/A _18724_/B vssd1 vssd1 vccd1 vccd1 _20962_/D sky130_fd_sc_hd__and2_1
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ input129/X input134/X _11241_/S vssd1 vssd1 vccd1 vccd1 _11059_/X sky130_fd_sc_hd__mux2_8
X_15936_ _21039_/Q _21007_/Q _15993_/S vssd1 vssd1 vccd1 vccd1 _15936_/X sky130_fd_sc_hd__mux2_1
XFILLER_260_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18655_ _19517_/Q _18683_/B vssd1 vssd1 vccd1 vccd1 _18655_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _15843_/A _15866_/X _15895_/S vssd1 vssd1 vccd1 vccd1 _15867_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17606_ _20364_/Q _17917_/A1 _17606_/S vssd1 vssd1 vccd1 vccd1 _20364_/D sky130_fd_sc_hd__mux2_1
XFILLER_252_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14818_ _09861_/B _10636_/Y _14822_/S vssd1 vssd1 vccd1 vccd1 _14818_/X sky130_fd_sc_hd__mux2_1
X_18586_ _18480_/X _18621_/A2 _18584_/Y _18585_/Y vssd1 vssd1 vccd1 vccd1 _18587_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ _20744_/Q _15934_/A2 _15934_/B1 _20776_/Q vssd1 vssd1 vccd1 vccd1 _15798_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_251_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_251_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ _17537_/A _17537_/B _17537_/C vssd1 vssd1 vccd1 vccd1 _20300_/D sky130_fd_sc_hd__and3_1
XFILLER_83_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14749_ _19499_/Q _14763_/B vssd1 vssd1 vccd1 vccd1 _14749_/X sky130_fd_sc_hd__or2_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_225_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17468_ _20269_/Q _17494_/B vssd1 vssd1 vccd1 vccd1 _17468_/Y sky130_fd_sc_hd__nand2_1
X_19207_ _20665_/CLK _19207_/D vssd1 vssd1 vccd1 vccd1 _19207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16419_ _18821_/A _16419_/B _16420_/B vssd1 vssd1 vccd1 vccd1 _19752_/D sky130_fd_sc_hd__nor3_1
X_17399_ _20248_/Q _17401_/A2 _17398_/X _17536_/D vssd1 vssd1 vccd1 vccd1 _20248_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_285_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19138_ _20291_/CLK _19138_/D vssd1 vssd1 vccd1 vccd1 _19138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19069_ _20414_/Q vssd1 vssd1 vccd1 vccd1 _20414_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput400 _13822_/X vssd1 vssd1 vccd1 vccd1 din0[31] sky130_fd_sc_hd__buf_4
Xoutput411 _19971_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[10] sky130_fd_sc_hd__buf_4
Xoutput422 _19981_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[20] sky130_fd_sc_hd__buf_4
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput433 _19991_/Q vssd1 vssd1 vccd1 vccd1 localMemory_wb_data_o[30] sky130_fd_sc_hd__buf_4
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput444 _13192_/Y vssd1 vssd1 vccd1 vccd1 probe_env[1] sky130_fd_sc_hd__buf_4
Xoutput455 _19508_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[14] sky130_fd_sc_hd__buf_4
XFILLER_271_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput466 _19518_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[24] sky130_fd_sc_hd__buf_4
XFILLER_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21031_ _21043_/CLK _21031_/D vssd1 vssd1 vccd1 vccd1 _21031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput477 _19499_/Q vssd1 vssd1 vccd1 vccd1 probe_programCounter[5] sky130_fd_sc_hd__buf_4
XFILLER_248_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09724_ _09709_/X _09723_/X _12153_/A1 vssd1 vssd1 vccd1 vccd1 _09724_/X sky130_fd_sc_hd__a21o_1
XFILLER_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_255_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09655_ _19695_/Q _19655_/Q vssd1 vssd1 vccd1 vccd1 _09655_/Y sky130_fd_sc_hd__nand2_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_283_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_271_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_283_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_243_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_271_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_215_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09586_ _09596_/A vssd1 vssd1 vccd1 vccd1 _09586_/Y sky130_fd_sc_hd__inv_2
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_250_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_270_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20815_ _20990_/CLK _20815_/D vssd1 vssd1 vccd1 vccd1 _20815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_270_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20746_ _20812_/CLK _20746_/D vssd1 vssd1 vccd1 vccd1 _20746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_259_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20677_ _20677_/CLK _20677_/D vssd1 vssd1 vccd1 vccd1 _20677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10430_ _10428_/X _10429_/X _10430_/S vssd1 vssd1 vccd1 vccd1 _10430_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10361_ _10340_/X _10348_/X _10354_/X _10360_/X vssd1 vssd1 vccd1 vccd1 _10361_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12100_ _20487_/Q _12097_/S _12100_/B1 vssd1 vssd1 vccd1 vccd1 _12100_/X sky130_fd_sc_hd__o21a_1
XFILLER_275_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ _13025_/Y _13368_/A _13367_/B vssd1 vssd1 vccd1 vccd1 _13270_/C sky130_fd_sc_hd__o21ai_4
X_10292_ _10035_/Y _10286_/X _10291_/X _10284_/X _10024_/X vssd1 vssd1 vccd1 vccd1
+ _10293_/B sky130_fd_sc_hd__a32o_2
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12031_ _15931_/A vssd1 vssd1 vccd1 vccd1 _12031_/Y sky130_fd_sc_hd__inv_2
XFILLER_278_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1603 _12063_/C1 vssd1 vssd1 vccd1 vccd1 _11995_/S sky130_fd_sc_hd__buf_8
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1614 _11988_/S vssd1 vssd1 vccd1 vccd1 _12134_/S sky130_fd_sc_hd__buf_6
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1625 _12376_/S vssd1 vssd1 vccd1 vccd1 _12395_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1636 _09614_/X vssd1 vssd1 vccd1 vccd1 _12073_/C1 sky130_fd_sc_hd__buf_4
Xfanout1647 _18955_/A vssd1 vssd1 vccd1 vccd1 _18975_/A sky130_fd_sc_hd__buf_6
XFILLER_265_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1658 _11239_/B1 vssd1 vssd1 vccd1 vccd1 _11228_/B1 sky130_fd_sc_hd__buf_8
Xfanout660 _14773_/B vssd1 vssd1 vccd1 vccd1 _14763_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout671 _13921_/B vssd1 vssd1 vccd1 vccd1 _13919_/S sky130_fd_sc_hd__buf_4
XFILLER_59_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1669 _14029_/A1 vssd1 vssd1 vccd1 vccd1 _14035_/A1 sky130_fd_sc_hd__buf_4
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_247_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout682 _13863_/B vssd1 vssd1 vccd1 vccd1 _13953_/A2 sky130_fd_sc_hd__buf_4
X_16770_ _16770_/A vssd1 vssd1 vccd1 vccd1 _16770_/Y sky130_fd_sc_hd__clkinv_4
X_13982_ _19193_/Q _14067_/C _14042_/S vssd1 vssd1 vccd1 vccd1 _13982_/X sky130_fd_sc_hd__mux2_1
Xfanout693 _13790_/X vssd1 vssd1 vccd1 vccd1 split9/A sky130_fd_sc_hd__buf_6
XFILLER_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_281_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15721_ _20965_/Q _15939_/A2 _15996_/B1 _20837_/Q _15720_/X vssd1 vssd1 vccd1 vccd1
+ _15721_/X sky130_fd_sc_hd__a221o_1
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12933_ _19261_/Q _12950_/B2 _16716_/A _20009_/Q vssd1 vssd1 vccd1 vccd1 _16720_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18440_ _18740_/A _18440_/B vssd1 vssd1 vccd1 vccd1 _20874_/D sky130_fd_sc_hd__and2_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15652_ _15652_/A _15652_/B _15981_/B vssd1 vssd1 vccd1 vccd1 _15652_/X sky130_fd_sc_hd__and3_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ _13300_/B _12864_/B vssd1 vssd1 vccd1 vccd1 _12864_/Y sky130_fd_sc_hd__nand2b_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _19367_/Q _17887_/A1 _14633_/S vssd1 vssd1 vccd1 vccd1 _19367_/D sky130_fd_sc_hd__mux2_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _18535_/B _18375_/B vssd1 vssd1 vccd1 vccd1 _18371_/Y sky130_fd_sc_hd__nand2_1
X_11815_ _20485_/Q _20325_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _11815_/X sky130_fd_sc_hd__mux2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _13426_/B _15982_/C _16056_/B1 vssd1 vssd1 vccd1 vccd1 _15583_/Y sky130_fd_sc_hd__a21oi_1
X_12795_ _13586_/A _12790_/D _12790_/C vssd1 vssd1 vccd1 vccd1 _12795_/X sky130_fd_sc_hd__o21ba_1
XFILLER_215_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _20213_/Q _17328_/A2 _17321_/X _18416_/A vssd1 vssd1 vccd1 vccd1 _20213_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ _19304_/Q _17679_/A1 _14563_/S vssd1 vssd1 vccd1 vccd1 _19304_/D sky130_fd_sc_hd__mux2_1
XFILLER_144_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11746_ _10018_/Y _11745_/X _13414_/A vssd1 vssd1 vccd1 vccd1 _15789_/A sky130_fd_sc_hd__a21o_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ _20190_/Q _17268_/A2 _17251_/X _17252_/X _17274_/C1 vssd1 vssd1 vccd1 vccd1
+ _20190_/D sky130_fd_sc_hd__o221a_1
X_14465_ _20228_/Q _19257_/Q _14469_/S vssd1 vssd1 vccd1 vccd1 _14466_/B sky130_fd_sc_hd__mux2_1
XFILLER_174_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11677_ _09806_/S _11676_/X _11675_/X _11680_/C1 vssd1 vssd1 vccd1 vccd1 _11677_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16204_ _19627_/Q _17890_/A1 _16231_/S vssd1 vssd1 vccd1 vccd1 _19627_/D sky130_fd_sc_hd__mux2_1
X_13416_ _13416_/A _13416_/B vssd1 vssd1 vccd1 vccd1 _13417_/A sky130_fd_sc_hd__xnor2_4
X_10628_ _19874_/Q _19775_/Q _10628_/S vssd1 vssd1 vccd1 vccd1 _10629_/B sky130_fd_sc_hd__mux2_1
XFILLER_128_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17184_ _17184_/A _17812_/A vssd1 vssd1 vccd1 vccd1 _17185_/C sky130_fd_sc_hd__nor2_1
X_14396_ _13139_/A _14395_/X _13218_/Y vssd1 vssd1 vccd1 vccd1 _14397_/C sky130_fd_sc_hd__a21bo_1
X_16135_ _19591_/Q _16196_/S _16134_/Y _16165_/C1 vssd1 vssd1 vccd1 vccd1 _19591_/D
+ sky130_fd_sc_hd__o211a_1
X_13347_ _13347_/A _13347_/B vssd1 vssd1 vccd1 vccd1 _13347_/Y sky130_fd_sc_hd__nand2_1
X_10559_ _10037_/Y _10558_/Y _09669_/X vssd1 vssd1 vccd1 vccd1 _10559_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13278_ _12701_/A _12701_/B _12791_/C _12791_/D vssd1 vssd1 vccd1 vccd1 _13279_/B
+ sky130_fd_sc_hd__a211oi_1
X_16066_ _16066_/A _16066_/B vssd1 vssd1 vccd1 vccd1 _16068_/C sky130_fd_sc_hd__nor2_2
XFILLER_64_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12229_ _12310_/C1 _12228_/X _12225_/X _12385_/C1 vssd1 vssd1 vccd1 vccd1 _12229_/X
+ sky130_fd_sc_hd__a211o_2
X_15017_ _15020_/A _15022_/D _15508_/S vssd1 vssd1 vccd1 vccd1 _15017_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_269_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_284_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19825_ _19956_/CLK _19825_/D vssd1 vssd1 vccd1 vccd1 _19825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_271_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_269_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19756_ _20962_/CLK _19756_/D vssd1 vssd1 vccd1 vccd1 _19756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16968_ _16950_/Y _16967_/X _16875_/B2 vssd1 vssd1 vccd1 vccd1 _16968_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_256_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_284_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_237_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18707_ _20954_/Q _18200_/Y _18707_/S vssd1 vssd1 vccd1 vccd1 _18708_/B sky130_fd_sc_hd__mux2_1
XFILLER_253_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15919_ _16024_/A1 _15917_/X _15918_/X _15898_/A _15975_/B2 vssd1 vssd1 vccd1 vccd1
+ _15919_/X sky130_fd_sc_hd__a32o_1
X_19687_ _20481_/CLK _19687_/D vssd1 vssd1 vccd1 vccd1 _19687_/Q sky130_fd_sc_hd__dfxtp_1
X_16899_ _16981_/A1 _15698_/X _16879_/X _16898_/X vssd1 vssd1 vccd1 vccd1 _16899_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_225_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18638_ _18891_/A _18638_/B vssd1 vssd1 vccd1 vccd1 _20932_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18569_ _20915_/Q _18619_/B vssd1 vssd1 vccd1 vccd1 _18569_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20600_ _20683_/CLK _20600_/D vssd1 vssd1 vccd1 vccd1 _20600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20531_ _20663_/CLK _20531_/D vssd1 vssd1 vccd1 vccd1 _20531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20462_ _20694_/CLK _20462_/D vssd1 vssd1 vccd1 vccd1 _20462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20393_ _20645_/CLK _20393_/D vssd1 vssd1 vccd1 vccd1 _20393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_279_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput285 _13827_/X vssd1 vssd1 vccd1 vccd1 addr0[0] sky130_fd_sc_hd__buf_4
XFILLER_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21014_ _21016_/CLK _21014_/D vssd1 vssd1 vccd1 vccd1 _21014_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput296 _13783_/X vssd1 vssd1 vccd1 vccd1 addr1[2] sky130_fd_sc_hd__buf_4
XFILLER_0_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_275_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_263_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09707_ _11903_/A1 _09700_/X _09701_/X vssd1 vssd1 vccd1 vccd1 _09707_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09638_ _18163_/B _11235_/A vssd1 vssd1 vccd1 vccd1 _09638_/Y sky130_fd_sc_hd__nand2_8
XFILLER_16_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_231_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09569_ _09569_/A _15442_/A vssd1 vssd1 vccd1 vccd1 _13657_/A sky130_fd_sc_hd__nor2_8
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11600_ _11980_/S _11599_/X _11598_/X _11600_/C1 vssd1 vssd1 vccd1 vccd1 _11600_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12580_ _12580_/A _12580_/B vssd1 vssd1 vccd1 vccd1 _12581_/B sky130_fd_sc_hd__nor2_4
XFILLER_230_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11531_ _11516_/X _11530_/X _12153_/A1 vssd1 vssd1 vccd1 vccd1 _11531_/X sky130_fd_sc_hd__a21o_2
X_20729_ _20763_/CLK _20729_/D vssd1 vssd1 vccd1 vccd1 _20729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_278_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14250_ _14250_/A _14250_/B _14250_/C vssd1 vssd1 vccd1 vccd1 _14252_/B sky130_fd_sc_hd__and3_1
XFILLER_139_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11462_ _19479_/Q _19447_/Q _12185_/S vssd1 vssd1 vccd1 vccd1 _11462_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _19238_/Q _19237_/Q _13390_/B _19239_/Q vssd1 vssd1 vccd1 vccd1 _13201_/Y
+ sky130_fd_sc_hd__a31oi_1
X_10413_ _19634_/Q _19940_/Q _19278_/Q _20065_/Q _10092_/S _12084_/C vssd1 vssd1 vccd1
+ vccd1 _10413_/X sky130_fd_sc_hd__mux4_1
XFILLER_171_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14181_ _14181_/A _14181_/B vssd1 vssd1 vccd1 vccd1 _14182_/B sky130_fd_sc_hd__xnor2_1
XFILLER_99_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11393_ _20405_/Q _20341_/Q _20633_/Q _20597_/Q _11393_/S0 _11391_/C vssd1 vssd1
+ vccd1 vccd1 _11393_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ _20943_/Q _13366_/C1 _18687_/B vssd1 vssd1 vccd1 vccd1 _13132_/Y sky130_fd_sc_hd__a21oi_1
X_10344_ _19676_/Q _20164_/Q _11295_/S vssd1 vssd1 vccd1 vccd1 _10344_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13063_ _20951_/Q _20885_/Q _13062_/Y vssd1 vssd1 vccd1 vccd1 _13064_/D sky130_fd_sc_hd__a21o_1
X_17940_ _20709_/Q _17940_/A1 _17948_/S vssd1 vssd1 vccd1 vccd1 _20709_/D sky130_fd_sc_hd__mux2_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10275_ _10277_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _15613_/S sky130_fd_sc_hd__nand2_4
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_285_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1400 _10092_/S vssd1 vssd1 vccd1 vccd1 _10400_/S sky130_fd_sc_hd__buf_6
X_12014_ _09752_/A _19489_/Q _19457_/Q _12013_/S _12016_/C1 vssd1 vssd1 vccd1 vccd1
+ _12014_/X sky130_fd_sc_hd__a221o_1
XFILLER_79_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_278_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1411 _10174_/S vssd1 vssd1 vccd1 vccd1 _11039_/S sky130_fd_sc_hd__buf_2
Xfanout1422 fanout1430/X vssd1 vssd1 vccd1 vccd1 fanout1422/X sky130_fd_sc_hd__clkbuf_8
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17871_ _20644_/Q _17871_/A1 _17880_/S vssd1 vssd1 vccd1 vccd1 _20644_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout1433 _11852_/B2 vssd1 vssd1 vccd1 vccd1 _12190_/C1 sky130_fd_sc_hd__buf_6
X_19610_ _19617_/CLK _19610_/D vssd1 vssd1 vccd1 vccd1 _19610_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout1444 _10611_/B vssd1 vssd1 vccd1 vccd1 _09986_/C sky130_fd_sc_hd__buf_8
XFILLER_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1455 _12411_/C vssd1 vssd1 vccd1 vccd1 _12406_/C sky130_fd_sc_hd__clkbuf_8
X_16822_ _16822_/A _16822_/B vssd1 vssd1 vccd1 vccd1 _16822_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1466 _11204_/S vssd1 vssd1 vccd1 vccd1 _11933_/S sky130_fd_sc_hd__buf_4
Xfanout1477 _09731_/Y vssd1 vssd1 vccd1 vccd1 _11204_/S sky130_fd_sc_hd__buf_12
XFILLER_94_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout490 _17934_/S vssd1 vssd1 vccd1 vccd1 _17951_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_266_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1488 _09729_/Y vssd1 vssd1 vccd1 vccd1 _11396_/S sky130_fd_sc_hd__buf_12
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1499 _12041_/B vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__buf_6
XFILLER_65_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19541_ _19541_/CLK _19541_/D vssd1 vssd1 vccd1 vccd1 _19541_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_235_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16753_ _19963_/Q _16822_/A _16752_/Y _18801_/A vssd1 vssd1 vccd1 vccd1 _19963_/D
+ sky130_fd_sc_hd__a211o_1
X_13965_ _19155_/Q _19050_/S _14043_/B1 _13964_/X _16097_/B1 vssd1 vssd1 vccd1 vccd1
+ _19155_/D sky130_fd_sc_hd__o221a_1
XFILLER_111_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15704_ _19168_/Q _15978_/A2 _13427_/A _15922_/B2 vssd1 vssd1 vccd1 vccd1 _15705_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19472_ _21047_/A _19472_/D vssd1 vssd1 vccd1 vccd1 _19472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12916_ _14433_/A _12916_/A2 _12915_/X _12916_/B2 vssd1 vssd1 vccd1 vccd1 _12917_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_80_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16684_ _19939_/Q _17896_/A1 _16705_/S vssd1 vssd1 vccd1 vccd1 _19939_/D sky130_fd_sc_hd__mux2_1
XFILLER_250_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13896_ _19114_/Q _14527_/A2 _13896_/B1 _12512_/B _16195_/A vssd1 vssd1 vccd1 vccd1
+ _19114_/D sky130_fd_sc_hd__o221a_1
XFILLER_62_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18423_ _20866_/Q _18240_/Y _18449_/S vssd1 vssd1 vccd1 vccd1 _18424_/B sky130_fd_sc_hd__mux2_1
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ _21028_/Q _20996_/Q _15993_/S vssd1 vssd1 vccd1 vccd1 _15635_/X sky130_fd_sc_hd__mux2_1
X_12847_ split8/X _12847_/A2 _15526_/A _12846_/Y vssd1 vssd1 vccd1 vccd1 _12847_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_250_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18354_ _20832_/Q _18363_/B _18353_/Y _18720_/A vssd1 vssd1 vccd1 vccd1 _20832_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_199_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _20896_/Q _15937_/A2 _15566_/B1 _15565_/X _15937_/C1 vssd1 vssd1 vccd1 vccd1
+ _15566_/X sky130_fd_sc_hd__a221o_1
XFILLER_221_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12776_/Y _12777_/X _11367_/A _13589_/A1 vssd1 vssd1 vccd1 vccd1 _13586_/A
+ sky130_fd_sc_hd__o211a_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17305_/A _17329_/S _17305_/C vssd1 vssd1 vccd1 vccd1 _17305_/X sky130_fd_sc_hd__and3_1
XFILLER_30_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14517_ _19295_/Q _17112_/A1 _14517_/S vssd1 vssd1 vccd1 vccd1 _19295_/D sky130_fd_sc_hd__mux2_1
XFILLER_187_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18285_ _18541_/B vssd1 vssd1 vccd1 vccd1 _18285_/Y sky130_fd_sc_hd__clkinv_2
X_11729_ _11729_/A _11733_/B vssd1 vssd1 vccd1 vccd1 _11730_/B sky130_fd_sc_hd__and2_4
XFILLER_175_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15497_ _14841_/S _15211_/X _15496_/X vssd1 vssd1 vccd1 vccd1 _15497_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17236_ _17236_/A _17337_/B vssd1 vssd1 vccd1 vccd1 _17236_/Y sky130_fd_sc_hd__nand2_1
X_14448_ _18702_/A _14448_/B vssd1 vssd1 vccd1 vccd1 _19248_/D sky130_fd_sc_hd__and2_1
XFILLER_163_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17167_ _20133_/Q _17692_/A1 _17183_/S vssd1 vssd1 vccd1 vccd1 _20133_/D sky130_fd_sc_hd__mux2_1
XFILLER_143_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14379_ _14437_/A _14437_/B _14379_/C vssd1 vssd1 vccd1 vccd1 _14379_/X sky130_fd_sc_hd__or3_1
XFILLER_155_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16118_ _11228_/X _16132_/A2 _16117_/X vssd1 vssd1 vccd1 vccd1 _19583_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17098_ _20068_/Q _17934_/A1 _17115_/S vssd1 vssd1 vccd1 vccd1 _20068_/D sky130_fd_sc_hd__mux2_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_282_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16049_ _16049_/A1 _16038_/X _16039_/X _16048_/X vssd1 vssd1 vccd1 vccd1 _16049_/X
+ sky130_fd_sc_hd__a22o_4
XFILLER_170_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_276_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_229_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19808_ _20539_/CLK _19808_/D vssd1 vssd1 vccd1 vccd1 _19808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_285_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19739_ _20759_/CLK _19739_/D vssd1 vssd1 vccd1 vccd1 _19739_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_272_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20514_ _20646_/CLK _20514_/D vssd1 vssd1 vccd1 vccd1 _20514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20445_ _20573_/CLK _20445_/D vssd1 vssd1 vccd1 vccd1 _20445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_256_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20376_ _20568_/CLK _20376_/D vssd1 vssd1 vccd1 vccd1 _20376_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_279_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_279_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_148_wb_clk_i clkbuf_4_7__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _21025_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _20637_/Q _12044_/B _11684_/A1 vssd1 vssd1 vccd1 vccd1 _10060_/X sky130_fd_sc_hd__a21o_1
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_263_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10962_ _11309_/A1 _10957_/X _10961_/X _11384_/S vssd1 vssd1 vccd1 vccd1 _10963_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13750_ _13765_/A _13750_/B vssd1 vssd1 vccd1 vccd1 _13750_/X sky130_fd_sc_hd__and2_2
XFILLER_44_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12701_ _12701_/A _12701_/B vssd1 vssd1 vccd1 vccd1 _13571_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10893_ _19563_/Q _09666_/B _09659_/X _10892_/Y vssd1 vssd1 vccd1 vccd1 _10893_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13681_ _13718_/A _13718_/B vssd1 vssd1 vccd1 vccd1 _13681_/Y sky130_fd_sc_hd__nor2_2
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15420_ _20859_/Q _15419_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15420_/X sky130_fd_sc_hd__mux2_1
XPHY_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12632_ _15331_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _12632_/Y sky130_fd_sc_hd__nand2_1
XPHY_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15351_ _11788_/A _15494_/B _15350_/Y vssd1 vssd1 vccd1 vccd1 _15351_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12563_ _13658_/A _13740_/B vssd1 vssd1 vccd1 vccd1 _12563_/Y sky130_fd_sc_hd__nor2_1
XFILLER_197_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11514_ _11514_/A1 _11507_/X _11508_/X vssd1 vssd1 vccd1 vccd1 _11514_/X sky130_fd_sc_hd__o21a_1
X_14302_ _14302_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14303_/B sky130_fd_sc_hd__nor2_1
X_18070_ _18080_/A _18070_/B _18071_/B vssd1 vssd1 vccd1 vccd1 _20763_/D sky130_fd_sc_hd__nor3_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12494_ _11219_/X _12738_/B _12493_/X vssd1 vssd1 vccd1 vccd1 _12496_/B sky130_fd_sc_hd__o21ai_4
X_15282_ _15282_/A _16774_/B vssd1 vssd1 vccd1 vccd1 _15282_/X sky130_fd_sc_hd__or2_1
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17021_ _19999_/Q input208/X _17849_/S vssd1 vssd1 vccd1 vccd1 _19999_/D sky130_fd_sc_hd__mux2_1
XFILLER_172_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11445_ _12143_/S _11444_/X _11443_/X _12144_/A1 vssd1 vssd1 vccd1 vccd1 _11445_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14233_ _14229_/B _14232_/X _14233_/S vssd1 vssd1 vccd1 vccd1 _14233_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ _18763_/A1 _14163_/X _13520_/X vssd1 vssd1 vccd1 vccd1 _14165_/C sky130_fd_sc_hd__a21o_1
XFILLER_171_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11376_ _12427_/A1 _19470_/Q _19438_/Q _11377_/S vssd1 vssd1 vccd1 vccd1 _11376_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10327_ _09689_/A _10319_/X _10326_/X _10310_/X vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_4_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13115_ _12998_/Y _13114_/X _13002_/A vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__a21o_1
X_14095_ _14107_/A _14099_/B _14095_/C vssd1 vssd1 vccd1 vccd1 _14095_/X sky130_fd_sc_hd__or3_1
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18972_ _18556_/X _18971_/B _18970_/X _18971_/Y vssd1 vssd1 vccd1 vccd1 _18973_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_180_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17923_ _20692_/Q _17923_/A1 _17951_/S vssd1 vssd1 vccd1 vccd1 _20692_/D sky130_fd_sc_hd__mux2_1
X_13046_ _20955_/Q _20889_/Q vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__and2_1
X_10258_ _10255_/X _10256_/X _10257_/X _12429_/A1 _12430_/S vssd1 vssd1 vccd1 vccd1
+ _10258_/X sky130_fd_sc_hd__a221o_1
XFILLER_285_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1230 _12493_/A vssd1 vssd1 vccd1 vccd1 _12731_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1241 _13661_/A vssd1 vssd1 vccd1 vccd1 _13653_/A sky130_fd_sc_hd__buf_12
X_17854_ _20627_/Q _17888_/A1 _17882_/S vssd1 vssd1 vccd1 vccd1 _20627_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10189_ _19379_/Q _11192_/A2 _10187_/X _15129_/A0 _10188_/X vssd1 vssd1 vccd1 vccd1
+ _10189_/X sky130_fd_sc_hd__o221a_1
XFILLER_182_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1252 _17371_/A2 vssd1 vssd1 vccd1 vccd1 _17363_/A2 sky130_fd_sc_hd__buf_6
XFILLER_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1263 _12075_/C1 vssd1 vssd1 vccd1 vccd1 _12153_/B1 sky130_fd_sc_hd__clkbuf_16
XFILLER_227_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1274 _15303_/A vssd1 vssd1 vccd1 vccd1 _15442_/A sky130_fd_sc_hd__buf_6
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16805_ _20622_/Q _16945_/B _16945_/C vssd1 vssd1 vccd1 vccd1 _16805_/X sky130_fd_sc_hd__and3_4
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1285 _15922_/B2 vssd1 vssd1 vccd1 vccd1 _16063_/B2 sky130_fd_sc_hd__buf_6
XFILLER_208_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1296 _12708_/B vssd1 vssd1 vccd1 vccd1 _12752_/B sky130_fd_sc_hd__buf_6
XFILLER_82_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17785_ _20562_/Q _17925_/A1 _17811_/S vssd1 vssd1 vccd1 vccd1 _20562_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14997_ _15019_/B _15019_/C _14997_/C vssd1 vssd1 vccd1 vccd1 _14997_/X sky130_fd_sc_hd__and3_1
XFILLER_226_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_254_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19524_ _20296_/CLK _19524_/D vssd1 vssd1 vccd1 vccd1 _19524_/Q sky130_fd_sc_hd__dfxtp_4
X_16736_ _17219_/B _16732_/Y _16734_/X _12952_/X vssd1 vssd1 vccd1 vccd1 _16736_/X
+ sky130_fd_sc_hd__a31o_1
X_13948_ _14002_/A1 _13960_/A2 _11238_/X _14002_/B1 _19831_/Q vssd1 vssd1 vccd1 vccd1
+ _14045_/C sky130_fd_sc_hd__o32a_1
XFILLER_47_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_208_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_262_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19455_ _20708_/CLK _19455_/D vssd1 vssd1 vccd1 vccd1 _19455_/Q sky130_fd_sc_hd__dfxtp_1
X_16667_ _19924_/Q _17111_/A1 _16668_/S vssd1 vssd1 vccd1 vccd1 _19924_/D sky130_fd_sc_hd__mux2_1
X_13879_ _12967_/B _14527_/A2 _13900_/A2 _19163_/Q _16195_/A vssd1 vssd1 vccd1 vccd1
+ _19097_/D sky130_fd_sc_hd__o221a_1
XFILLER_201_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_250_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18406_ _18418_/A _18406_/B vssd1 vssd1 vccd1 vccd1 _20857_/D sky130_fd_sc_hd__and2_1
XFILLER_250_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15618_ _11757_/Y _16028_/C _15617_/X _15890_/B vssd1 vssd1 vccd1 vccd1 _15618_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_195_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19386_ _20585_/CLK _19386_/D vssd1 vssd1 vccd1 vccd1 _19386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16598_ _16598_/A _16598_/B _16598_/C vssd1 vssd1 vccd1 vccd1 _16598_/X sky130_fd_sc_hd__or3_2
XFILLER_50_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_277_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18337_ _18483_/B _18343_/B vssd1 vssd1 vccd1 vccd1 _18337_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15549_ _15984_/A2 _15264_/B _15549_/S vssd1 vssd1 vccd1 vccd1 _15549_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18268_ _19549_/Q _18308_/B vssd1 vssd1 vccd1 vccd1 _18268_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_148_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _17219_/A _17219_/B _17219_/C vssd1 vssd1 vccd1 vccd1 _17219_/Y sky130_fd_sc_hd__nand3_2
X_18199_ _18199_/A1 _14198_/B _18198_/Y vssd1 vssd1 vccd1 vccd1 _18490_/B sky130_fd_sc_hd__o21ai_4
XFILLER_144_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20230_ _21016_/CLK _20230_/D vssd1 vssd1 vccd1 vccd1 _20230_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20161_ _20711_/CLK _20161_/D vssd1 vssd1 vccd1 vccd1 _20161_/Q sky130_fd_sc_hd__dfxtp_1
X_09972_ _12134_/S _09971_/X _09970_/X _12147_/C1 vssd1 vssd1 vccd1 vccd1 _09972_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_277_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20092_ _20563_/CLK _20092_/D vssd1 vssd1 vccd1 vccd1 _20092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_276_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_269_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_285_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_258_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_285_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_268_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_608 input217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_619 _20000_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20994_ _21024_/CLK _20994_/D vssd1 vssd1 vccd1 vccd1 _20994_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_272_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_240_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_275_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_267_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _11230_/A _11236_/C vssd1 vssd1 vccd1 vccd1 _11230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20428_ _20428_/CLK _20428_/D vssd1 vssd1 vccd1 vccd1 _20428_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _20398_/Q _20334_/Q _11161_/S vssd1 vssd1 vccd1 vccd1 _11161_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20359_ _20683_/CLK _20359_/D vssd1 vssd1 vccd1 vccd1 _20359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_283_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10112_ _10112_/A _11412_/B vssd1 vssd1 vccd1 vccd1 _15500_/S sky130_fd_sc_hd__nand2_2
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11092_ _20024_/Q _19899_/Q _11093_/S vssd1 vssd1 vccd1 vccd1 _11092_/X sky130_fd_sc_hd__mux2_1
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xsplit7 split7/A vssd1 vssd1 vccd1 vccd1 split7/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14920_ _14920_/A _15022_/A _14951_/C vssd1 vssd1 vccd1 vccd1 _14980_/B sky130_fd_sc_hd__or3_2
X_10043_ _10034_/X _10035_/Y _10042_/X _10028_/X _10024_/X vssd1 vssd1 vccd1 vccd1
+ _10044_/B sky130_fd_sc_hd__a32o_2
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_275_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14851_ _14849_/X _14850_/X _15058_/S vssd1 vssd1 vccd1 vccd1 _14851_/X sky130_fd_sc_hd__mux2_1
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13802_ _13802_/A1 _13683_/B _13805_/B1 input217/X vssd1 vssd1 vccd1 vccd1 _13802_/X
+ sky130_fd_sc_hd__a22o_1
X_17570_ _20330_/Q _17706_/A1 _17570_/S vssd1 vssd1 vccd1 vccd1 _20330_/D sky130_fd_sc_hd__mux2_1
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14782_ _19138_/Q _14802_/A2 _14781_/X _17393_/C1 vssd1 vssd1 vccd1 vccd1 _19515_/D
+ sky130_fd_sc_hd__o211a_1
X_11994_ _19294_/Q _20081_/Q _11994_/S vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__mux2_1
XFILLER_216_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16521_ _19828_/Q _17114_/A1 _16521_/S vssd1 vssd1 vccd1 vccd1 _19828_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13733_ _13780_/A _13733_/B vssd1 vssd1 vccd1 vccd1 _13733_/X sky130_fd_sc_hd__and2_1
X_10945_ _10943_/X _10944_/X _11033_/S vssd1 vssd1 vccd1 vccd1 _10945_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_wb_clk_i clkbuf_4_8__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20565_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_204_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19240_ _19520_/CLK _19240_/D vssd1 vssd1 vccd1 vccd1 _19240_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16452_ _19765_/Q _16451_/C _16451_/A vssd1 vssd1 vccd1 vccd1 _16452_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_189_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13664_ _13664_/A _13684_/B vssd1 vssd1 vccd1 vccd1 _13665_/A sky130_fd_sc_hd__and2_4
XFILLER_232_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10876_ _19403_/Q _20562_/Q _12344_/S vssd1 vssd1 vccd1 vccd1 _10876_/X sky130_fd_sc_hd__mux2_1
X_15403_ _19535_/Q _15402_/A _15402_/Y _16143_/A vssd1 vssd1 vccd1 vccd1 _19535_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19171_ _20426_/CLK _19171_/D vssd1 vssd1 vccd1 vccd1 _19171_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _19524_/Q _12624_/A vssd1 vssd1 vccd1 vccd1 _12914_/B sky130_fd_sc_hd__nand2_2
X_16383_ _19739_/Q _16386_/C _18056_/A vssd1 vssd1 vccd1 vccd1 _16383_/Y sky130_fd_sc_hd__a21oi_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _13595_/A _13921_/A vssd1 vssd1 vccd1 vccd1 _13595_/Y sky130_fd_sc_hd__nor2_2
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18122_ _20783_/Q _20782_/Q _18122_/C vssd1 vssd1 vccd1 vccd1 _18125_/B sky130_fd_sc_hd__and3_1
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15334_ input8/X _15334_/B vssd1 vssd1 vccd1 vccd1 _15334_/X sky130_fd_sc_hd__or2_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12546_ _20876_/Q _12548_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12550_/D sky130_fd_sc_hd__and3_1
X_18053_ _20757_/Q _20756_/Q _18053_/C vssd1 vssd1 vccd1 vccd1 _18055_/B sky130_fd_sc_hd__and3_2
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15265_ _14837_/S _15262_/Y _15263_/Y _10885_/B _15260_/X vssd1 vssd1 vccd1 vccd1
+ _15265_/X sky130_fd_sc_hd__o221a_1
X_12477_ _14895_/A _12468_/C _12500_/D _12480_/A vssd1 vssd1 vccd1 vccd1 _12477_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_4 _15238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ _20428_/Q _17004_/A2 _17004_/B1 vssd1 vssd1 vccd1 vccd1 _17004_/X sky130_fd_sc_hd__a21o_1
X_14216_ _20276_/Q _14117_/A _14216_/B1 input216/X vssd1 vssd1 vccd1 vccd1 _14218_/B
+ sky130_fd_sc_hd__a22o_4
XFILLER_160_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11428_ _19946_/Q _12131_/B vssd1 vssd1 vccd1 vccd1 _11428_/X sky130_fd_sc_hd__or2_1
X_15196_ _20853_/Q _15195_/X _15601_/S vssd1 vssd1 vccd1 vccd1 _15196_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11359_ _11357_/X _11358_/X _11359_/S vssd1 vssd1 vccd1 vccd1 _11359_/X sky130_fd_sc_hd__mux2_1
X_14147_ _19497_/Q _14148_/B vssd1 vssd1 vccd1 vccd1 _14161_/A sky130_fd_sc_hd__nor2_1
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_259_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14078_ _19198_/Q _14104_/A2 _14077_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1 _19198_/D
+ sky130_fd_sc_hd__o211a_1
X_18955_ _18955_/A _18955_/B vssd1 vssd1 vccd1 vccd1 _18955_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17906_ _20677_/Q _17906_/A1 _17914_/S vssd1 vssd1 vccd1 vccd1 _20677_/D sky130_fd_sc_hd__mux2_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13029_ _20964_/Q _20898_/Q vssd1 vssd1 vccd1 vccd1 _13029_/Y sky130_fd_sc_hd__nor2_2
X_18886_ _18975_/A _18886_/B vssd1 vssd1 vccd1 vccd1 _18886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_267_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1060 _10813_/X vssd1 vssd1 vccd1 vccd1 _17891_/A1 sky130_fd_sc_hd__buf_2
XFILLER_239_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1071 _09748_/Y vssd1 vssd1 vccd1 vccd1 _12433_/A1 sky130_fd_sc_hd__buf_6
X_17837_ _20612_/Q _17909_/A1 _17842_/S vssd1 vssd1 vccd1 vccd1 _20612_/D sky130_fd_sc_hd__mux2_1
Xfanout1082 _15326_/A vssd1 vssd1 vccd1 vccd1 _15527_/B sky130_fd_sc_hd__buf_2
Xfanout1093 _17706_/A1 vssd1 vssd1 vccd1 vccd1 _17881_/A1 sky130_fd_sc_hd__clkbuf_2
XFILLER_227_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_254_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17768_ _20547_/Q _17908_/A1 _17772_/S vssd1 vssd1 vccd1 vccd1 _20547_/D sky130_fd_sc_hd__mux2_1
XFILLER_214_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_282_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_270_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16719_ _16719_/A _16719_/B _16720_/D _12959_/B vssd1 vssd1 vccd1 vccd1 _16719_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19507_ _20930_/CLK _19507_/D vssd1 vssd1 vccd1 vccd1 _19507_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17699_ _20483_/Q _17802_/A1 _17703_/S vssd1 vssd1 vccd1 vccd1 _20483_/D sky130_fd_sc_hd__mux2_1
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_223_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19438_ _20718_/CLK _19438_/D vssd1 vssd1 vccd1 vccd1 _19438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19369_ _20657_/CLK _19369_/D vssd1 vssd1 vccd1 vccd1 _19369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20213_ _20766_/CLK _20213_/D vssd1 vssd1 vccd1 vccd1 _20213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_278_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_278_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_249_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20144_ _20579_/CLK _20144_/D vssd1 vssd1 vccd1 vccd1 _20144_/Q sky130_fd_sc_hd__dfxtp_1
X_09955_ _20481_/Q _20321_/Q _11899_/S vssd1 vssd1 vccd1 vccd1 _09955_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20075_ _20075_/CLK _20075_/D vssd1 vssd1 vccd1 vccd1 _20075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09886_ _09878_/X _09879_/X _11902_/S vssd1 vssd1 vccd1 vccd1 _09886_/X sky130_fd_sc_hd__mux2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_405 _16943_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_416 _18565_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_427 _12328_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_260_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_226_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_438 _13721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20977_ _21006_/CLK _20977_/D vssd1 vssd1 vccd1 vccd1 _20977_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_449 _13775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10730_ _19871_/Q _19772_/Q _12397_/S vssd1 vssd1 vccd1 vccd1 _10730_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_281_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10661_ _10659_/X _10660_/X _12391_/S vssd1 vssd1 vccd1 vccd1 _10662_/B sky130_fd_sc_hd__mux2_1
XFILLER_241_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12400_ _12400_/A1 _12392_/X _12399_/X _12385_/X vssd1 vssd1 vccd1 vccd1 _12400_/X
+ sky130_fd_sc_hd__o31a_4
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13380_ _14110_/B _13403_/B _13378_/Y _13379_/Y vssd1 vssd1 vccd1 vccd1 _13380_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_178_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10592_ _11995_/S _10590_/X _10591_/X _11684_/A1 vssd1 vssd1 vccd1 vccd1 _10592_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_222_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _12332_/A _19928_/Q _12334_/S0 _20053_/Q vssd1 vssd1 vccd1 vccd1 _12331_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_163_wb_clk_i clkbuf_4_5__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _20913_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12262_ _19427_/Q _20586_/Q _12428_/S vssd1 vssd1 vccd1 vccd1 _12262_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15050_ _15042_/X _15049_/X _15407_/S vssd1 vssd1 vccd1 vccd1 _15050_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14001_ _12504_/A _14043_/A2 _14040_/B1 _14000_/X _14088_/C1 vssd1 vssd1 vccd1 vccd1
+ _19167_/D sky130_fd_sc_hd__o221a_1
X_11213_ _20302_/Q _11213_/B vssd1 vssd1 vccd1 vccd1 _11213_/X sky130_fd_sc_hd__or2_1
X_12193_ _12012_/S _12168_/X _12176_/X _12192_/X vssd1 vssd1 vccd1 vccd1 _12193_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11144_ _14524_/B1 _16071_/A _11143_/Y vssd1 vssd1 vccd1 vccd1 _11144_/X sky130_fd_sc_hd__o21a_1
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18740_ _18740_/A _18740_/B vssd1 vssd1 vccd1 vccd1 _20970_/D sky130_fd_sc_hd__and2_1
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11075_ _11073_/X _11074_/X _12376_/S vssd1 vssd1 vccd1 vccd1 _11075_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15952_ _16007_/A _15952_/B vssd1 vssd1 vccd1 vccd1 _15952_/Y sky130_fd_sc_hd__nand2_1
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput130 dout1[30] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__clkbuf_2
XFILLER_283_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput141 dout1[40] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__buf_2
Xinput152 dout1[50] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__buf_2
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10026_ _11228_/A1 _09664_/B _10025_/X _11239_/B1 _19843_/Q vssd1 vssd1 vccd1 vccd1
+ _10026_/X sky130_fd_sc_hd__o32a_1
X_14903_ _18198_/B _18152_/B _16133_/C _16878_/A vssd1 vssd1 vccd1 vccd1 _14903_/Y
+ sky130_fd_sc_hd__a31oi_4
Xinput163 dout1[60] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_hd__clkbuf_2
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18671_ _19521_/Q _18671_/B vssd1 vssd1 vccd1 vccd1 _18671_/Y sky130_fd_sc_hd__nand2_1
XFILLER_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15883_ _15973_/A1 _15882_/X _15870_/X vssd1 vssd1 vccd1 vccd1 _15883_/X sky130_fd_sc_hd__a21o_1
XFILLER_237_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 irq[12] vssd1 vssd1 vccd1 vccd1 _12542_/C sky130_fd_sc_hd__clkbuf_2
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput185 irq[8] vssd1 vssd1 vccd1 vccd1 _12537_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_237_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput196 localMemory_wb_adr_i[15] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_hd__clkbuf_2
X_17622_ _20378_/Q _17933_/A1 _17623_/S vssd1 vssd1 vccd1 vccd1 _20378_/D sky130_fd_sc_hd__mux2_1
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ _11136_/B _12282_/B _14837_/S vssd1 vssd1 vccd1 vccd1 _14834_/X sky130_fd_sc_hd__mux2_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ _20313_/Q _17689_/A1 _17570_/S vssd1 vssd1 vccd1 vccd1 _20313_/D sky130_fd_sc_hd__mux2_1
XFILLER_251_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _19507_/Q _14773_/B vssd1 vssd1 vccd1 vccd1 _14765_/X sky130_fd_sc_hd__or2_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11977_ _11977_/A1 _19457_/Q _11979_/S _11976_/X vssd1 vssd1 vccd1 vccd1 _11977_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_204_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16504_ _19811_/Q _17097_/A1 _16521_/S vssd1 vssd1 vccd1 vccd1 _19811_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_260_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13716_ _16598_/C _13716_/B vssd1 vssd1 vccd1 vccd1 _13716_/Y sky130_fd_sc_hd__nor2_1
X_17484_ _20277_/Q _17486_/B vssd1 vssd1 vccd1 vccd1 _17484_/Y sky130_fd_sc_hd__nand2_1
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10928_ _11012_/A _10928_/B _10928_/C vssd1 vssd1 vccd1 vccd1 _10928_/X sky130_fd_sc_hd__or3_4
XFILLER_220_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14696_ _19455_/Q _17911_/A1 _14698_/S vssd1 vssd1 vccd1 vccd1 _19455_/D sky130_fd_sc_hd__mux2_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19223_ _19223_/CLK _19223_/D vssd1 vssd1 vccd1 vccd1 _19223_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_177_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16435_ _18863_/A _16435_/B _16437_/B vssd1 vssd1 vccd1 vccd1 _19758_/D sky130_fd_sc_hd__nor3_1
XFILLER_189_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13647_ _13663_/A _13663_/B _13676_/B vssd1 vssd1 vccd1 vccd1 _13647_/X sky130_fd_sc_hd__and3_4
X_10859_ _19371_/Q _12412_/A2 _10857_/X _12412_/B2 _10858_/X vssd1 vssd1 vccd1 vccd1
+ _10859_/X sky130_fd_sc_hd__o221a_1
XFILLER_220_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_258_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19154_ _19574_/CLK _19154_/D vssd1 vssd1 vccd1 vccd1 _19154_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_188_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16370_/C _16366_/B vssd1 vssd1 vccd1 vccd1 _19732_/D sky130_fd_sc_hd__nor2_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13047_/X _13048_/Y _13066_/X _13564_/B vssd1 vssd1 vccd1 vccd1 _13578_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18105_ _20776_/Q _18103_/B _18104_/Y vssd1 vssd1 vccd1 vccd1 _20776_/D sky130_fd_sc_hd__o21a_1
X_15317_ _15012_/B _14977_/Y _14978_/Y input7/X _15316_/X vssd1 vssd1 vccd1 vccd1
+ _15317_/X sky130_fd_sc_hd__o221a_1
XFILLER_173_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19085_ _19620_/CLK _19085_/D vssd1 vssd1 vccd1 vccd1 _19085_/Q sky130_fd_sc_hd__dfxtp_2
X_12529_ _12527_/X _12528_/X _18476_/A vssd1 vssd1 vccd1 vccd1 _12529_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16297_ _19707_/Q _16300_/C vssd1 vssd1 vccd1 vccd1 _16298_/B sky130_fd_sc_hd__and2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_258_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18036_ _20751_/Q _20750_/Q _18036_/C vssd1 vssd1 vccd1 vccd1 _18039_/B sky130_fd_sc_hd__and3_2
XFILLER_184_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15248_ _15248_/A _15248_/B _15248_/C vssd1 vssd1 vccd1 vccd1 _15248_/X sky130_fd_sc_hd__and3_1
X_15179_ _11053_/Y _15500_/A0 _15178_/Y _11055_/B vssd1 vssd1 vccd1 vccd1 _15179_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_259_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19987_ _19992_/CLK _19987_/D vssd1 vssd1 vccd1 vccd1 _19987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09740_ _16454_/B _12426_/S vssd1 vssd1 vccd1 vccd1 _09746_/A sky130_fd_sc_hd__xnor2_1
X_18938_ _18541_/X _18964_/B _18936_/X _18937_/Y vssd1 vssd1 vccd1 vccd1 _18939_/B
+ sky130_fd_sc_hd__o211a_1
.ends

