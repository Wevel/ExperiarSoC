magic
tech sky130A
magscale 1 2
timestamp 1683814369
<< obsli1 >>
rect 1104 2159 68816 217617
<< obsm1 >>
rect 14 892 69078 219292
<< metal2 >>
rect 3698 219200 3754 220000
rect 4342 219200 4398 220000
rect 4986 219200 5042 220000
rect 5630 219200 5686 220000
rect 6274 219200 6330 220000
rect 6918 219200 6974 220000
rect 7562 219200 7618 220000
rect 8206 219200 8262 220000
rect 8850 219200 8906 220000
rect 9494 219200 9550 220000
rect 10138 219200 10194 220000
rect 10782 219200 10838 220000
rect 11426 219200 11482 220000
rect 12070 219200 12126 220000
rect 12714 219200 12770 220000
rect 13358 219200 13414 220000
rect 14002 219200 14058 220000
rect 14646 219200 14702 220000
rect 15290 219200 15346 220000
rect 15934 219200 15990 220000
rect 16578 219200 16634 220000
rect 17222 219200 17278 220000
rect 17866 219200 17922 220000
rect 18510 219200 18566 220000
rect 19154 219200 19210 220000
rect 19798 219200 19854 220000
rect 20442 219200 20498 220000
rect 21086 219200 21142 220000
rect 21730 219200 21786 220000
rect 22374 219200 22430 220000
rect 23018 219200 23074 220000
rect 23662 219200 23718 220000
rect 24306 219200 24362 220000
rect 24950 219200 25006 220000
rect 25594 219200 25650 220000
rect 26238 219200 26294 220000
rect 26882 219200 26938 220000
rect 27526 219200 27582 220000
rect 28170 219200 28226 220000
rect 28814 219200 28870 220000
rect 29458 219200 29514 220000
rect 30102 219200 30158 220000
rect 30746 219200 30802 220000
rect 31390 219200 31446 220000
rect 32034 219200 32090 220000
rect 32678 219200 32734 220000
rect 33322 219200 33378 220000
rect 33966 219200 34022 220000
rect 34610 219200 34666 220000
rect 35254 219200 35310 220000
rect 35898 219200 35954 220000
rect 36542 219200 36598 220000
rect 37186 219200 37242 220000
rect 37830 219200 37886 220000
rect 38474 219200 38530 220000
rect 39118 219200 39174 220000
rect 39762 219200 39818 220000
rect 40406 219200 40462 220000
rect 41050 219200 41106 220000
rect 41694 219200 41750 220000
rect 42338 219200 42394 220000
rect 42982 219200 43038 220000
rect 43626 219200 43682 220000
rect 44270 219200 44326 220000
rect 44914 219200 44970 220000
rect 45558 219200 45614 220000
rect 46202 219200 46258 220000
rect 46846 219200 46902 220000
rect 47490 219200 47546 220000
rect 48134 219200 48190 220000
rect 48778 219200 48834 220000
rect 49422 219200 49478 220000
rect 50066 219200 50122 220000
rect 50710 219200 50766 220000
rect 51354 219200 51410 220000
rect 51998 219200 52054 220000
rect 52642 219200 52698 220000
rect 53286 219200 53342 220000
rect 53930 219200 53986 220000
rect 54574 219200 54630 220000
rect 55218 219200 55274 220000
rect 55862 219200 55918 220000
rect 56506 219200 56562 220000
rect 57150 219200 57206 220000
rect 57794 219200 57850 220000
rect 58438 219200 58494 220000
rect 59082 219200 59138 220000
rect 59726 219200 59782 220000
rect 60370 219200 60426 220000
rect 61014 219200 61070 220000
rect 61658 219200 61714 220000
rect 62302 219200 62358 220000
rect 62946 219200 63002 220000
rect 63590 219200 63646 220000
rect 64234 219200 64290 220000
rect 64878 219200 64934 220000
rect 65522 219200 65578 220000
rect 66166 219200 66222 220000
rect 2134 0 2190 800
rect 2686 0 2742 800
rect 3238 0 3294 800
rect 3790 0 3846 800
rect 4342 0 4398 800
rect 4894 0 4950 800
rect 5446 0 5502 800
rect 5998 0 6054 800
rect 6550 0 6606 800
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8206 0 8262 800
rect 8758 0 8814 800
rect 9310 0 9366 800
rect 9862 0 9918 800
rect 10414 0 10470 800
rect 10966 0 11022 800
rect 11518 0 11574 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17590 0 17646 800
rect 18142 0 18198 800
rect 18694 0 18750 800
rect 19246 0 19302 800
rect 19798 0 19854 800
rect 20350 0 20406 800
rect 20902 0 20958 800
rect 21454 0 21510 800
rect 22006 0 22062 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23662 0 23718 800
rect 24214 0 24270 800
rect 24766 0 24822 800
rect 25318 0 25374 800
rect 25870 0 25926 800
rect 26422 0 26478 800
rect 26974 0 27030 800
rect 27526 0 27582 800
rect 28078 0 28134 800
rect 28630 0 28686 800
rect 29182 0 29238 800
rect 29734 0 29790 800
rect 30286 0 30342 800
rect 30838 0 30894 800
rect 31390 0 31446 800
rect 31942 0 31998 800
rect 32494 0 32550 800
rect 33046 0 33102 800
rect 33598 0 33654 800
rect 34150 0 34206 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36358 0 36414 800
rect 36910 0 36966 800
rect 37462 0 37518 800
rect 38014 0 38070 800
rect 38566 0 38622 800
rect 39118 0 39174 800
rect 39670 0 39726 800
rect 40222 0 40278 800
rect 40774 0 40830 800
rect 41326 0 41382 800
rect 41878 0 41934 800
rect 42430 0 42486 800
rect 42982 0 43038 800
rect 43534 0 43590 800
rect 44086 0 44142 800
rect 44638 0 44694 800
rect 45190 0 45246 800
rect 45742 0 45798 800
rect 46294 0 46350 800
rect 46846 0 46902 800
rect 47398 0 47454 800
rect 47950 0 48006 800
rect 48502 0 48558 800
rect 49054 0 49110 800
rect 49606 0 49662 800
rect 50158 0 50214 800
rect 50710 0 50766 800
rect 51262 0 51318 800
rect 51814 0 51870 800
rect 52366 0 52422 800
rect 52918 0 52974 800
rect 53470 0 53526 800
rect 54022 0 54078 800
rect 54574 0 54630 800
rect 55126 0 55182 800
rect 55678 0 55734 800
rect 56230 0 56286 800
rect 56782 0 56838 800
rect 57334 0 57390 800
rect 57886 0 57942 800
rect 58438 0 58494 800
rect 58990 0 59046 800
rect 59542 0 59598 800
rect 60094 0 60150 800
rect 60646 0 60702 800
rect 61198 0 61254 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62854 0 62910 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64510 0 64566 800
rect 65062 0 65118 800
rect 65614 0 65670 800
rect 66166 0 66222 800
rect 66718 0 66774 800
rect 67270 0 67326 800
rect 67822 0 67878 800
<< obsm2 >>
rect 20 219144 3642 219450
rect 3810 219144 4286 219450
rect 4454 219144 4930 219450
rect 5098 219144 5574 219450
rect 5742 219144 6218 219450
rect 6386 219144 6862 219450
rect 7030 219144 7506 219450
rect 7674 219144 8150 219450
rect 8318 219144 8794 219450
rect 8962 219144 9438 219450
rect 9606 219144 10082 219450
rect 10250 219144 10726 219450
rect 10894 219144 11370 219450
rect 11538 219144 12014 219450
rect 12182 219144 12658 219450
rect 12826 219144 13302 219450
rect 13470 219144 13946 219450
rect 14114 219144 14590 219450
rect 14758 219144 15234 219450
rect 15402 219144 15878 219450
rect 16046 219144 16522 219450
rect 16690 219144 17166 219450
rect 17334 219144 17810 219450
rect 17978 219144 18454 219450
rect 18622 219144 19098 219450
rect 19266 219144 19742 219450
rect 19910 219144 20386 219450
rect 20554 219144 21030 219450
rect 21198 219144 21674 219450
rect 21842 219144 22318 219450
rect 22486 219144 22962 219450
rect 23130 219144 23606 219450
rect 23774 219144 24250 219450
rect 24418 219144 24894 219450
rect 25062 219144 25538 219450
rect 25706 219144 26182 219450
rect 26350 219144 26826 219450
rect 26994 219144 27470 219450
rect 27638 219144 28114 219450
rect 28282 219144 28758 219450
rect 28926 219144 29402 219450
rect 29570 219144 30046 219450
rect 30214 219144 30690 219450
rect 30858 219144 31334 219450
rect 31502 219144 31978 219450
rect 32146 219144 32622 219450
rect 32790 219144 33266 219450
rect 33434 219144 33910 219450
rect 34078 219144 34554 219450
rect 34722 219144 35198 219450
rect 35366 219144 35842 219450
rect 36010 219144 36486 219450
rect 36654 219144 37130 219450
rect 37298 219144 37774 219450
rect 37942 219144 38418 219450
rect 38586 219144 39062 219450
rect 39230 219144 39706 219450
rect 39874 219144 40350 219450
rect 40518 219144 40994 219450
rect 41162 219144 41638 219450
rect 41806 219144 42282 219450
rect 42450 219144 42926 219450
rect 43094 219144 43570 219450
rect 43738 219144 44214 219450
rect 44382 219144 44858 219450
rect 45026 219144 45502 219450
rect 45670 219144 46146 219450
rect 46314 219144 46790 219450
rect 46958 219144 47434 219450
rect 47602 219144 48078 219450
rect 48246 219144 48722 219450
rect 48890 219144 49366 219450
rect 49534 219144 50010 219450
rect 50178 219144 50654 219450
rect 50822 219144 51298 219450
rect 51466 219144 51942 219450
rect 52110 219144 52586 219450
rect 52754 219144 53230 219450
rect 53398 219144 53874 219450
rect 54042 219144 54518 219450
rect 54686 219144 55162 219450
rect 55330 219144 55806 219450
rect 55974 219144 56450 219450
rect 56618 219144 57094 219450
rect 57262 219144 57738 219450
rect 57906 219144 58382 219450
rect 58550 219144 59026 219450
rect 59194 219144 59670 219450
rect 59838 219144 60314 219450
rect 60482 219144 60958 219450
rect 61126 219144 61602 219450
rect 61770 219144 62246 219450
rect 62414 219144 62890 219450
rect 63058 219144 63534 219450
rect 63702 219144 64178 219450
rect 64346 219144 64822 219450
rect 64990 219144 65466 219450
rect 65634 219144 66110 219450
rect 66278 219144 69074 219450
rect 20 856 69074 219144
rect 20 734 2078 856
rect 2246 734 2630 856
rect 2798 734 3182 856
rect 3350 734 3734 856
rect 3902 734 4286 856
rect 4454 734 4838 856
rect 5006 734 5390 856
rect 5558 734 5942 856
rect 6110 734 6494 856
rect 6662 734 7046 856
rect 7214 734 7598 856
rect 7766 734 8150 856
rect 8318 734 8702 856
rect 8870 734 9254 856
rect 9422 734 9806 856
rect 9974 734 10358 856
rect 10526 734 10910 856
rect 11078 734 11462 856
rect 11630 734 12014 856
rect 12182 734 12566 856
rect 12734 734 13118 856
rect 13286 734 13670 856
rect 13838 734 14222 856
rect 14390 734 14774 856
rect 14942 734 15326 856
rect 15494 734 15878 856
rect 16046 734 16430 856
rect 16598 734 16982 856
rect 17150 734 17534 856
rect 17702 734 18086 856
rect 18254 734 18638 856
rect 18806 734 19190 856
rect 19358 734 19742 856
rect 19910 734 20294 856
rect 20462 734 20846 856
rect 21014 734 21398 856
rect 21566 734 21950 856
rect 22118 734 22502 856
rect 22670 734 23054 856
rect 23222 734 23606 856
rect 23774 734 24158 856
rect 24326 734 24710 856
rect 24878 734 25262 856
rect 25430 734 25814 856
rect 25982 734 26366 856
rect 26534 734 26918 856
rect 27086 734 27470 856
rect 27638 734 28022 856
rect 28190 734 28574 856
rect 28742 734 29126 856
rect 29294 734 29678 856
rect 29846 734 30230 856
rect 30398 734 30782 856
rect 30950 734 31334 856
rect 31502 734 31886 856
rect 32054 734 32438 856
rect 32606 734 32990 856
rect 33158 734 33542 856
rect 33710 734 34094 856
rect 34262 734 34646 856
rect 34814 734 35198 856
rect 35366 734 35750 856
rect 35918 734 36302 856
rect 36470 734 36854 856
rect 37022 734 37406 856
rect 37574 734 37958 856
rect 38126 734 38510 856
rect 38678 734 39062 856
rect 39230 734 39614 856
rect 39782 734 40166 856
rect 40334 734 40718 856
rect 40886 734 41270 856
rect 41438 734 41822 856
rect 41990 734 42374 856
rect 42542 734 42926 856
rect 43094 734 43478 856
rect 43646 734 44030 856
rect 44198 734 44582 856
rect 44750 734 45134 856
rect 45302 734 45686 856
rect 45854 734 46238 856
rect 46406 734 46790 856
rect 46958 734 47342 856
rect 47510 734 47894 856
rect 48062 734 48446 856
rect 48614 734 48998 856
rect 49166 734 49550 856
rect 49718 734 50102 856
rect 50270 734 50654 856
rect 50822 734 51206 856
rect 51374 734 51758 856
rect 51926 734 52310 856
rect 52478 734 52862 856
rect 53030 734 53414 856
rect 53582 734 53966 856
rect 54134 734 54518 856
rect 54686 734 55070 856
rect 55238 734 55622 856
rect 55790 734 56174 856
rect 56342 734 56726 856
rect 56894 734 57278 856
rect 57446 734 57830 856
rect 57998 734 58382 856
rect 58550 734 58934 856
rect 59102 734 59486 856
rect 59654 734 60038 856
rect 60206 734 60590 856
rect 60758 734 61142 856
rect 61310 734 61694 856
rect 61862 734 62246 856
rect 62414 734 62798 856
rect 62966 734 63350 856
rect 63518 734 63902 856
rect 64070 734 64454 856
rect 64622 734 65006 856
rect 65174 734 65558 856
rect 65726 734 66110 856
rect 66278 734 66662 856
rect 66830 734 67214 856
rect 67382 734 67766 856
rect 67934 734 69074 856
<< metal3 >>
rect 0 218424 800 218544
rect 0 217880 800 218000
rect 0 217336 800 217456
rect 0 216792 800 216912
rect 0 216248 800 216368
rect 69200 215976 70000 216096
rect 0 215704 800 215824
rect 0 215160 800 215280
rect 69200 214888 70000 215008
rect 0 214616 800 214736
rect 0 214072 800 214192
rect 69200 213800 70000 213920
rect 0 213528 800 213648
rect 0 212984 800 213104
rect 69200 212712 70000 212832
rect 0 212440 800 212560
rect 0 211896 800 212016
rect 69200 211624 70000 211744
rect 0 211352 800 211472
rect 0 210808 800 210928
rect 69200 210536 70000 210656
rect 0 210264 800 210384
rect 0 209720 800 209840
rect 69200 209448 70000 209568
rect 0 209176 800 209296
rect 0 208632 800 208752
rect 69200 208360 70000 208480
rect 0 208088 800 208208
rect 0 207544 800 207664
rect 69200 207272 70000 207392
rect 0 207000 800 207120
rect 0 206456 800 206576
rect 69200 206184 70000 206304
rect 0 205912 800 206032
rect 0 205368 800 205488
rect 69200 205096 70000 205216
rect 0 204824 800 204944
rect 0 204280 800 204400
rect 69200 204008 70000 204128
rect 0 203736 800 203856
rect 0 203192 800 203312
rect 69200 202920 70000 203040
rect 0 202648 800 202768
rect 0 202104 800 202224
rect 69200 201832 70000 201952
rect 0 201560 800 201680
rect 0 201016 800 201136
rect 69200 200744 70000 200864
rect 0 200472 800 200592
rect 0 199928 800 200048
rect 69200 199656 70000 199776
rect 0 199384 800 199504
rect 0 198840 800 198960
rect 69200 198568 70000 198688
rect 0 198296 800 198416
rect 0 197752 800 197872
rect 69200 197480 70000 197600
rect 0 197208 800 197328
rect 0 196664 800 196784
rect 69200 196392 70000 196512
rect 0 196120 800 196240
rect 0 195576 800 195696
rect 69200 195304 70000 195424
rect 0 195032 800 195152
rect 0 194488 800 194608
rect 69200 194216 70000 194336
rect 0 193944 800 194064
rect 0 193400 800 193520
rect 69200 193128 70000 193248
rect 0 192856 800 192976
rect 0 192312 800 192432
rect 69200 192040 70000 192160
rect 0 191768 800 191888
rect 0 191224 800 191344
rect 69200 190952 70000 191072
rect 0 190680 800 190800
rect 0 190136 800 190256
rect 69200 189864 70000 189984
rect 0 189592 800 189712
rect 0 189048 800 189168
rect 69200 188776 70000 188896
rect 0 188504 800 188624
rect 0 187960 800 188080
rect 69200 187688 70000 187808
rect 0 187416 800 187536
rect 0 186872 800 186992
rect 69200 186600 70000 186720
rect 0 186328 800 186448
rect 0 185784 800 185904
rect 69200 185512 70000 185632
rect 0 185240 800 185360
rect 0 184696 800 184816
rect 69200 184424 70000 184544
rect 0 184152 800 184272
rect 0 183608 800 183728
rect 69200 183336 70000 183456
rect 0 183064 800 183184
rect 0 182520 800 182640
rect 69200 182248 70000 182368
rect 0 181976 800 182096
rect 0 181432 800 181552
rect 69200 181160 70000 181280
rect 0 180888 800 181008
rect 0 180344 800 180464
rect 69200 180072 70000 180192
rect 0 179800 800 179920
rect 0 179256 800 179376
rect 69200 178984 70000 179104
rect 0 178712 800 178832
rect 0 178168 800 178288
rect 69200 177896 70000 178016
rect 0 177624 800 177744
rect 0 177080 800 177200
rect 69200 176808 70000 176928
rect 0 176536 800 176656
rect 0 175992 800 176112
rect 69200 175720 70000 175840
rect 0 175448 800 175568
rect 0 174904 800 175024
rect 69200 174632 70000 174752
rect 0 174360 800 174480
rect 0 173816 800 173936
rect 69200 173544 70000 173664
rect 0 173272 800 173392
rect 0 172728 800 172848
rect 69200 172456 70000 172576
rect 0 172184 800 172304
rect 0 171640 800 171760
rect 69200 171368 70000 171488
rect 0 171096 800 171216
rect 0 170552 800 170672
rect 69200 170280 70000 170400
rect 0 170008 800 170128
rect 0 169464 800 169584
rect 69200 169192 70000 169312
rect 0 168920 800 169040
rect 0 168376 800 168496
rect 69200 168104 70000 168224
rect 0 167832 800 167952
rect 0 167288 800 167408
rect 69200 167016 70000 167136
rect 0 166744 800 166864
rect 0 166200 800 166320
rect 69200 165928 70000 166048
rect 0 165656 800 165776
rect 0 165112 800 165232
rect 69200 164840 70000 164960
rect 0 164568 800 164688
rect 0 164024 800 164144
rect 69200 163752 70000 163872
rect 0 163480 800 163600
rect 0 162936 800 163056
rect 69200 162664 70000 162784
rect 0 162392 800 162512
rect 0 161848 800 161968
rect 69200 161576 70000 161696
rect 0 161304 800 161424
rect 0 160760 800 160880
rect 69200 160488 70000 160608
rect 0 160216 800 160336
rect 0 159672 800 159792
rect 69200 159400 70000 159520
rect 0 159128 800 159248
rect 0 158584 800 158704
rect 69200 158312 70000 158432
rect 0 158040 800 158160
rect 0 157496 800 157616
rect 69200 157224 70000 157344
rect 0 156952 800 157072
rect 0 156408 800 156528
rect 69200 156136 70000 156256
rect 0 155864 800 155984
rect 0 155320 800 155440
rect 69200 155048 70000 155168
rect 0 154776 800 154896
rect 0 154232 800 154352
rect 69200 153960 70000 154080
rect 0 153688 800 153808
rect 0 153144 800 153264
rect 69200 152872 70000 152992
rect 0 152600 800 152720
rect 0 152056 800 152176
rect 69200 151784 70000 151904
rect 0 151512 800 151632
rect 0 150968 800 151088
rect 69200 150696 70000 150816
rect 0 150424 800 150544
rect 0 149880 800 150000
rect 69200 149608 70000 149728
rect 0 149336 800 149456
rect 0 148792 800 148912
rect 69200 148520 70000 148640
rect 0 148248 800 148368
rect 0 147704 800 147824
rect 69200 147432 70000 147552
rect 0 147160 800 147280
rect 0 146616 800 146736
rect 69200 146344 70000 146464
rect 0 146072 800 146192
rect 0 145528 800 145648
rect 69200 145256 70000 145376
rect 0 144984 800 145104
rect 0 144440 800 144560
rect 69200 144168 70000 144288
rect 0 143896 800 144016
rect 0 143352 800 143472
rect 69200 143080 70000 143200
rect 0 142808 800 142928
rect 0 142264 800 142384
rect 69200 141992 70000 142112
rect 0 141720 800 141840
rect 0 141176 800 141296
rect 69200 140904 70000 141024
rect 0 140632 800 140752
rect 0 140088 800 140208
rect 69200 139816 70000 139936
rect 0 139544 800 139664
rect 0 139000 800 139120
rect 69200 138728 70000 138848
rect 0 138456 800 138576
rect 0 137912 800 138032
rect 69200 137640 70000 137760
rect 0 137368 800 137488
rect 0 136824 800 136944
rect 69200 136552 70000 136672
rect 0 136280 800 136400
rect 0 135736 800 135856
rect 69200 135464 70000 135584
rect 0 135192 800 135312
rect 0 134648 800 134768
rect 69200 134376 70000 134496
rect 0 134104 800 134224
rect 0 133560 800 133680
rect 69200 133288 70000 133408
rect 0 133016 800 133136
rect 0 132472 800 132592
rect 69200 132200 70000 132320
rect 0 131928 800 132048
rect 0 131384 800 131504
rect 69200 131112 70000 131232
rect 0 130840 800 130960
rect 0 130296 800 130416
rect 69200 130024 70000 130144
rect 0 129752 800 129872
rect 0 129208 800 129328
rect 69200 128936 70000 129056
rect 0 128664 800 128784
rect 0 128120 800 128240
rect 69200 127848 70000 127968
rect 0 127576 800 127696
rect 0 127032 800 127152
rect 69200 126760 70000 126880
rect 0 126488 800 126608
rect 0 125944 800 126064
rect 69200 125672 70000 125792
rect 0 125400 800 125520
rect 0 124856 800 124976
rect 69200 124584 70000 124704
rect 0 124312 800 124432
rect 0 123768 800 123888
rect 69200 123496 70000 123616
rect 0 123224 800 123344
rect 0 122680 800 122800
rect 69200 122408 70000 122528
rect 0 122136 800 122256
rect 0 121592 800 121712
rect 69200 121320 70000 121440
rect 0 121048 800 121168
rect 0 120504 800 120624
rect 69200 120232 70000 120352
rect 0 119960 800 120080
rect 0 119416 800 119536
rect 69200 119144 70000 119264
rect 0 118872 800 118992
rect 0 118328 800 118448
rect 69200 118056 70000 118176
rect 0 117784 800 117904
rect 0 117240 800 117360
rect 69200 116968 70000 117088
rect 0 116696 800 116816
rect 0 116152 800 116272
rect 69200 115880 70000 116000
rect 0 115608 800 115728
rect 0 115064 800 115184
rect 69200 114792 70000 114912
rect 0 114520 800 114640
rect 0 113976 800 114096
rect 69200 113704 70000 113824
rect 0 113432 800 113552
rect 0 112888 800 113008
rect 69200 112616 70000 112736
rect 0 112344 800 112464
rect 0 111800 800 111920
rect 69200 111528 70000 111648
rect 0 111256 800 111376
rect 0 110712 800 110832
rect 69200 110440 70000 110560
rect 0 110168 800 110288
rect 0 109624 800 109744
rect 69200 109352 70000 109472
rect 0 109080 800 109200
rect 0 108536 800 108656
rect 69200 108264 70000 108384
rect 0 107992 800 108112
rect 0 107448 800 107568
rect 69200 107176 70000 107296
rect 0 106904 800 107024
rect 0 106360 800 106480
rect 69200 106088 70000 106208
rect 0 105816 800 105936
rect 0 105272 800 105392
rect 69200 105000 70000 105120
rect 0 104728 800 104848
rect 0 104184 800 104304
rect 69200 103912 70000 104032
rect 0 103640 800 103760
rect 0 103096 800 103216
rect 69200 102824 70000 102944
rect 0 102552 800 102672
rect 0 102008 800 102128
rect 69200 101736 70000 101856
rect 0 101464 800 101584
rect 0 100920 800 101040
rect 69200 100648 70000 100768
rect 0 100376 800 100496
rect 0 99832 800 99952
rect 69200 99560 70000 99680
rect 0 99288 800 99408
rect 0 98744 800 98864
rect 69200 98472 70000 98592
rect 0 98200 800 98320
rect 0 97656 800 97776
rect 69200 97384 70000 97504
rect 0 97112 800 97232
rect 0 96568 800 96688
rect 69200 96296 70000 96416
rect 0 96024 800 96144
rect 0 95480 800 95600
rect 69200 95208 70000 95328
rect 0 94936 800 95056
rect 0 94392 800 94512
rect 69200 94120 70000 94240
rect 0 93848 800 93968
rect 0 93304 800 93424
rect 69200 93032 70000 93152
rect 0 92760 800 92880
rect 0 92216 800 92336
rect 69200 91944 70000 92064
rect 0 91672 800 91792
rect 0 91128 800 91248
rect 69200 90856 70000 90976
rect 0 90584 800 90704
rect 0 90040 800 90160
rect 69200 89768 70000 89888
rect 0 89496 800 89616
rect 0 88952 800 89072
rect 69200 88680 70000 88800
rect 0 88408 800 88528
rect 0 87864 800 87984
rect 69200 87592 70000 87712
rect 0 87320 800 87440
rect 0 86776 800 86896
rect 69200 86504 70000 86624
rect 0 86232 800 86352
rect 0 85688 800 85808
rect 69200 85416 70000 85536
rect 0 85144 800 85264
rect 0 84600 800 84720
rect 69200 84328 70000 84448
rect 0 84056 800 84176
rect 0 83512 800 83632
rect 69200 83240 70000 83360
rect 0 82968 800 83088
rect 0 82424 800 82544
rect 69200 82152 70000 82272
rect 0 81880 800 82000
rect 0 81336 800 81456
rect 69200 81064 70000 81184
rect 0 80792 800 80912
rect 0 80248 800 80368
rect 69200 79976 70000 80096
rect 0 79704 800 79824
rect 0 79160 800 79280
rect 69200 78888 70000 79008
rect 0 78616 800 78736
rect 0 78072 800 78192
rect 69200 77800 70000 77920
rect 0 77528 800 77648
rect 0 76984 800 77104
rect 69200 76712 70000 76832
rect 0 76440 800 76560
rect 0 75896 800 76016
rect 69200 75624 70000 75744
rect 0 75352 800 75472
rect 0 74808 800 74928
rect 69200 74536 70000 74656
rect 0 74264 800 74384
rect 0 73720 800 73840
rect 69200 73448 70000 73568
rect 0 73176 800 73296
rect 0 72632 800 72752
rect 69200 72360 70000 72480
rect 0 72088 800 72208
rect 0 71544 800 71664
rect 69200 71272 70000 71392
rect 0 71000 800 71120
rect 0 70456 800 70576
rect 69200 70184 70000 70304
rect 0 69912 800 70032
rect 0 69368 800 69488
rect 69200 69096 70000 69216
rect 0 68824 800 68944
rect 0 68280 800 68400
rect 69200 68008 70000 68128
rect 0 67736 800 67856
rect 0 67192 800 67312
rect 69200 66920 70000 67040
rect 0 66648 800 66768
rect 0 66104 800 66224
rect 69200 65832 70000 65952
rect 0 65560 800 65680
rect 0 65016 800 65136
rect 69200 64744 70000 64864
rect 0 64472 800 64592
rect 0 63928 800 64048
rect 69200 63656 70000 63776
rect 0 63384 800 63504
rect 0 62840 800 62960
rect 69200 62568 70000 62688
rect 0 62296 800 62416
rect 0 61752 800 61872
rect 69200 61480 70000 61600
rect 0 61208 800 61328
rect 0 60664 800 60784
rect 69200 60392 70000 60512
rect 0 60120 800 60240
rect 0 59576 800 59696
rect 69200 59304 70000 59424
rect 0 59032 800 59152
rect 0 58488 800 58608
rect 69200 58216 70000 58336
rect 0 57944 800 58064
rect 0 57400 800 57520
rect 69200 57128 70000 57248
rect 0 56856 800 56976
rect 0 56312 800 56432
rect 69200 56040 70000 56160
rect 0 55768 800 55888
rect 0 55224 800 55344
rect 69200 54952 70000 55072
rect 0 54680 800 54800
rect 0 54136 800 54256
rect 69200 53864 70000 53984
rect 0 53592 800 53712
rect 0 53048 800 53168
rect 69200 52776 70000 52896
rect 0 52504 800 52624
rect 0 51960 800 52080
rect 69200 51688 70000 51808
rect 0 51416 800 51536
rect 0 50872 800 50992
rect 69200 50600 70000 50720
rect 0 50328 800 50448
rect 0 49784 800 49904
rect 69200 49512 70000 49632
rect 0 49240 800 49360
rect 0 48696 800 48816
rect 69200 48424 70000 48544
rect 0 48152 800 48272
rect 0 47608 800 47728
rect 69200 47336 70000 47456
rect 0 47064 800 47184
rect 0 46520 800 46640
rect 69200 46248 70000 46368
rect 0 45976 800 46096
rect 0 45432 800 45552
rect 69200 45160 70000 45280
rect 0 44888 800 45008
rect 0 44344 800 44464
rect 69200 44072 70000 44192
rect 0 43800 800 43920
rect 0 43256 800 43376
rect 69200 42984 70000 43104
rect 0 42712 800 42832
rect 0 42168 800 42288
rect 69200 41896 70000 42016
rect 0 41624 800 41744
rect 0 41080 800 41200
rect 69200 40808 70000 40928
rect 0 40536 800 40656
rect 0 39992 800 40112
rect 69200 39720 70000 39840
rect 0 39448 800 39568
rect 0 38904 800 39024
rect 69200 38632 70000 38752
rect 0 38360 800 38480
rect 0 37816 800 37936
rect 69200 37544 70000 37664
rect 0 37272 800 37392
rect 0 36728 800 36848
rect 69200 36456 70000 36576
rect 0 36184 800 36304
rect 0 35640 800 35760
rect 69200 35368 70000 35488
rect 0 35096 800 35216
rect 0 34552 800 34672
rect 69200 34280 70000 34400
rect 0 34008 800 34128
rect 0 33464 800 33584
rect 69200 33192 70000 33312
rect 0 32920 800 33040
rect 0 32376 800 32496
rect 69200 32104 70000 32224
rect 0 31832 800 31952
rect 0 31288 800 31408
rect 69200 31016 70000 31136
rect 0 30744 800 30864
rect 0 30200 800 30320
rect 69200 29928 70000 30048
rect 0 29656 800 29776
rect 0 29112 800 29232
rect 69200 28840 70000 28960
rect 0 28568 800 28688
rect 0 28024 800 28144
rect 69200 27752 70000 27872
rect 0 27480 800 27600
rect 0 26936 800 27056
rect 69200 26664 70000 26784
rect 0 26392 800 26512
rect 0 25848 800 25968
rect 69200 25576 70000 25696
rect 0 25304 800 25424
rect 0 24760 800 24880
rect 69200 24488 70000 24608
rect 0 24216 800 24336
rect 0 23672 800 23792
rect 69200 23400 70000 23520
rect 0 23128 800 23248
rect 0 22584 800 22704
rect 69200 22312 70000 22432
rect 0 22040 800 22160
rect 0 21496 800 21616
rect 69200 21224 70000 21344
rect 0 20952 800 21072
rect 0 20408 800 20528
rect 69200 20136 70000 20256
rect 0 19864 800 19984
rect 0 19320 800 19440
rect 69200 19048 70000 19168
rect 0 18776 800 18896
rect 0 18232 800 18352
rect 69200 17960 70000 18080
rect 0 17688 800 17808
rect 0 17144 800 17264
rect 69200 16872 70000 16992
rect 0 16600 800 16720
rect 0 16056 800 16176
rect 69200 15784 70000 15904
rect 0 15512 800 15632
rect 0 14968 800 15088
rect 69200 14696 70000 14816
rect 0 14424 800 14544
rect 0 13880 800 14000
rect 69200 13608 70000 13728
rect 0 13336 800 13456
rect 0 12792 800 12912
rect 69200 12520 70000 12640
rect 0 12248 800 12368
rect 0 11704 800 11824
rect 69200 11432 70000 11552
rect 0 11160 800 11280
rect 0 10616 800 10736
rect 69200 10344 70000 10464
rect 0 10072 800 10192
rect 0 9528 800 9648
rect 69200 9256 70000 9376
rect 0 8984 800 9104
rect 0 8440 800 8560
rect 69200 8168 70000 8288
rect 0 7896 800 8016
rect 0 7352 800 7472
rect 69200 7080 70000 7200
rect 0 6808 800 6928
rect 0 6264 800 6384
rect 69200 5992 70000 6112
rect 0 5720 800 5840
rect 0 5176 800 5296
rect 69200 4904 70000 5024
rect 0 4632 800 4752
rect 0 4088 800 4208
rect 69200 3816 70000 3936
rect 0 3544 800 3664
rect 0 3000 800 3120
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 0 1368 800 1488
<< obsm3 >>
rect 880 218344 69200 218517
rect 790 218080 69200 218344
rect 880 217800 69200 218080
rect 790 217536 69200 217800
rect 880 217256 69200 217536
rect 790 216992 69200 217256
rect 880 216712 69200 216992
rect 790 216448 69200 216712
rect 880 216176 69200 216448
rect 880 216168 69120 216176
rect 790 215904 69120 216168
rect 880 215896 69120 215904
rect 880 215624 69200 215896
rect 790 215360 69200 215624
rect 880 215088 69200 215360
rect 880 215080 69120 215088
rect 790 214816 69120 215080
rect 880 214808 69120 214816
rect 880 214536 69200 214808
rect 790 214272 69200 214536
rect 880 214000 69200 214272
rect 880 213992 69120 214000
rect 790 213728 69120 213992
rect 880 213720 69120 213728
rect 880 213448 69200 213720
rect 790 213184 69200 213448
rect 880 212912 69200 213184
rect 880 212904 69120 212912
rect 790 212640 69120 212904
rect 880 212632 69120 212640
rect 880 212360 69200 212632
rect 790 212096 69200 212360
rect 880 211824 69200 212096
rect 880 211816 69120 211824
rect 790 211552 69120 211816
rect 880 211544 69120 211552
rect 880 211272 69200 211544
rect 790 211008 69200 211272
rect 880 210736 69200 211008
rect 880 210728 69120 210736
rect 790 210464 69120 210728
rect 880 210456 69120 210464
rect 880 210184 69200 210456
rect 790 209920 69200 210184
rect 880 209648 69200 209920
rect 880 209640 69120 209648
rect 790 209376 69120 209640
rect 880 209368 69120 209376
rect 880 209096 69200 209368
rect 790 208832 69200 209096
rect 880 208560 69200 208832
rect 880 208552 69120 208560
rect 790 208288 69120 208552
rect 880 208280 69120 208288
rect 880 208008 69200 208280
rect 790 207744 69200 208008
rect 880 207472 69200 207744
rect 880 207464 69120 207472
rect 790 207200 69120 207464
rect 880 207192 69120 207200
rect 880 206920 69200 207192
rect 790 206656 69200 206920
rect 880 206384 69200 206656
rect 880 206376 69120 206384
rect 790 206112 69120 206376
rect 880 206104 69120 206112
rect 880 205832 69200 206104
rect 790 205568 69200 205832
rect 880 205296 69200 205568
rect 880 205288 69120 205296
rect 790 205024 69120 205288
rect 880 205016 69120 205024
rect 880 204744 69200 205016
rect 790 204480 69200 204744
rect 880 204208 69200 204480
rect 880 204200 69120 204208
rect 790 203936 69120 204200
rect 880 203928 69120 203936
rect 880 203656 69200 203928
rect 790 203392 69200 203656
rect 880 203120 69200 203392
rect 880 203112 69120 203120
rect 790 202848 69120 203112
rect 880 202840 69120 202848
rect 880 202568 69200 202840
rect 790 202304 69200 202568
rect 880 202032 69200 202304
rect 880 202024 69120 202032
rect 790 201760 69120 202024
rect 880 201752 69120 201760
rect 880 201480 69200 201752
rect 790 201216 69200 201480
rect 880 200944 69200 201216
rect 880 200936 69120 200944
rect 790 200672 69120 200936
rect 880 200664 69120 200672
rect 880 200392 69200 200664
rect 790 200128 69200 200392
rect 880 199856 69200 200128
rect 880 199848 69120 199856
rect 790 199584 69120 199848
rect 880 199576 69120 199584
rect 880 199304 69200 199576
rect 790 199040 69200 199304
rect 880 198768 69200 199040
rect 880 198760 69120 198768
rect 790 198496 69120 198760
rect 880 198488 69120 198496
rect 880 198216 69200 198488
rect 790 197952 69200 198216
rect 880 197680 69200 197952
rect 880 197672 69120 197680
rect 790 197408 69120 197672
rect 880 197400 69120 197408
rect 880 197128 69200 197400
rect 790 196864 69200 197128
rect 880 196592 69200 196864
rect 880 196584 69120 196592
rect 790 196320 69120 196584
rect 880 196312 69120 196320
rect 880 196040 69200 196312
rect 790 195776 69200 196040
rect 880 195504 69200 195776
rect 880 195496 69120 195504
rect 790 195232 69120 195496
rect 880 195224 69120 195232
rect 880 194952 69200 195224
rect 790 194688 69200 194952
rect 880 194416 69200 194688
rect 880 194408 69120 194416
rect 790 194144 69120 194408
rect 880 194136 69120 194144
rect 880 193864 69200 194136
rect 790 193600 69200 193864
rect 880 193328 69200 193600
rect 880 193320 69120 193328
rect 790 193056 69120 193320
rect 880 193048 69120 193056
rect 880 192776 69200 193048
rect 790 192512 69200 192776
rect 880 192240 69200 192512
rect 880 192232 69120 192240
rect 790 191968 69120 192232
rect 880 191960 69120 191968
rect 880 191688 69200 191960
rect 790 191424 69200 191688
rect 880 191152 69200 191424
rect 880 191144 69120 191152
rect 790 190880 69120 191144
rect 880 190872 69120 190880
rect 880 190600 69200 190872
rect 790 190336 69200 190600
rect 880 190064 69200 190336
rect 880 190056 69120 190064
rect 790 189792 69120 190056
rect 880 189784 69120 189792
rect 880 189512 69200 189784
rect 790 189248 69200 189512
rect 880 188976 69200 189248
rect 880 188968 69120 188976
rect 790 188704 69120 188968
rect 880 188696 69120 188704
rect 880 188424 69200 188696
rect 790 188160 69200 188424
rect 880 187888 69200 188160
rect 880 187880 69120 187888
rect 790 187616 69120 187880
rect 880 187608 69120 187616
rect 880 187336 69200 187608
rect 790 187072 69200 187336
rect 880 186800 69200 187072
rect 880 186792 69120 186800
rect 790 186528 69120 186792
rect 880 186520 69120 186528
rect 880 186248 69200 186520
rect 790 185984 69200 186248
rect 880 185712 69200 185984
rect 880 185704 69120 185712
rect 790 185440 69120 185704
rect 880 185432 69120 185440
rect 880 185160 69200 185432
rect 790 184896 69200 185160
rect 880 184624 69200 184896
rect 880 184616 69120 184624
rect 790 184352 69120 184616
rect 880 184344 69120 184352
rect 880 184072 69200 184344
rect 790 183808 69200 184072
rect 880 183536 69200 183808
rect 880 183528 69120 183536
rect 790 183264 69120 183528
rect 880 183256 69120 183264
rect 880 182984 69200 183256
rect 790 182720 69200 182984
rect 880 182448 69200 182720
rect 880 182440 69120 182448
rect 790 182176 69120 182440
rect 880 182168 69120 182176
rect 880 181896 69200 182168
rect 790 181632 69200 181896
rect 880 181360 69200 181632
rect 880 181352 69120 181360
rect 790 181088 69120 181352
rect 880 181080 69120 181088
rect 880 180808 69200 181080
rect 790 180544 69200 180808
rect 880 180272 69200 180544
rect 880 180264 69120 180272
rect 790 180000 69120 180264
rect 880 179992 69120 180000
rect 880 179720 69200 179992
rect 790 179456 69200 179720
rect 880 179184 69200 179456
rect 880 179176 69120 179184
rect 790 178912 69120 179176
rect 880 178904 69120 178912
rect 880 178632 69200 178904
rect 790 178368 69200 178632
rect 880 178096 69200 178368
rect 880 178088 69120 178096
rect 790 177824 69120 178088
rect 880 177816 69120 177824
rect 880 177544 69200 177816
rect 790 177280 69200 177544
rect 880 177008 69200 177280
rect 880 177000 69120 177008
rect 790 176736 69120 177000
rect 880 176728 69120 176736
rect 880 176456 69200 176728
rect 790 176192 69200 176456
rect 880 175920 69200 176192
rect 880 175912 69120 175920
rect 790 175648 69120 175912
rect 880 175640 69120 175648
rect 880 175368 69200 175640
rect 790 175104 69200 175368
rect 880 174832 69200 175104
rect 880 174824 69120 174832
rect 790 174560 69120 174824
rect 880 174552 69120 174560
rect 880 174280 69200 174552
rect 790 174016 69200 174280
rect 880 173744 69200 174016
rect 880 173736 69120 173744
rect 790 173472 69120 173736
rect 880 173464 69120 173472
rect 880 173192 69200 173464
rect 790 172928 69200 173192
rect 880 172656 69200 172928
rect 880 172648 69120 172656
rect 790 172384 69120 172648
rect 880 172376 69120 172384
rect 880 172104 69200 172376
rect 790 171840 69200 172104
rect 880 171568 69200 171840
rect 880 171560 69120 171568
rect 790 171296 69120 171560
rect 880 171288 69120 171296
rect 880 171016 69200 171288
rect 790 170752 69200 171016
rect 880 170480 69200 170752
rect 880 170472 69120 170480
rect 790 170208 69120 170472
rect 880 170200 69120 170208
rect 880 169928 69200 170200
rect 790 169664 69200 169928
rect 880 169392 69200 169664
rect 880 169384 69120 169392
rect 790 169120 69120 169384
rect 880 169112 69120 169120
rect 880 168840 69200 169112
rect 790 168576 69200 168840
rect 880 168304 69200 168576
rect 880 168296 69120 168304
rect 790 168032 69120 168296
rect 880 168024 69120 168032
rect 880 167752 69200 168024
rect 790 167488 69200 167752
rect 880 167216 69200 167488
rect 880 167208 69120 167216
rect 790 166944 69120 167208
rect 880 166936 69120 166944
rect 880 166664 69200 166936
rect 790 166400 69200 166664
rect 880 166128 69200 166400
rect 880 166120 69120 166128
rect 790 165856 69120 166120
rect 880 165848 69120 165856
rect 880 165576 69200 165848
rect 790 165312 69200 165576
rect 880 165040 69200 165312
rect 880 165032 69120 165040
rect 790 164768 69120 165032
rect 880 164760 69120 164768
rect 880 164488 69200 164760
rect 790 164224 69200 164488
rect 880 163952 69200 164224
rect 880 163944 69120 163952
rect 790 163680 69120 163944
rect 880 163672 69120 163680
rect 880 163400 69200 163672
rect 790 163136 69200 163400
rect 880 162864 69200 163136
rect 880 162856 69120 162864
rect 790 162592 69120 162856
rect 880 162584 69120 162592
rect 880 162312 69200 162584
rect 790 162048 69200 162312
rect 880 161776 69200 162048
rect 880 161768 69120 161776
rect 790 161504 69120 161768
rect 880 161496 69120 161504
rect 880 161224 69200 161496
rect 790 160960 69200 161224
rect 880 160688 69200 160960
rect 880 160680 69120 160688
rect 790 160416 69120 160680
rect 880 160408 69120 160416
rect 880 160136 69200 160408
rect 790 159872 69200 160136
rect 880 159600 69200 159872
rect 880 159592 69120 159600
rect 790 159328 69120 159592
rect 880 159320 69120 159328
rect 880 159048 69200 159320
rect 790 158784 69200 159048
rect 880 158512 69200 158784
rect 880 158504 69120 158512
rect 790 158240 69120 158504
rect 880 158232 69120 158240
rect 880 157960 69200 158232
rect 790 157696 69200 157960
rect 880 157424 69200 157696
rect 880 157416 69120 157424
rect 790 157152 69120 157416
rect 880 157144 69120 157152
rect 880 156872 69200 157144
rect 790 156608 69200 156872
rect 880 156336 69200 156608
rect 880 156328 69120 156336
rect 790 156064 69120 156328
rect 880 156056 69120 156064
rect 880 155784 69200 156056
rect 790 155520 69200 155784
rect 880 155248 69200 155520
rect 880 155240 69120 155248
rect 790 154976 69120 155240
rect 880 154968 69120 154976
rect 880 154696 69200 154968
rect 790 154432 69200 154696
rect 880 154160 69200 154432
rect 880 154152 69120 154160
rect 790 153888 69120 154152
rect 880 153880 69120 153888
rect 880 153608 69200 153880
rect 790 153344 69200 153608
rect 880 153072 69200 153344
rect 880 153064 69120 153072
rect 790 152800 69120 153064
rect 880 152792 69120 152800
rect 880 152520 69200 152792
rect 790 152256 69200 152520
rect 880 151984 69200 152256
rect 880 151976 69120 151984
rect 790 151712 69120 151976
rect 880 151704 69120 151712
rect 880 151432 69200 151704
rect 790 151168 69200 151432
rect 880 150896 69200 151168
rect 880 150888 69120 150896
rect 790 150624 69120 150888
rect 880 150616 69120 150624
rect 880 150344 69200 150616
rect 790 150080 69200 150344
rect 880 149808 69200 150080
rect 880 149800 69120 149808
rect 790 149536 69120 149800
rect 880 149528 69120 149536
rect 880 149256 69200 149528
rect 790 148992 69200 149256
rect 880 148720 69200 148992
rect 880 148712 69120 148720
rect 790 148448 69120 148712
rect 880 148440 69120 148448
rect 880 148168 69200 148440
rect 790 147904 69200 148168
rect 880 147632 69200 147904
rect 880 147624 69120 147632
rect 790 147360 69120 147624
rect 880 147352 69120 147360
rect 880 147080 69200 147352
rect 790 146816 69200 147080
rect 880 146544 69200 146816
rect 880 146536 69120 146544
rect 790 146272 69120 146536
rect 880 146264 69120 146272
rect 880 145992 69200 146264
rect 790 145728 69200 145992
rect 880 145456 69200 145728
rect 880 145448 69120 145456
rect 790 145184 69120 145448
rect 880 145176 69120 145184
rect 880 144904 69200 145176
rect 790 144640 69200 144904
rect 880 144368 69200 144640
rect 880 144360 69120 144368
rect 790 144096 69120 144360
rect 880 144088 69120 144096
rect 880 143816 69200 144088
rect 790 143552 69200 143816
rect 880 143280 69200 143552
rect 880 143272 69120 143280
rect 790 143008 69120 143272
rect 880 143000 69120 143008
rect 880 142728 69200 143000
rect 790 142464 69200 142728
rect 880 142192 69200 142464
rect 880 142184 69120 142192
rect 790 141920 69120 142184
rect 880 141912 69120 141920
rect 880 141640 69200 141912
rect 790 141376 69200 141640
rect 880 141104 69200 141376
rect 880 141096 69120 141104
rect 790 140832 69120 141096
rect 880 140824 69120 140832
rect 880 140552 69200 140824
rect 790 140288 69200 140552
rect 880 140016 69200 140288
rect 880 140008 69120 140016
rect 790 139744 69120 140008
rect 880 139736 69120 139744
rect 880 139464 69200 139736
rect 790 139200 69200 139464
rect 880 138928 69200 139200
rect 880 138920 69120 138928
rect 790 138656 69120 138920
rect 880 138648 69120 138656
rect 880 138376 69200 138648
rect 790 138112 69200 138376
rect 880 137840 69200 138112
rect 880 137832 69120 137840
rect 790 137568 69120 137832
rect 880 137560 69120 137568
rect 880 137288 69200 137560
rect 790 137024 69200 137288
rect 880 136752 69200 137024
rect 880 136744 69120 136752
rect 790 136480 69120 136744
rect 880 136472 69120 136480
rect 880 136200 69200 136472
rect 790 135936 69200 136200
rect 880 135664 69200 135936
rect 880 135656 69120 135664
rect 790 135392 69120 135656
rect 880 135384 69120 135392
rect 880 135112 69200 135384
rect 790 134848 69200 135112
rect 880 134576 69200 134848
rect 880 134568 69120 134576
rect 790 134304 69120 134568
rect 880 134296 69120 134304
rect 880 134024 69200 134296
rect 790 133760 69200 134024
rect 880 133488 69200 133760
rect 880 133480 69120 133488
rect 790 133216 69120 133480
rect 880 133208 69120 133216
rect 880 132936 69200 133208
rect 790 132672 69200 132936
rect 880 132400 69200 132672
rect 880 132392 69120 132400
rect 790 132128 69120 132392
rect 880 132120 69120 132128
rect 880 131848 69200 132120
rect 790 131584 69200 131848
rect 880 131312 69200 131584
rect 880 131304 69120 131312
rect 790 131040 69120 131304
rect 880 131032 69120 131040
rect 880 130760 69200 131032
rect 790 130496 69200 130760
rect 880 130224 69200 130496
rect 880 130216 69120 130224
rect 790 129952 69120 130216
rect 880 129944 69120 129952
rect 880 129672 69200 129944
rect 790 129408 69200 129672
rect 880 129136 69200 129408
rect 880 129128 69120 129136
rect 790 128864 69120 129128
rect 880 128856 69120 128864
rect 880 128584 69200 128856
rect 790 128320 69200 128584
rect 880 128048 69200 128320
rect 880 128040 69120 128048
rect 790 127776 69120 128040
rect 880 127768 69120 127776
rect 880 127496 69200 127768
rect 790 127232 69200 127496
rect 880 126960 69200 127232
rect 880 126952 69120 126960
rect 790 126688 69120 126952
rect 880 126680 69120 126688
rect 880 126408 69200 126680
rect 790 126144 69200 126408
rect 880 125872 69200 126144
rect 880 125864 69120 125872
rect 790 125600 69120 125864
rect 880 125592 69120 125600
rect 880 125320 69200 125592
rect 790 125056 69200 125320
rect 880 124784 69200 125056
rect 880 124776 69120 124784
rect 790 124512 69120 124776
rect 880 124504 69120 124512
rect 880 124232 69200 124504
rect 790 123968 69200 124232
rect 880 123696 69200 123968
rect 880 123688 69120 123696
rect 790 123424 69120 123688
rect 880 123416 69120 123424
rect 880 123144 69200 123416
rect 790 122880 69200 123144
rect 880 122608 69200 122880
rect 880 122600 69120 122608
rect 790 122336 69120 122600
rect 880 122328 69120 122336
rect 880 122056 69200 122328
rect 790 121792 69200 122056
rect 880 121520 69200 121792
rect 880 121512 69120 121520
rect 790 121248 69120 121512
rect 880 121240 69120 121248
rect 880 120968 69200 121240
rect 790 120704 69200 120968
rect 880 120432 69200 120704
rect 880 120424 69120 120432
rect 790 120160 69120 120424
rect 880 120152 69120 120160
rect 880 119880 69200 120152
rect 790 119616 69200 119880
rect 880 119344 69200 119616
rect 880 119336 69120 119344
rect 790 119072 69120 119336
rect 880 119064 69120 119072
rect 880 118792 69200 119064
rect 790 118528 69200 118792
rect 880 118256 69200 118528
rect 880 118248 69120 118256
rect 790 117984 69120 118248
rect 880 117976 69120 117984
rect 880 117704 69200 117976
rect 790 117440 69200 117704
rect 880 117168 69200 117440
rect 880 117160 69120 117168
rect 790 116896 69120 117160
rect 880 116888 69120 116896
rect 880 116616 69200 116888
rect 790 116352 69200 116616
rect 880 116080 69200 116352
rect 880 116072 69120 116080
rect 790 115808 69120 116072
rect 880 115800 69120 115808
rect 880 115528 69200 115800
rect 790 115264 69200 115528
rect 880 114992 69200 115264
rect 880 114984 69120 114992
rect 790 114720 69120 114984
rect 880 114712 69120 114720
rect 880 114440 69200 114712
rect 790 114176 69200 114440
rect 880 113904 69200 114176
rect 880 113896 69120 113904
rect 790 113632 69120 113896
rect 880 113624 69120 113632
rect 880 113352 69200 113624
rect 790 113088 69200 113352
rect 880 112816 69200 113088
rect 880 112808 69120 112816
rect 790 112544 69120 112808
rect 880 112536 69120 112544
rect 880 112264 69200 112536
rect 790 112000 69200 112264
rect 880 111728 69200 112000
rect 880 111720 69120 111728
rect 790 111456 69120 111720
rect 880 111448 69120 111456
rect 880 111176 69200 111448
rect 790 110912 69200 111176
rect 880 110640 69200 110912
rect 880 110632 69120 110640
rect 790 110368 69120 110632
rect 880 110360 69120 110368
rect 880 110088 69200 110360
rect 790 109824 69200 110088
rect 880 109552 69200 109824
rect 880 109544 69120 109552
rect 790 109280 69120 109544
rect 880 109272 69120 109280
rect 880 109000 69200 109272
rect 790 108736 69200 109000
rect 880 108464 69200 108736
rect 880 108456 69120 108464
rect 790 108192 69120 108456
rect 880 108184 69120 108192
rect 880 107912 69200 108184
rect 790 107648 69200 107912
rect 880 107376 69200 107648
rect 880 107368 69120 107376
rect 790 107104 69120 107368
rect 880 107096 69120 107104
rect 880 106824 69200 107096
rect 790 106560 69200 106824
rect 880 106288 69200 106560
rect 880 106280 69120 106288
rect 790 106016 69120 106280
rect 880 106008 69120 106016
rect 880 105736 69200 106008
rect 790 105472 69200 105736
rect 880 105200 69200 105472
rect 880 105192 69120 105200
rect 790 104928 69120 105192
rect 880 104920 69120 104928
rect 880 104648 69200 104920
rect 790 104384 69200 104648
rect 880 104112 69200 104384
rect 880 104104 69120 104112
rect 790 103840 69120 104104
rect 880 103832 69120 103840
rect 880 103560 69200 103832
rect 790 103296 69200 103560
rect 880 103024 69200 103296
rect 880 103016 69120 103024
rect 790 102752 69120 103016
rect 880 102744 69120 102752
rect 880 102472 69200 102744
rect 790 102208 69200 102472
rect 880 101936 69200 102208
rect 880 101928 69120 101936
rect 790 101664 69120 101928
rect 880 101656 69120 101664
rect 880 101384 69200 101656
rect 790 101120 69200 101384
rect 880 100848 69200 101120
rect 880 100840 69120 100848
rect 790 100576 69120 100840
rect 880 100568 69120 100576
rect 880 100296 69200 100568
rect 790 100032 69200 100296
rect 880 99760 69200 100032
rect 880 99752 69120 99760
rect 790 99488 69120 99752
rect 880 99480 69120 99488
rect 880 99208 69200 99480
rect 790 98944 69200 99208
rect 880 98672 69200 98944
rect 880 98664 69120 98672
rect 790 98400 69120 98664
rect 880 98392 69120 98400
rect 880 98120 69200 98392
rect 790 97856 69200 98120
rect 880 97584 69200 97856
rect 880 97576 69120 97584
rect 790 97312 69120 97576
rect 880 97304 69120 97312
rect 880 97032 69200 97304
rect 790 96768 69200 97032
rect 880 96496 69200 96768
rect 880 96488 69120 96496
rect 790 96224 69120 96488
rect 880 96216 69120 96224
rect 880 95944 69200 96216
rect 790 95680 69200 95944
rect 880 95408 69200 95680
rect 880 95400 69120 95408
rect 790 95136 69120 95400
rect 880 95128 69120 95136
rect 880 94856 69200 95128
rect 790 94592 69200 94856
rect 880 94320 69200 94592
rect 880 94312 69120 94320
rect 790 94048 69120 94312
rect 880 94040 69120 94048
rect 880 93768 69200 94040
rect 790 93504 69200 93768
rect 880 93232 69200 93504
rect 880 93224 69120 93232
rect 790 92960 69120 93224
rect 880 92952 69120 92960
rect 880 92680 69200 92952
rect 790 92416 69200 92680
rect 880 92144 69200 92416
rect 880 92136 69120 92144
rect 790 91872 69120 92136
rect 880 91864 69120 91872
rect 880 91592 69200 91864
rect 790 91328 69200 91592
rect 880 91056 69200 91328
rect 880 91048 69120 91056
rect 790 90784 69120 91048
rect 880 90776 69120 90784
rect 880 90504 69200 90776
rect 790 90240 69200 90504
rect 880 89968 69200 90240
rect 880 89960 69120 89968
rect 790 89696 69120 89960
rect 880 89688 69120 89696
rect 880 89416 69200 89688
rect 790 89152 69200 89416
rect 880 88880 69200 89152
rect 880 88872 69120 88880
rect 790 88608 69120 88872
rect 880 88600 69120 88608
rect 880 88328 69200 88600
rect 790 88064 69200 88328
rect 880 87792 69200 88064
rect 880 87784 69120 87792
rect 790 87520 69120 87784
rect 880 87512 69120 87520
rect 880 87240 69200 87512
rect 790 86976 69200 87240
rect 880 86704 69200 86976
rect 880 86696 69120 86704
rect 790 86432 69120 86696
rect 880 86424 69120 86432
rect 880 86152 69200 86424
rect 790 85888 69200 86152
rect 880 85616 69200 85888
rect 880 85608 69120 85616
rect 790 85344 69120 85608
rect 880 85336 69120 85344
rect 880 85064 69200 85336
rect 790 84800 69200 85064
rect 880 84528 69200 84800
rect 880 84520 69120 84528
rect 790 84256 69120 84520
rect 880 84248 69120 84256
rect 880 83976 69200 84248
rect 790 83712 69200 83976
rect 880 83440 69200 83712
rect 880 83432 69120 83440
rect 790 83168 69120 83432
rect 880 83160 69120 83168
rect 880 82888 69200 83160
rect 790 82624 69200 82888
rect 880 82352 69200 82624
rect 880 82344 69120 82352
rect 790 82080 69120 82344
rect 880 82072 69120 82080
rect 880 81800 69200 82072
rect 790 81536 69200 81800
rect 880 81264 69200 81536
rect 880 81256 69120 81264
rect 790 80992 69120 81256
rect 880 80984 69120 80992
rect 880 80712 69200 80984
rect 790 80448 69200 80712
rect 880 80176 69200 80448
rect 880 80168 69120 80176
rect 790 79904 69120 80168
rect 880 79896 69120 79904
rect 880 79624 69200 79896
rect 790 79360 69200 79624
rect 880 79088 69200 79360
rect 880 79080 69120 79088
rect 790 78816 69120 79080
rect 880 78808 69120 78816
rect 880 78536 69200 78808
rect 790 78272 69200 78536
rect 880 78000 69200 78272
rect 880 77992 69120 78000
rect 790 77728 69120 77992
rect 880 77720 69120 77728
rect 880 77448 69200 77720
rect 790 77184 69200 77448
rect 880 76912 69200 77184
rect 880 76904 69120 76912
rect 790 76640 69120 76904
rect 880 76632 69120 76640
rect 880 76360 69200 76632
rect 790 76096 69200 76360
rect 880 75824 69200 76096
rect 880 75816 69120 75824
rect 790 75552 69120 75816
rect 880 75544 69120 75552
rect 880 75272 69200 75544
rect 790 75008 69200 75272
rect 880 74736 69200 75008
rect 880 74728 69120 74736
rect 790 74464 69120 74728
rect 880 74456 69120 74464
rect 880 74184 69200 74456
rect 790 73920 69200 74184
rect 880 73648 69200 73920
rect 880 73640 69120 73648
rect 790 73376 69120 73640
rect 880 73368 69120 73376
rect 880 73096 69200 73368
rect 790 72832 69200 73096
rect 880 72560 69200 72832
rect 880 72552 69120 72560
rect 790 72288 69120 72552
rect 880 72280 69120 72288
rect 880 72008 69200 72280
rect 790 71744 69200 72008
rect 880 71472 69200 71744
rect 880 71464 69120 71472
rect 790 71200 69120 71464
rect 880 71192 69120 71200
rect 880 70920 69200 71192
rect 790 70656 69200 70920
rect 880 70384 69200 70656
rect 880 70376 69120 70384
rect 790 70112 69120 70376
rect 880 70104 69120 70112
rect 880 69832 69200 70104
rect 790 69568 69200 69832
rect 880 69296 69200 69568
rect 880 69288 69120 69296
rect 790 69024 69120 69288
rect 880 69016 69120 69024
rect 880 68744 69200 69016
rect 790 68480 69200 68744
rect 880 68208 69200 68480
rect 880 68200 69120 68208
rect 790 67936 69120 68200
rect 880 67928 69120 67936
rect 880 67656 69200 67928
rect 790 67392 69200 67656
rect 880 67120 69200 67392
rect 880 67112 69120 67120
rect 790 66848 69120 67112
rect 880 66840 69120 66848
rect 880 66568 69200 66840
rect 790 66304 69200 66568
rect 880 66032 69200 66304
rect 880 66024 69120 66032
rect 790 65760 69120 66024
rect 880 65752 69120 65760
rect 880 65480 69200 65752
rect 790 65216 69200 65480
rect 880 64944 69200 65216
rect 880 64936 69120 64944
rect 790 64672 69120 64936
rect 880 64664 69120 64672
rect 880 64392 69200 64664
rect 790 64128 69200 64392
rect 880 63856 69200 64128
rect 880 63848 69120 63856
rect 790 63584 69120 63848
rect 880 63576 69120 63584
rect 880 63304 69200 63576
rect 790 63040 69200 63304
rect 880 62768 69200 63040
rect 880 62760 69120 62768
rect 790 62496 69120 62760
rect 880 62488 69120 62496
rect 880 62216 69200 62488
rect 790 61952 69200 62216
rect 880 61680 69200 61952
rect 880 61672 69120 61680
rect 790 61408 69120 61672
rect 880 61400 69120 61408
rect 880 61128 69200 61400
rect 790 60864 69200 61128
rect 880 60592 69200 60864
rect 880 60584 69120 60592
rect 790 60320 69120 60584
rect 880 60312 69120 60320
rect 880 60040 69200 60312
rect 790 59776 69200 60040
rect 880 59504 69200 59776
rect 880 59496 69120 59504
rect 790 59232 69120 59496
rect 880 59224 69120 59232
rect 880 58952 69200 59224
rect 790 58688 69200 58952
rect 880 58416 69200 58688
rect 880 58408 69120 58416
rect 790 58144 69120 58408
rect 880 58136 69120 58144
rect 880 57864 69200 58136
rect 790 57600 69200 57864
rect 880 57328 69200 57600
rect 880 57320 69120 57328
rect 790 57056 69120 57320
rect 880 57048 69120 57056
rect 880 56776 69200 57048
rect 790 56512 69200 56776
rect 880 56240 69200 56512
rect 880 56232 69120 56240
rect 790 55968 69120 56232
rect 880 55960 69120 55968
rect 880 55688 69200 55960
rect 790 55424 69200 55688
rect 880 55152 69200 55424
rect 880 55144 69120 55152
rect 790 54880 69120 55144
rect 880 54872 69120 54880
rect 880 54600 69200 54872
rect 790 54336 69200 54600
rect 880 54064 69200 54336
rect 880 54056 69120 54064
rect 790 53792 69120 54056
rect 880 53784 69120 53792
rect 880 53512 69200 53784
rect 790 53248 69200 53512
rect 880 52976 69200 53248
rect 880 52968 69120 52976
rect 790 52704 69120 52968
rect 880 52696 69120 52704
rect 880 52424 69200 52696
rect 790 52160 69200 52424
rect 880 51888 69200 52160
rect 880 51880 69120 51888
rect 790 51616 69120 51880
rect 880 51608 69120 51616
rect 880 51336 69200 51608
rect 790 51072 69200 51336
rect 880 50800 69200 51072
rect 880 50792 69120 50800
rect 790 50528 69120 50792
rect 880 50520 69120 50528
rect 880 50248 69200 50520
rect 790 49984 69200 50248
rect 880 49712 69200 49984
rect 880 49704 69120 49712
rect 790 49440 69120 49704
rect 880 49432 69120 49440
rect 880 49160 69200 49432
rect 790 48896 69200 49160
rect 880 48624 69200 48896
rect 880 48616 69120 48624
rect 790 48352 69120 48616
rect 880 48344 69120 48352
rect 880 48072 69200 48344
rect 790 47808 69200 48072
rect 880 47536 69200 47808
rect 880 47528 69120 47536
rect 790 47264 69120 47528
rect 880 47256 69120 47264
rect 880 46984 69200 47256
rect 790 46720 69200 46984
rect 880 46448 69200 46720
rect 880 46440 69120 46448
rect 790 46176 69120 46440
rect 880 46168 69120 46176
rect 880 45896 69200 46168
rect 790 45632 69200 45896
rect 880 45360 69200 45632
rect 880 45352 69120 45360
rect 790 45088 69120 45352
rect 880 45080 69120 45088
rect 880 44808 69200 45080
rect 790 44544 69200 44808
rect 880 44272 69200 44544
rect 880 44264 69120 44272
rect 790 44000 69120 44264
rect 880 43992 69120 44000
rect 880 43720 69200 43992
rect 790 43456 69200 43720
rect 880 43184 69200 43456
rect 880 43176 69120 43184
rect 790 42912 69120 43176
rect 880 42904 69120 42912
rect 880 42632 69200 42904
rect 790 42368 69200 42632
rect 880 42096 69200 42368
rect 880 42088 69120 42096
rect 790 41824 69120 42088
rect 880 41816 69120 41824
rect 880 41544 69200 41816
rect 790 41280 69200 41544
rect 880 41008 69200 41280
rect 880 41000 69120 41008
rect 790 40736 69120 41000
rect 880 40728 69120 40736
rect 880 40456 69200 40728
rect 790 40192 69200 40456
rect 880 39920 69200 40192
rect 880 39912 69120 39920
rect 790 39648 69120 39912
rect 880 39640 69120 39648
rect 880 39368 69200 39640
rect 790 39104 69200 39368
rect 880 38832 69200 39104
rect 880 38824 69120 38832
rect 790 38560 69120 38824
rect 880 38552 69120 38560
rect 880 38280 69200 38552
rect 790 38016 69200 38280
rect 880 37744 69200 38016
rect 880 37736 69120 37744
rect 790 37472 69120 37736
rect 880 37464 69120 37472
rect 880 37192 69200 37464
rect 790 36928 69200 37192
rect 880 36656 69200 36928
rect 880 36648 69120 36656
rect 790 36384 69120 36648
rect 880 36376 69120 36384
rect 880 36104 69200 36376
rect 790 35840 69200 36104
rect 880 35568 69200 35840
rect 880 35560 69120 35568
rect 790 35296 69120 35560
rect 880 35288 69120 35296
rect 880 35016 69200 35288
rect 790 34752 69200 35016
rect 880 34480 69200 34752
rect 880 34472 69120 34480
rect 790 34208 69120 34472
rect 880 34200 69120 34208
rect 880 33928 69200 34200
rect 790 33664 69200 33928
rect 880 33392 69200 33664
rect 880 33384 69120 33392
rect 790 33120 69120 33384
rect 880 33112 69120 33120
rect 880 32840 69200 33112
rect 790 32576 69200 32840
rect 880 32304 69200 32576
rect 880 32296 69120 32304
rect 790 32032 69120 32296
rect 880 32024 69120 32032
rect 880 31752 69200 32024
rect 790 31488 69200 31752
rect 880 31216 69200 31488
rect 880 31208 69120 31216
rect 790 30944 69120 31208
rect 880 30936 69120 30944
rect 880 30664 69200 30936
rect 790 30400 69200 30664
rect 880 30128 69200 30400
rect 880 30120 69120 30128
rect 790 29856 69120 30120
rect 880 29848 69120 29856
rect 880 29576 69200 29848
rect 790 29312 69200 29576
rect 880 29040 69200 29312
rect 880 29032 69120 29040
rect 790 28768 69120 29032
rect 880 28760 69120 28768
rect 880 28488 69200 28760
rect 790 28224 69200 28488
rect 880 27952 69200 28224
rect 880 27944 69120 27952
rect 790 27680 69120 27944
rect 880 27672 69120 27680
rect 880 27400 69200 27672
rect 790 27136 69200 27400
rect 880 26864 69200 27136
rect 880 26856 69120 26864
rect 790 26592 69120 26856
rect 880 26584 69120 26592
rect 880 26312 69200 26584
rect 790 26048 69200 26312
rect 880 25776 69200 26048
rect 880 25768 69120 25776
rect 790 25504 69120 25768
rect 880 25496 69120 25504
rect 880 25224 69200 25496
rect 790 24960 69200 25224
rect 880 24688 69200 24960
rect 880 24680 69120 24688
rect 790 24416 69120 24680
rect 880 24408 69120 24416
rect 880 24136 69200 24408
rect 790 23872 69200 24136
rect 880 23600 69200 23872
rect 880 23592 69120 23600
rect 790 23328 69120 23592
rect 880 23320 69120 23328
rect 880 23048 69200 23320
rect 790 22784 69200 23048
rect 880 22512 69200 22784
rect 880 22504 69120 22512
rect 790 22240 69120 22504
rect 880 22232 69120 22240
rect 880 21960 69200 22232
rect 790 21696 69200 21960
rect 880 21424 69200 21696
rect 880 21416 69120 21424
rect 790 21152 69120 21416
rect 880 21144 69120 21152
rect 880 20872 69200 21144
rect 790 20608 69200 20872
rect 880 20336 69200 20608
rect 880 20328 69120 20336
rect 790 20064 69120 20328
rect 880 20056 69120 20064
rect 880 19784 69200 20056
rect 790 19520 69200 19784
rect 880 19248 69200 19520
rect 880 19240 69120 19248
rect 790 18976 69120 19240
rect 880 18968 69120 18976
rect 880 18696 69200 18968
rect 790 18432 69200 18696
rect 880 18160 69200 18432
rect 880 18152 69120 18160
rect 790 17888 69120 18152
rect 880 17880 69120 17888
rect 880 17608 69200 17880
rect 790 17344 69200 17608
rect 880 17072 69200 17344
rect 880 17064 69120 17072
rect 790 16800 69120 17064
rect 880 16792 69120 16800
rect 880 16520 69200 16792
rect 790 16256 69200 16520
rect 880 15984 69200 16256
rect 880 15976 69120 15984
rect 790 15712 69120 15976
rect 880 15704 69120 15712
rect 880 15432 69200 15704
rect 790 15168 69200 15432
rect 880 14896 69200 15168
rect 880 14888 69120 14896
rect 790 14624 69120 14888
rect 880 14616 69120 14624
rect 880 14344 69200 14616
rect 790 14080 69200 14344
rect 880 13808 69200 14080
rect 880 13800 69120 13808
rect 790 13536 69120 13800
rect 880 13528 69120 13536
rect 880 13256 69200 13528
rect 790 12992 69200 13256
rect 880 12720 69200 12992
rect 880 12712 69120 12720
rect 790 12448 69120 12712
rect 880 12440 69120 12448
rect 880 12168 69200 12440
rect 790 11904 69200 12168
rect 880 11632 69200 11904
rect 880 11624 69120 11632
rect 790 11360 69120 11624
rect 880 11352 69120 11360
rect 880 11080 69200 11352
rect 790 10816 69200 11080
rect 880 10544 69200 10816
rect 880 10536 69120 10544
rect 790 10272 69120 10536
rect 880 10264 69120 10272
rect 880 9992 69200 10264
rect 790 9728 69200 9992
rect 880 9456 69200 9728
rect 880 9448 69120 9456
rect 790 9184 69120 9448
rect 880 9176 69120 9184
rect 880 8904 69200 9176
rect 790 8640 69200 8904
rect 880 8368 69200 8640
rect 880 8360 69120 8368
rect 790 8096 69120 8360
rect 880 8088 69120 8096
rect 880 7816 69200 8088
rect 790 7552 69200 7816
rect 880 7280 69200 7552
rect 880 7272 69120 7280
rect 790 7008 69120 7272
rect 880 7000 69120 7008
rect 880 6728 69200 7000
rect 790 6464 69200 6728
rect 880 6192 69200 6464
rect 880 6184 69120 6192
rect 790 5920 69120 6184
rect 880 5912 69120 5920
rect 880 5640 69200 5912
rect 790 5376 69200 5640
rect 880 5104 69200 5376
rect 880 5096 69120 5104
rect 790 4832 69120 5096
rect 880 4824 69120 4832
rect 880 4552 69200 4824
rect 790 4288 69200 4552
rect 880 4016 69200 4288
rect 880 4008 69120 4016
rect 790 3744 69120 4008
rect 880 3736 69120 3744
rect 880 3464 69200 3736
rect 790 3200 69200 3464
rect 880 2920 69200 3200
rect 790 2656 69200 2920
rect 880 2376 69200 2656
rect 790 2112 69200 2376
rect 880 1832 69200 2112
rect 790 1568 69200 1832
rect 880 1395 69200 1568
<< metal4 >>
rect 4208 2128 4528 217648
rect 19568 2128 19888 217648
rect 34928 2128 35248 217648
rect 50288 2128 50608 217648
rect 65648 2128 65968 217648
<< obsm4 >>
rect 795 3979 4128 217429
rect 4608 3979 19488 217429
rect 19968 3979 34848 217429
rect 35328 3979 50208 217429
rect 50688 3979 64525 217429
<< labels >>
rlabel metal2 s 12070 0 12126 800 6 master0_wb_ack_i
port 1 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 master0_wb_adr_o[0]
port 2 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 master0_wb_adr_o[10]
port 3 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 master0_wb_adr_o[11]
port 4 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 master0_wb_adr_o[12]
port 5 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 master0_wb_adr_o[13]
port 6 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 master0_wb_adr_o[14]
port 7 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 master0_wb_adr_o[15]
port 8 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 master0_wb_adr_o[16]
port 9 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 master0_wb_adr_o[17]
port 10 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 master0_wb_adr_o[18]
port 11 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 master0_wb_adr_o[19]
port 12 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 master0_wb_adr_o[1]
port 13 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 master0_wb_adr_o[20]
port 14 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 master0_wb_adr_o[21]
port 15 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 master0_wb_adr_o[22]
port 16 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 master0_wb_adr_o[23]
port 17 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 master0_wb_adr_o[24]
port 18 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 master0_wb_adr_o[25]
port 19 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 master0_wb_adr_o[26]
port 20 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 master0_wb_adr_o[27]
port 21 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 master0_wb_adr_o[2]
port 22 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 master0_wb_adr_o[3]
port 23 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 master0_wb_adr_o[4]
port 24 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 master0_wb_adr_o[5]
port 25 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 master0_wb_adr_o[6]
port 26 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 master0_wb_adr_o[7]
port 27 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 master0_wb_adr_o[8]
port 28 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 master0_wb_adr_o[9]
port 29 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 master0_wb_cyc_o
port 30 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 master0_wb_data_i[0]
port 31 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 master0_wb_data_i[10]
port 32 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 master0_wb_data_i[11]
port 33 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 master0_wb_data_i[12]
port 34 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 master0_wb_data_i[13]
port 35 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 master0_wb_data_i[14]
port 36 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 master0_wb_data_i[15]
port 37 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 master0_wb_data_i[16]
port 38 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 master0_wb_data_i[17]
port 39 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 master0_wb_data_i[18]
port 40 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 master0_wb_data_i[19]
port 41 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 master0_wb_data_i[1]
port 42 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 master0_wb_data_i[20]
port 43 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 master0_wb_data_i[21]
port 44 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 master0_wb_data_i[22]
port 45 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 master0_wb_data_i[23]
port 46 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 master0_wb_data_i[24]
port 47 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 master0_wb_data_i[25]
port 48 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 master0_wb_data_i[26]
port 49 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 master0_wb_data_i[27]
port 50 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 master0_wb_data_i[28]
port 51 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 master0_wb_data_i[29]
port 52 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 master0_wb_data_i[2]
port 53 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 master0_wb_data_i[30]
port 54 nsew signal output
rlabel metal2 s 67270 0 67326 800 6 master0_wb_data_i[31]
port 55 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 master0_wb_data_i[3]
port 56 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 master0_wb_data_i[4]
port 57 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 master0_wb_data_i[5]
port 58 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 master0_wb_data_i[6]
port 59 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 master0_wb_data_i[7]
port 60 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 master0_wb_data_i[8]
port 61 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 master0_wb_data_i[9]
port 62 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 master0_wb_data_o[0]
port 63 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 master0_wb_data_o[10]
port 64 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 master0_wb_data_o[11]
port 65 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 master0_wb_data_o[12]
port 66 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 master0_wb_data_o[13]
port 67 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 master0_wb_data_o[14]
port 68 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 master0_wb_data_o[15]
port 69 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 master0_wb_data_o[16]
port 70 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 master0_wb_data_o[17]
port 71 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 master0_wb_data_o[18]
port 72 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 master0_wb_data_o[19]
port 73 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 master0_wb_data_o[1]
port 74 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 master0_wb_data_o[20]
port 75 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 master0_wb_data_o[21]
port 76 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 master0_wb_data_o[22]
port 77 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 master0_wb_data_o[23]
port 78 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 master0_wb_data_o[24]
port 79 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 master0_wb_data_o[25]
port 80 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 master0_wb_data_o[26]
port 81 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 master0_wb_data_o[27]
port 82 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 master0_wb_data_o[28]
port 83 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 master0_wb_data_o[29]
port 84 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 master0_wb_data_o[2]
port 85 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 master0_wb_data_o[30]
port 86 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 master0_wb_data_o[31]
port 87 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 master0_wb_data_o[3]
port 88 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 master0_wb_data_o[4]
port 89 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 master0_wb_data_o[5]
port 90 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 master0_wb_data_o[6]
port 91 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 master0_wb_data_o[7]
port 92 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 master0_wb_data_o[8]
port 93 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 master0_wb_data_o[9]
port 94 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 master0_wb_error_i
port 95 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 master0_wb_sel_o[0]
port 96 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 master0_wb_sel_o[1]
port 97 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 master0_wb_sel_o[2]
port 98 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 master0_wb_sel_o[3]
port 99 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 master0_wb_stall_i
port 100 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 master0_wb_stb_o
port 101 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 master0_wb_we_o
port 102 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 master1_wb_ack_i
port 103 nsew signal output
rlabel metal3 s 0 113432 800 113552 6 master1_wb_adr_o[0]
port 104 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 master1_wb_adr_o[10]
port 105 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 master1_wb_adr_o[11]
port 106 nsew signal input
rlabel metal3 s 0 135192 800 135312 6 master1_wb_adr_o[12]
port 107 nsew signal input
rlabel metal3 s 0 136824 800 136944 6 master1_wb_adr_o[13]
port 108 nsew signal input
rlabel metal3 s 0 138456 800 138576 6 master1_wb_adr_o[14]
port 109 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 master1_wb_adr_o[15]
port 110 nsew signal input
rlabel metal3 s 0 141720 800 141840 6 master1_wb_adr_o[16]
port 111 nsew signal input
rlabel metal3 s 0 143352 800 143472 6 master1_wb_adr_o[17]
port 112 nsew signal input
rlabel metal3 s 0 144984 800 145104 6 master1_wb_adr_o[18]
port 113 nsew signal input
rlabel metal3 s 0 146616 800 146736 6 master1_wb_adr_o[19]
port 114 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 master1_wb_adr_o[1]
port 115 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 master1_wb_adr_o[20]
port 116 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 master1_wb_adr_o[21]
port 117 nsew signal input
rlabel metal3 s 0 151512 800 151632 6 master1_wb_adr_o[22]
port 118 nsew signal input
rlabel metal3 s 0 153144 800 153264 6 master1_wb_adr_o[23]
port 119 nsew signal input
rlabel metal3 s 0 154776 800 154896 6 master1_wb_adr_o[24]
port 120 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 master1_wb_adr_o[25]
port 121 nsew signal input
rlabel metal3 s 0 158040 800 158160 6 master1_wb_adr_o[26]
port 122 nsew signal input
rlabel metal3 s 0 159672 800 159792 6 master1_wb_adr_o[27]
port 123 nsew signal input
rlabel metal3 s 0 117784 800 117904 6 master1_wb_adr_o[2]
port 124 nsew signal input
rlabel metal3 s 0 119960 800 120080 6 master1_wb_adr_o[3]
port 125 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 master1_wb_adr_o[4]
port 126 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 master1_wb_adr_o[5]
port 127 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 master1_wb_adr_o[6]
port 128 nsew signal input
rlabel metal3 s 0 127032 800 127152 6 master1_wb_adr_o[7]
port 129 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 master1_wb_adr_o[8]
port 130 nsew signal input
rlabel metal3 s 0 130296 800 130416 6 master1_wb_adr_o[9]
port 131 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 master1_wb_cyc_o
port 132 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 master1_wb_data_i[0]
port 133 nsew signal output
rlabel metal3 s 0 132472 800 132592 6 master1_wb_data_i[10]
port 134 nsew signal output
rlabel metal3 s 0 134104 800 134224 6 master1_wb_data_i[11]
port 135 nsew signal output
rlabel metal3 s 0 135736 800 135856 6 master1_wb_data_i[12]
port 136 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 master1_wb_data_i[13]
port 137 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 master1_wb_data_i[14]
port 138 nsew signal output
rlabel metal3 s 0 140632 800 140752 6 master1_wb_data_i[15]
port 139 nsew signal output
rlabel metal3 s 0 142264 800 142384 6 master1_wb_data_i[16]
port 140 nsew signal output
rlabel metal3 s 0 143896 800 144016 6 master1_wb_data_i[17]
port 141 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 master1_wb_data_i[18]
port 142 nsew signal output
rlabel metal3 s 0 147160 800 147280 6 master1_wb_data_i[19]
port 143 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 master1_wb_data_i[1]
port 144 nsew signal output
rlabel metal3 s 0 148792 800 148912 6 master1_wb_data_i[20]
port 145 nsew signal output
rlabel metal3 s 0 150424 800 150544 6 master1_wb_data_i[21]
port 146 nsew signal output
rlabel metal3 s 0 152056 800 152176 6 master1_wb_data_i[22]
port 147 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 master1_wb_data_i[23]
port 148 nsew signal output
rlabel metal3 s 0 155320 800 155440 6 master1_wb_data_i[24]
port 149 nsew signal output
rlabel metal3 s 0 156952 800 157072 6 master1_wb_data_i[25]
port 150 nsew signal output
rlabel metal3 s 0 158584 800 158704 6 master1_wb_data_i[26]
port 151 nsew signal output
rlabel metal3 s 0 160216 800 160336 6 master1_wb_data_i[27]
port 152 nsew signal output
rlabel metal3 s 0 161304 800 161424 6 master1_wb_data_i[28]
port 153 nsew signal output
rlabel metal3 s 0 162392 800 162512 6 master1_wb_data_i[29]
port 154 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 master1_wb_data_i[2]
port 155 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 master1_wb_data_i[30]
port 156 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 master1_wb_data_i[31]
port 157 nsew signal output
rlabel metal3 s 0 120504 800 120624 6 master1_wb_data_i[3]
port 158 nsew signal output
rlabel metal3 s 0 122680 800 122800 6 master1_wb_data_i[4]
port 159 nsew signal output
rlabel metal3 s 0 124312 800 124432 6 master1_wb_data_i[5]
port 160 nsew signal output
rlabel metal3 s 0 125944 800 126064 6 master1_wb_data_i[6]
port 161 nsew signal output
rlabel metal3 s 0 127576 800 127696 6 master1_wb_data_i[7]
port 162 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 master1_wb_data_i[8]
port 163 nsew signal output
rlabel metal3 s 0 130840 800 130960 6 master1_wb_data_i[9]
port 164 nsew signal output
rlabel metal3 s 0 114520 800 114640 6 master1_wb_data_o[0]
port 165 nsew signal input
rlabel metal3 s 0 133016 800 133136 6 master1_wb_data_o[10]
port 166 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 master1_wb_data_o[11]
port 167 nsew signal input
rlabel metal3 s 0 136280 800 136400 6 master1_wb_data_o[12]
port 168 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 master1_wb_data_o[13]
port 169 nsew signal input
rlabel metal3 s 0 139544 800 139664 6 master1_wb_data_o[14]
port 170 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 master1_wb_data_o[15]
port 171 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 master1_wb_data_o[16]
port 172 nsew signal input
rlabel metal3 s 0 144440 800 144560 6 master1_wb_data_o[17]
port 173 nsew signal input
rlabel metal3 s 0 146072 800 146192 6 master1_wb_data_o[18]
port 174 nsew signal input
rlabel metal3 s 0 147704 800 147824 6 master1_wb_data_o[19]
port 175 nsew signal input
rlabel metal3 s 0 116696 800 116816 6 master1_wb_data_o[1]
port 176 nsew signal input
rlabel metal3 s 0 149336 800 149456 6 master1_wb_data_o[20]
port 177 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 master1_wb_data_o[21]
port 178 nsew signal input
rlabel metal3 s 0 152600 800 152720 6 master1_wb_data_o[22]
port 179 nsew signal input
rlabel metal3 s 0 154232 800 154352 6 master1_wb_data_o[23]
port 180 nsew signal input
rlabel metal3 s 0 155864 800 155984 6 master1_wb_data_o[24]
port 181 nsew signal input
rlabel metal3 s 0 157496 800 157616 6 master1_wb_data_o[25]
port 182 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 master1_wb_data_o[26]
port 183 nsew signal input
rlabel metal3 s 0 160760 800 160880 6 master1_wb_data_o[27]
port 184 nsew signal input
rlabel metal3 s 0 161848 800 161968 6 master1_wb_data_o[28]
port 185 nsew signal input
rlabel metal3 s 0 162936 800 163056 6 master1_wb_data_o[29]
port 186 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 master1_wb_data_o[2]
port 187 nsew signal input
rlabel metal3 s 0 164024 800 164144 6 master1_wb_data_o[30]
port 188 nsew signal input
rlabel metal3 s 0 165112 800 165232 6 master1_wb_data_o[31]
port 189 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 master1_wb_data_o[3]
port 190 nsew signal input
rlabel metal3 s 0 123224 800 123344 6 master1_wb_data_o[4]
port 191 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 master1_wb_data_o[5]
port 192 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 master1_wb_data_o[6]
port 193 nsew signal input
rlabel metal3 s 0 128120 800 128240 6 master1_wb_data_o[7]
port 194 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 master1_wb_data_o[8]
port 195 nsew signal input
rlabel metal3 s 0 131384 800 131504 6 master1_wb_data_o[9]
port 196 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 master1_wb_error_i
port 197 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 master1_wb_sel_o[0]
port 198 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 master1_wb_sel_o[1]
port 199 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 master1_wb_sel_o[2]
port 200 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 master1_wb_sel_o[3]
port 201 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 master1_wb_stall_i
port 202 nsew signal output
rlabel metal3 s 0 112344 800 112464 6 master1_wb_stb_o
port 203 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 master1_wb_we_o
port 204 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 master2_wb_ack_i
port 205 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 master2_wb_adr_o[0]
port 206 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 master2_wb_adr_o[10]
port 207 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 master2_wb_adr_o[11]
port 208 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 master2_wb_adr_o[12]
port 209 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 master2_wb_adr_o[13]
port 210 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 master2_wb_adr_o[14]
port 211 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 master2_wb_adr_o[15]
port 212 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 master2_wb_adr_o[16]
port 213 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 master2_wb_adr_o[17]
port 214 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 master2_wb_adr_o[18]
port 215 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 master2_wb_adr_o[19]
port 216 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 master2_wb_adr_o[1]
port 217 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 master2_wb_adr_o[20]
port 218 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 master2_wb_adr_o[21]
port 219 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 master2_wb_adr_o[22]
port 220 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 master2_wb_adr_o[23]
port 221 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 master2_wb_adr_o[24]
port 222 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 master2_wb_adr_o[25]
port 223 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 master2_wb_adr_o[26]
port 224 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 master2_wb_adr_o[27]
port 225 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 master2_wb_adr_o[2]
port 226 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 master2_wb_adr_o[3]
port 227 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 master2_wb_adr_o[4]
port 228 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 master2_wb_adr_o[5]
port 229 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 master2_wb_adr_o[6]
port 230 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 master2_wb_adr_o[7]
port 231 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 master2_wb_adr_o[8]
port 232 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 master2_wb_adr_o[9]
port 233 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 master2_wb_cyc_o
port 234 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 master2_wb_data_i[0]
port 235 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 master2_wb_data_i[10]
port 236 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 master2_wb_data_i[11]
port 237 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 master2_wb_data_i[12]
port 238 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 master2_wb_data_i[13]
port 239 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 master2_wb_data_i[14]
port 240 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 master2_wb_data_i[15]
port 241 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 master2_wb_data_i[16]
port 242 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 master2_wb_data_i[17]
port 243 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 master2_wb_data_i[18]
port 244 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 master2_wb_data_i[19]
port 245 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 master2_wb_data_i[1]
port 246 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 master2_wb_data_i[20]
port 247 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 master2_wb_data_i[21]
port 248 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 master2_wb_data_i[22]
port 249 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 master2_wb_data_i[23]
port 250 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 master2_wb_data_i[24]
port 251 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 master2_wb_data_i[25]
port 252 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 master2_wb_data_i[26]
port 253 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 master2_wb_data_i[27]
port 254 nsew signal output
rlabel metal3 s 0 52504 800 52624 6 master2_wb_data_i[28]
port 255 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 master2_wb_data_i[29]
port 256 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 master2_wb_data_i[2]
port 257 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 master2_wb_data_i[30]
port 258 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 master2_wb_data_i[31]
port 259 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 master2_wb_data_i[3]
port 260 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 master2_wb_data_i[4]
port 261 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 master2_wb_data_i[5]
port 262 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 master2_wb_data_i[6]
port 263 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 master2_wb_data_i[7]
port 264 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 master2_wb_data_i[8]
port 265 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 master2_wb_data_i[9]
port 266 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 master2_wb_data_o[0]
port 267 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 master2_wb_data_o[10]
port 268 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 master2_wb_data_o[11]
port 269 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 master2_wb_data_o[12]
port 270 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 master2_wb_data_o[13]
port 271 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 master2_wb_data_o[14]
port 272 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 master2_wb_data_o[15]
port 273 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 master2_wb_data_o[16]
port 274 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 master2_wb_data_o[17]
port 275 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 master2_wb_data_o[18]
port 276 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 master2_wb_data_o[19]
port 277 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 master2_wb_data_o[1]
port 278 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 master2_wb_data_o[20]
port 279 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 master2_wb_data_o[21]
port 280 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 master2_wb_data_o[22]
port 281 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 master2_wb_data_o[23]
port 282 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 master2_wb_data_o[24]
port 283 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 master2_wb_data_o[25]
port 284 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 master2_wb_data_o[26]
port 285 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 master2_wb_data_o[27]
port 286 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 master2_wb_data_o[28]
port 287 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 master2_wb_data_o[29]
port 288 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 master2_wb_data_o[2]
port 289 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 master2_wb_data_o[30]
port 290 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 master2_wb_data_o[31]
port 291 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 master2_wb_data_o[3]
port 292 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 master2_wb_data_o[4]
port 293 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 master2_wb_data_o[5]
port 294 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 master2_wb_data_o[6]
port 295 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 master2_wb_data_o[7]
port 296 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 master2_wb_data_o[8]
port 297 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 master2_wb_data_o[9]
port 298 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 master2_wb_error_i
port 299 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 master2_wb_sel_o[0]
port 300 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 master2_wb_sel_o[1]
port 301 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 master2_wb_sel_o[2]
port 302 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 master2_wb_sel_o[3]
port 303 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 master2_wb_stall_i
port 304 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 master2_wb_stb_o
port 305 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 master2_wb_we_o
port 306 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 probe_master0_currentSlave[0]
port 307 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 probe_master0_currentSlave[1]
port 308 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 probe_master1_currentSlave[0]
port 309 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 probe_master1_currentSlave[1]
port 310 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 probe_master2_currentSlave[0]
port 311 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 probe_master2_currentSlave[1]
port 312 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 probe_master3_currentSlave[0]
port 313 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 probe_master3_currentSlave[1]
port 314 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 probe_slave0_currentMaster[0]
port 315 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 probe_slave0_currentMaster[1]
port 316 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 probe_slave1_currentMaster[0]
port 317 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 probe_slave1_currentMaster[1]
port 318 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 probe_slave2_currentMaster[0]
port 319 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 probe_slave2_currentMaster[1]
port 320 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 probe_slave3_currentMaster[0]
port 321 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 probe_slave3_currentMaster[1]
port 322 nsew signal output
rlabel metal3 s 0 165656 800 165776 6 slave0_wb_ack_o
port 323 nsew signal input
rlabel metal3 s 0 168920 800 169040 6 slave0_wb_adr_i[0]
port 324 nsew signal output
rlabel metal3 s 0 187416 800 187536 6 slave0_wb_adr_i[10]
port 325 nsew signal output
rlabel metal3 s 0 189048 800 189168 6 slave0_wb_adr_i[11]
port 326 nsew signal output
rlabel metal3 s 0 190680 800 190800 6 slave0_wb_adr_i[12]
port 327 nsew signal output
rlabel metal3 s 0 192312 800 192432 6 slave0_wb_adr_i[13]
port 328 nsew signal output
rlabel metal3 s 0 193944 800 194064 6 slave0_wb_adr_i[14]
port 329 nsew signal output
rlabel metal3 s 0 195576 800 195696 6 slave0_wb_adr_i[15]
port 330 nsew signal output
rlabel metal3 s 0 197208 800 197328 6 slave0_wb_adr_i[16]
port 331 nsew signal output
rlabel metal3 s 0 198840 800 198960 6 slave0_wb_adr_i[17]
port 332 nsew signal output
rlabel metal3 s 0 200472 800 200592 6 slave0_wb_adr_i[18]
port 333 nsew signal output
rlabel metal3 s 0 202104 800 202224 6 slave0_wb_adr_i[19]
port 334 nsew signal output
rlabel metal3 s 0 171096 800 171216 6 slave0_wb_adr_i[1]
port 335 nsew signal output
rlabel metal3 s 0 203736 800 203856 6 slave0_wb_adr_i[20]
port 336 nsew signal output
rlabel metal3 s 0 205368 800 205488 6 slave0_wb_adr_i[21]
port 337 nsew signal output
rlabel metal3 s 0 207000 800 207120 6 slave0_wb_adr_i[22]
port 338 nsew signal output
rlabel metal3 s 0 208632 800 208752 6 slave0_wb_adr_i[23]
port 339 nsew signal output
rlabel metal3 s 0 173272 800 173392 6 slave0_wb_adr_i[2]
port 340 nsew signal output
rlabel metal3 s 0 175448 800 175568 6 slave0_wb_adr_i[3]
port 341 nsew signal output
rlabel metal3 s 0 177624 800 177744 6 slave0_wb_adr_i[4]
port 342 nsew signal output
rlabel metal3 s 0 179256 800 179376 6 slave0_wb_adr_i[5]
port 343 nsew signal output
rlabel metal3 s 0 180888 800 181008 6 slave0_wb_adr_i[6]
port 344 nsew signal output
rlabel metal3 s 0 182520 800 182640 6 slave0_wb_adr_i[7]
port 345 nsew signal output
rlabel metal3 s 0 184152 800 184272 6 slave0_wb_adr_i[8]
port 346 nsew signal output
rlabel metal3 s 0 185784 800 185904 6 slave0_wb_adr_i[9]
port 347 nsew signal output
rlabel metal3 s 0 166200 800 166320 6 slave0_wb_cyc_i
port 348 nsew signal output
rlabel metal3 s 0 169464 800 169584 6 slave0_wb_data_i[0]
port 349 nsew signal output
rlabel metal3 s 0 187960 800 188080 6 slave0_wb_data_i[10]
port 350 nsew signal output
rlabel metal3 s 0 189592 800 189712 6 slave0_wb_data_i[11]
port 351 nsew signal output
rlabel metal3 s 0 191224 800 191344 6 slave0_wb_data_i[12]
port 352 nsew signal output
rlabel metal3 s 0 192856 800 192976 6 slave0_wb_data_i[13]
port 353 nsew signal output
rlabel metal3 s 0 194488 800 194608 6 slave0_wb_data_i[14]
port 354 nsew signal output
rlabel metal3 s 0 196120 800 196240 6 slave0_wb_data_i[15]
port 355 nsew signal output
rlabel metal3 s 0 197752 800 197872 6 slave0_wb_data_i[16]
port 356 nsew signal output
rlabel metal3 s 0 199384 800 199504 6 slave0_wb_data_i[17]
port 357 nsew signal output
rlabel metal3 s 0 201016 800 201136 6 slave0_wb_data_i[18]
port 358 nsew signal output
rlabel metal3 s 0 202648 800 202768 6 slave0_wb_data_i[19]
port 359 nsew signal output
rlabel metal3 s 0 171640 800 171760 6 slave0_wb_data_i[1]
port 360 nsew signal output
rlabel metal3 s 0 204280 800 204400 6 slave0_wb_data_i[20]
port 361 nsew signal output
rlabel metal3 s 0 205912 800 206032 6 slave0_wb_data_i[21]
port 362 nsew signal output
rlabel metal3 s 0 207544 800 207664 6 slave0_wb_data_i[22]
port 363 nsew signal output
rlabel metal3 s 0 209176 800 209296 6 slave0_wb_data_i[23]
port 364 nsew signal output
rlabel metal3 s 0 210264 800 210384 6 slave0_wb_data_i[24]
port 365 nsew signal output
rlabel metal3 s 0 211352 800 211472 6 slave0_wb_data_i[25]
port 366 nsew signal output
rlabel metal3 s 0 212440 800 212560 6 slave0_wb_data_i[26]
port 367 nsew signal output
rlabel metal3 s 0 213528 800 213648 6 slave0_wb_data_i[27]
port 368 nsew signal output
rlabel metal3 s 0 214616 800 214736 6 slave0_wb_data_i[28]
port 369 nsew signal output
rlabel metal3 s 0 215704 800 215824 6 slave0_wb_data_i[29]
port 370 nsew signal output
rlabel metal3 s 0 173816 800 173936 6 slave0_wb_data_i[2]
port 371 nsew signal output
rlabel metal3 s 0 216792 800 216912 6 slave0_wb_data_i[30]
port 372 nsew signal output
rlabel metal3 s 0 217880 800 218000 6 slave0_wb_data_i[31]
port 373 nsew signal output
rlabel metal3 s 0 175992 800 176112 6 slave0_wb_data_i[3]
port 374 nsew signal output
rlabel metal3 s 0 178168 800 178288 6 slave0_wb_data_i[4]
port 375 nsew signal output
rlabel metal3 s 0 179800 800 179920 6 slave0_wb_data_i[5]
port 376 nsew signal output
rlabel metal3 s 0 181432 800 181552 6 slave0_wb_data_i[6]
port 377 nsew signal output
rlabel metal3 s 0 183064 800 183184 6 slave0_wb_data_i[7]
port 378 nsew signal output
rlabel metal3 s 0 184696 800 184816 6 slave0_wb_data_i[8]
port 379 nsew signal output
rlabel metal3 s 0 186328 800 186448 6 slave0_wb_data_i[9]
port 380 nsew signal output
rlabel metal3 s 0 170008 800 170128 6 slave0_wb_data_o[0]
port 381 nsew signal input
rlabel metal3 s 0 188504 800 188624 6 slave0_wb_data_o[10]
port 382 nsew signal input
rlabel metal3 s 0 190136 800 190256 6 slave0_wb_data_o[11]
port 383 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 slave0_wb_data_o[12]
port 384 nsew signal input
rlabel metal3 s 0 193400 800 193520 6 slave0_wb_data_o[13]
port 385 nsew signal input
rlabel metal3 s 0 195032 800 195152 6 slave0_wb_data_o[14]
port 386 nsew signal input
rlabel metal3 s 0 196664 800 196784 6 slave0_wb_data_o[15]
port 387 nsew signal input
rlabel metal3 s 0 198296 800 198416 6 slave0_wb_data_o[16]
port 388 nsew signal input
rlabel metal3 s 0 199928 800 200048 6 slave0_wb_data_o[17]
port 389 nsew signal input
rlabel metal3 s 0 201560 800 201680 6 slave0_wb_data_o[18]
port 390 nsew signal input
rlabel metal3 s 0 203192 800 203312 6 slave0_wb_data_o[19]
port 391 nsew signal input
rlabel metal3 s 0 172184 800 172304 6 slave0_wb_data_o[1]
port 392 nsew signal input
rlabel metal3 s 0 204824 800 204944 6 slave0_wb_data_o[20]
port 393 nsew signal input
rlabel metal3 s 0 206456 800 206576 6 slave0_wb_data_o[21]
port 394 nsew signal input
rlabel metal3 s 0 208088 800 208208 6 slave0_wb_data_o[22]
port 395 nsew signal input
rlabel metal3 s 0 209720 800 209840 6 slave0_wb_data_o[23]
port 396 nsew signal input
rlabel metal3 s 0 210808 800 210928 6 slave0_wb_data_o[24]
port 397 nsew signal input
rlabel metal3 s 0 211896 800 212016 6 slave0_wb_data_o[25]
port 398 nsew signal input
rlabel metal3 s 0 212984 800 213104 6 slave0_wb_data_o[26]
port 399 nsew signal input
rlabel metal3 s 0 214072 800 214192 6 slave0_wb_data_o[27]
port 400 nsew signal input
rlabel metal3 s 0 215160 800 215280 6 slave0_wb_data_o[28]
port 401 nsew signal input
rlabel metal3 s 0 216248 800 216368 6 slave0_wb_data_o[29]
port 402 nsew signal input
rlabel metal3 s 0 174360 800 174480 6 slave0_wb_data_o[2]
port 403 nsew signal input
rlabel metal3 s 0 217336 800 217456 6 slave0_wb_data_o[30]
port 404 nsew signal input
rlabel metal3 s 0 218424 800 218544 6 slave0_wb_data_o[31]
port 405 nsew signal input
rlabel metal3 s 0 176536 800 176656 6 slave0_wb_data_o[3]
port 406 nsew signal input
rlabel metal3 s 0 178712 800 178832 6 slave0_wb_data_o[4]
port 407 nsew signal input
rlabel metal3 s 0 180344 800 180464 6 slave0_wb_data_o[5]
port 408 nsew signal input
rlabel metal3 s 0 181976 800 182096 6 slave0_wb_data_o[6]
port 409 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 slave0_wb_data_o[7]
port 410 nsew signal input
rlabel metal3 s 0 185240 800 185360 6 slave0_wb_data_o[8]
port 411 nsew signal input
rlabel metal3 s 0 186872 800 186992 6 slave0_wb_data_o[9]
port 412 nsew signal input
rlabel metal3 s 0 166744 800 166864 6 slave0_wb_error_o
port 413 nsew signal input
rlabel metal3 s 0 170552 800 170672 6 slave0_wb_sel_i[0]
port 414 nsew signal output
rlabel metal3 s 0 172728 800 172848 6 slave0_wb_sel_i[1]
port 415 nsew signal output
rlabel metal3 s 0 174904 800 175024 6 slave0_wb_sel_i[2]
port 416 nsew signal output
rlabel metal3 s 0 177080 800 177200 6 slave0_wb_sel_i[3]
port 417 nsew signal output
rlabel metal3 s 0 167288 800 167408 6 slave0_wb_stall_o
port 418 nsew signal input
rlabel metal3 s 0 167832 800 167952 6 slave0_wb_stb_i
port 419 nsew signal output
rlabel metal3 s 0 168376 800 168496 6 slave0_wb_we_i
port 420 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 slave1_wb_ack_o
port 421 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 slave1_wb_adr_i[0]
port 422 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 slave1_wb_adr_i[10]
port 423 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 slave1_wb_adr_i[11]
port 424 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 slave1_wb_adr_i[12]
port 425 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 slave1_wb_adr_i[13]
port 426 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 slave1_wb_adr_i[14]
port 427 nsew signal output
rlabel metal3 s 0 86776 800 86896 6 slave1_wb_adr_i[15]
port 428 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 slave1_wb_adr_i[16]
port 429 nsew signal output
rlabel metal3 s 0 90040 800 90160 6 slave1_wb_adr_i[17]
port 430 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 slave1_wb_adr_i[18]
port 431 nsew signal output
rlabel metal3 s 0 93304 800 93424 6 slave1_wb_adr_i[19]
port 432 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 slave1_wb_adr_i[1]
port 433 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 slave1_wb_adr_i[20]
port 434 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 slave1_wb_adr_i[21]
port 435 nsew signal output
rlabel metal3 s 0 98200 800 98320 6 slave1_wb_adr_i[22]
port 436 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 slave1_wb_adr_i[23]
port 437 nsew signal output
rlabel metal3 s 0 64472 800 64592 6 slave1_wb_adr_i[2]
port 438 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 slave1_wb_adr_i[3]
port 439 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 slave1_wb_adr_i[4]
port 440 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 slave1_wb_adr_i[5]
port 441 nsew signal output
rlabel metal3 s 0 72088 800 72208 6 slave1_wb_adr_i[6]
port 442 nsew signal output
rlabel metal3 s 0 73720 800 73840 6 slave1_wb_adr_i[7]
port 443 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 slave1_wb_adr_i[8]
port 444 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 slave1_wb_adr_i[9]
port 445 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 slave1_wb_cyc_i
port 446 nsew signal output
rlabel metal3 s 0 60664 800 60784 6 slave1_wb_data_i[0]
port 447 nsew signal output
rlabel metal3 s 0 79160 800 79280 6 slave1_wb_data_i[10]
port 448 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 slave1_wb_data_i[11]
port 449 nsew signal output
rlabel metal3 s 0 82424 800 82544 6 slave1_wb_data_i[12]
port 450 nsew signal output
rlabel metal3 s 0 84056 800 84176 6 slave1_wb_data_i[13]
port 451 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 slave1_wb_data_i[14]
port 452 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 slave1_wb_data_i[15]
port 453 nsew signal output
rlabel metal3 s 0 88952 800 89072 6 slave1_wb_data_i[16]
port 454 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 slave1_wb_data_i[17]
port 455 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 slave1_wb_data_i[18]
port 456 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 slave1_wb_data_i[19]
port 457 nsew signal output
rlabel metal3 s 0 62840 800 62960 6 slave1_wb_data_i[1]
port 458 nsew signal output
rlabel metal3 s 0 95480 800 95600 6 slave1_wb_data_i[20]
port 459 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 slave1_wb_data_i[21]
port 460 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 slave1_wb_data_i[22]
port 461 nsew signal output
rlabel metal3 s 0 100376 800 100496 6 slave1_wb_data_i[23]
port 462 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 slave1_wb_data_i[24]
port 463 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 slave1_wb_data_i[25]
port 464 nsew signal output
rlabel metal3 s 0 103640 800 103760 6 slave1_wb_data_i[26]
port 465 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 slave1_wb_data_i[27]
port 466 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 slave1_wb_data_i[28]
port 467 nsew signal output
rlabel metal3 s 0 106904 800 107024 6 slave1_wb_data_i[29]
port 468 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 slave1_wb_data_i[2]
port 469 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 slave1_wb_data_i[30]
port 470 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 slave1_wb_data_i[31]
port 471 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 slave1_wb_data_i[3]
port 472 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 slave1_wb_data_i[4]
port 473 nsew signal output
rlabel metal3 s 0 71000 800 71120 6 slave1_wb_data_i[5]
port 474 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 slave1_wb_data_i[6]
port 475 nsew signal output
rlabel metal3 s 0 74264 800 74384 6 slave1_wb_data_i[7]
port 476 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 slave1_wb_data_i[8]
port 477 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 slave1_wb_data_i[9]
port 478 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 slave1_wb_data_o[0]
port 479 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 slave1_wb_data_o[10]
port 480 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 slave1_wb_data_o[11]
port 481 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 slave1_wb_data_o[12]
port 482 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 slave1_wb_data_o[13]
port 483 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 slave1_wb_data_o[14]
port 484 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 slave1_wb_data_o[15]
port 485 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 slave1_wb_data_o[16]
port 486 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 slave1_wb_data_o[17]
port 487 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 slave1_wb_data_o[18]
port 488 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 slave1_wb_data_o[19]
port 489 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 slave1_wb_data_o[1]
port 490 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 slave1_wb_data_o[20]
port 491 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 slave1_wb_data_o[21]
port 492 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 slave1_wb_data_o[22]
port 493 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 slave1_wb_data_o[23]
port 494 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 slave1_wb_data_o[24]
port 495 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 slave1_wb_data_o[25]
port 496 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 slave1_wb_data_o[26]
port 497 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 slave1_wb_data_o[27]
port 498 nsew signal input
rlabel metal3 s 0 106360 800 106480 6 slave1_wb_data_o[28]
port 499 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 slave1_wb_data_o[29]
port 500 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 slave1_wb_data_o[2]
port 501 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 slave1_wb_data_o[30]
port 502 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 slave1_wb_data_o[31]
port 503 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 slave1_wb_data_o[3]
port 504 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 slave1_wb_data_o[4]
port 505 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 slave1_wb_data_o[5]
port 506 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 slave1_wb_data_o[6]
port 507 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 slave1_wb_data_o[7]
port 508 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 slave1_wb_data_o[8]
port 509 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 slave1_wb_data_o[9]
port 510 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 slave1_wb_error_o
port 511 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 slave1_wb_sel_i[0]
port 512 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 slave1_wb_sel_i[1]
port 513 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 slave1_wb_sel_i[2]
port 514 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 slave1_wb_sel_i[3]
port 515 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 slave1_wb_stall_o
port 516 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 slave1_wb_stb_i
port 517 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 slave1_wb_we_i
port 518 nsew signal output
rlabel metal2 s 3698 219200 3754 220000 6 slave2_wb_ack_o
port 519 nsew signal input
rlabel metal2 s 7562 219200 7618 220000 6 slave2_wb_adr_i[0]
port 520 nsew signal output
rlabel metal2 s 29458 219200 29514 220000 6 slave2_wb_adr_i[10]
port 521 nsew signal output
rlabel metal2 s 31390 219200 31446 220000 6 slave2_wb_adr_i[11]
port 522 nsew signal output
rlabel metal2 s 33322 219200 33378 220000 6 slave2_wb_adr_i[12]
port 523 nsew signal output
rlabel metal2 s 35254 219200 35310 220000 6 slave2_wb_adr_i[13]
port 524 nsew signal output
rlabel metal2 s 37186 219200 37242 220000 6 slave2_wb_adr_i[14]
port 525 nsew signal output
rlabel metal2 s 39118 219200 39174 220000 6 slave2_wb_adr_i[15]
port 526 nsew signal output
rlabel metal2 s 41050 219200 41106 220000 6 slave2_wb_adr_i[16]
port 527 nsew signal output
rlabel metal2 s 42982 219200 43038 220000 6 slave2_wb_adr_i[17]
port 528 nsew signal output
rlabel metal2 s 44914 219200 44970 220000 6 slave2_wb_adr_i[18]
port 529 nsew signal output
rlabel metal2 s 46846 219200 46902 220000 6 slave2_wb_adr_i[19]
port 530 nsew signal output
rlabel metal2 s 10138 219200 10194 220000 6 slave2_wb_adr_i[1]
port 531 nsew signal output
rlabel metal2 s 48778 219200 48834 220000 6 slave2_wb_adr_i[20]
port 532 nsew signal output
rlabel metal2 s 50710 219200 50766 220000 6 slave2_wb_adr_i[21]
port 533 nsew signal output
rlabel metal2 s 52642 219200 52698 220000 6 slave2_wb_adr_i[22]
port 534 nsew signal output
rlabel metal2 s 54574 219200 54630 220000 6 slave2_wb_adr_i[23]
port 535 nsew signal output
rlabel metal2 s 12714 219200 12770 220000 6 slave2_wb_adr_i[2]
port 536 nsew signal output
rlabel metal2 s 15290 219200 15346 220000 6 slave2_wb_adr_i[3]
port 537 nsew signal output
rlabel metal2 s 17866 219200 17922 220000 6 slave2_wb_adr_i[4]
port 538 nsew signal output
rlabel metal2 s 19798 219200 19854 220000 6 slave2_wb_adr_i[5]
port 539 nsew signal output
rlabel metal2 s 21730 219200 21786 220000 6 slave2_wb_adr_i[6]
port 540 nsew signal output
rlabel metal2 s 23662 219200 23718 220000 6 slave2_wb_adr_i[7]
port 541 nsew signal output
rlabel metal2 s 25594 219200 25650 220000 6 slave2_wb_adr_i[8]
port 542 nsew signal output
rlabel metal2 s 27526 219200 27582 220000 6 slave2_wb_adr_i[9]
port 543 nsew signal output
rlabel metal2 s 4342 219200 4398 220000 6 slave2_wb_cyc_i
port 544 nsew signal output
rlabel metal2 s 8206 219200 8262 220000 6 slave2_wb_data_i[0]
port 545 nsew signal output
rlabel metal2 s 30102 219200 30158 220000 6 slave2_wb_data_i[10]
port 546 nsew signal output
rlabel metal2 s 32034 219200 32090 220000 6 slave2_wb_data_i[11]
port 547 nsew signal output
rlabel metal2 s 33966 219200 34022 220000 6 slave2_wb_data_i[12]
port 548 nsew signal output
rlabel metal2 s 35898 219200 35954 220000 6 slave2_wb_data_i[13]
port 549 nsew signal output
rlabel metal2 s 37830 219200 37886 220000 6 slave2_wb_data_i[14]
port 550 nsew signal output
rlabel metal2 s 39762 219200 39818 220000 6 slave2_wb_data_i[15]
port 551 nsew signal output
rlabel metal2 s 41694 219200 41750 220000 6 slave2_wb_data_i[16]
port 552 nsew signal output
rlabel metal2 s 43626 219200 43682 220000 6 slave2_wb_data_i[17]
port 553 nsew signal output
rlabel metal2 s 45558 219200 45614 220000 6 slave2_wb_data_i[18]
port 554 nsew signal output
rlabel metal2 s 47490 219200 47546 220000 6 slave2_wb_data_i[19]
port 555 nsew signal output
rlabel metal2 s 10782 219200 10838 220000 6 slave2_wb_data_i[1]
port 556 nsew signal output
rlabel metal2 s 49422 219200 49478 220000 6 slave2_wb_data_i[20]
port 557 nsew signal output
rlabel metal2 s 51354 219200 51410 220000 6 slave2_wb_data_i[21]
port 558 nsew signal output
rlabel metal2 s 53286 219200 53342 220000 6 slave2_wb_data_i[22]
port 559 nsew signal output
rlabel metal2 s 55218 219200 55274 220000 6 slave2_wb_data_i[23]
port 560 nsew signal output
rlabel metal2 s 56506 219200 56562 220000 6 slave2_wb_data_i[24]
port 561 nsew signal output
rlabel metal2 s 57794 219200 57850 220000 6 slave2_wb_data_i[25]
port 562 nsew signal output
rlabel metal2 s 59082 219200 59138 220000 6 slave2_wb_data_i[26]
port 563 nsew signal output
rlabel metal2 s 60370 219200 60426 220000 6 slave2_wb_data_i[27]
port 564 nsew signal output
rlabel metal2 s 61658 219200 61714 220000 6 slave2_wb_data_i[28]
port 565 nsew signal output
rlabel metal2 s 62946 219200 63002 220000 6 slave2_wb_data_i[29]
port 566 nsew signal output
rlabel metal2 s 13358 219200 13414 220000 6 slave2_wb_data_i[2]
port 567 nsew signal output
rlabel metal2 s 64234 219200 64290 220000 6 slave2_wb_data_i[30]
port 568 nsew signal output
rlabel metal2 s 65522 219200 65578 220000 6 slave2_wb_data_i[31]
port 569 nsew signal output
rlabel metal2 s 15934 219200 15990 220000 6 slave2_wb_data_i[3]
port 570 nsew signal output
rlabel metal2 s 18510 219200 18566 220000 6 slave2_wb_data_i[4]
port 571 nsew signal output
rlabel metal2 s 20442 219200 20498 220000 6 slave2_wb_data_i[5]
port 572 nsew signal output
rlabel metal2 s 22374 219200 22430 220000 6 slave2_wb_data_i[6]
port 573 nsew signal output
rlabel metal2 s 24306 219200 24362 220000 6 slave2_wb_data_i[7]
port 574 nsew signal output
rlabel metal2 s 26238 219200 26294 220000 6 slave2_wb_data_i[8]
port 575 nsew signal output
rlabel metal2 s 28170 219200 28226 220000 6 slave2_wb_data_i[9]
port 576 nsew signal output
rlabel metal2 s 8850 219200 8906 220000 6 slave2_wb_data_o[0]
port 577 nsew signal input
rlabel metal2 s 30746 219200 30802 220000 6 slave2_wb_data_o[10]
port 578 nsew signal input
rlabel metal2 s 32678 219200 32734 220000 6 slave2_wb_data_o[11]
port 579 nsew signal input
rlabel metal2 s 34610 219200 34666 220000 6 slave2_wb_data_o[12]
port 580 nsew signal input
rlabel metal2 s 36542 219200 36598 220000 6 slave2_wb_data_o[13]
port 581 nsew signal input
rlabel metal2 s 38474 219200 38530 220000 6 slave2_wb_data_o[14]
port 582 nsew signal input
rlabel metal2 s 40406 219200 40462 220000 6 slave2_wb_data_o[15]
port 583 nsew signal input
rlabel metal2 s 42338 219200 42394 220000 6 slave2_wb_data_o[16]
port 584 nsew signal input
rlabel metal2 s 44270 219200 44326 220000 6 slave2_wb_data_o[17]
port 585 nsew signal input
rlabel metal2 s 46202 219200 46258 220000 6 slave2_wb_data_o[18]
port 586 nsew signal input
rlabel metal2 s 48134 219200 48190 220000 6 slave2_wb_data_o[19]
port 587 nsew signal input
rlabel metal2 s 11426 219200 11482 220000 6 slave2_wb_data_o[1]
port 588 nsew signal input
rlabel metal2 s 50066 219200 50122 220000 6 slave2_wb_data_o[20]
port 589 nsew signal input
rlabel metal2 s 51998 219200 52054 220000 6 slave2_wb_data_o[21]
port 590 nsew signal input
rlabel metal2 s 53930 219200 53986 220000 6 slave2_wb_data_o[22]
port 591 nsew signal input
rlabel metal2 s 55862 219200 55918 220000 6 slave2_wb_data_o[23]
port 592 nsew signal input
rlabel metal2 s 57150 219200 57206 220000 6 slave2_wb_data_o[24]
port 593 nsew signal input
rlabel metal2 s 58438 219200 58494 220000 6 slave2_wb_data_o[25]
port 594 nsew signal input
rlabel metal2 s 59726 219200 59782 220000 6 slave2_wb_data_o[26]
port 595 nsew signal input
rlabel metal2 s 61014 219200 61070 220000 6 slave2_wb_data_o[27]
port 596 nsew signal input
rlabel metal2 s 62302 219200 62358 220000 6 slave2_wb_data_o[28]
port 597 nsew signal input
rlabel metal2 s 63590 219200 63646 220000 6 slave2_wb_data_o[29]
port 598 nsew signal input
rlabel metal2 s 14002 219200 14058 220000 6 slave2_wb_data_o[2]
port 599 nsew signal input
rlabel metal2 s 64878 219200 64934 220000 6 slave2_wb_data_o[30]
port 600 nsew signal input
rlabel metal2 s 66166 219200 66222 220000 6 slave2_wb_data_o[31]
port 601 nsew signal input
rlabel metal2 s 16578 219200 16634 220000 6 slave2_wb_data_o[3]
port 602 nsew signal input
rlabel metal2 s 19154 219200 19210 220000 6 slave2_wb_data_o[4]
port 603 nsew signal input
rlabel metal2 s 21086 219200 21142 220000 6 slave2_wb_data_o[5]
port 604 nsew signal input
rlabel metal2 s 23018 219200 23074 220000 6 slave2_wb_data_o[6]
port 605 nsew signal input
rlabel metal2 s 24950 219200 25006 220000 6 slave2_wb_data_o[7]
port 606 nsew signal input
rlabel metal2 s 26882 219200 26938 220000 6 slave2_wb_data_o[8]
port 607 nsew signal input
rlabel metal2 s 28814 219200 28870 220000 6 slave2_wb_data_o[9]
port 608 nsew signal input
rlabel metal2 s 4986 219200 5042 220000 6 slave2_wb_error_o
port 609 nsew signal input
rlabel metal2 s 9494 219200 9550 220000 6 slave2_wb_sel_i[0]
port 610 nsew signal output
rlabel metal2 s 12070 219200 12126 220000 6 slave2_wb_sel_i[1]
port 611 nsew signal output
rlabel metal2 s 14646 219200 14702 220000 6 slave2_wb_sel_i[2]
port 612 nsew signal output
rlabel metal2 s 17222 219200 17278 220000 6 slave2_wb_sel_i[3]
port 613 nsew signal output
rlabel metal2 s 5630 219200 5686 220000 6 slave2_wb_stall_o
port 614 nsew signal input
rlabel metal2 s 6274 219200 6330 220000 6 slave2_wb_stb_i
port 615 nsew signal output
rlabel metal2 s 6918 219200 6974 220000 6 slave2_wb_we_i
port 616 nsew signal output
rlabel metal3 s 69200 110440 70000 110560 6 slave3_wb_ack_o
port 617 nsew signal input
rlabel metal3 s 69200 116968 70000 117088 6 slave3_wb_adr_i[0]
port 618 nsew signal output
rlabel metal3 s 69200 153960 70000 154080 6 slave3_wb_adr_i[10]
port 619 nsew signal output
rlabel metal3 s 69200 157224 70000 157344 6 slave3_wb_adr_i[11]
port 620 nsew signal output
rlabel metal3 s 69200 160488 70000 160608 6 slave3_wb_adr_i[12]
port 621 nsew signal output
rlabel metal3 s 69200 163752 70000 163872 6 slave3_wb_adr_i[13]
port 622 nsew signal output
rlabel metal3 s 69200 167016 70000 167136 6 slave3_wb_adr_i[14]
port 623 nsew signal output
rlabel metal3 s 69200 170280 70000 170400 6 slave3_wb_adr_i[15]
port 624 nsew signal output
rlabel metal3 s 69200 173544 70000 173664 6 slave3_wb_adr_i[16]
port 625 nsew signal output
rlabel metal3 s 69200 176808 70000 176928 6 slave3_wb_adr_i[17]
port 626 nsew signal output
rlabel metal3 s 69200 180072 70000 180192 6 slave3_wb_adr_i[18]
port 627 nsew signal output
rlabel metal3 s 69200 183336 70000 183456 6 slave3_wb_adr_i[19]
port 628 nsew signal output
rlabel metal3 s 69200 121320 70000 121440 6 slave3_wb_adr_i[1]
port 629 nsew signal output
rlabel metal3 s 69200 186600 70000 186720 6 slave3_wb_adr_i[20]
port 630 nsew signal output
rlabel metal3 s 69200 189864 70000 189984 6 slave3_wb_adr_i[21]
port 631 nsew signal output
rlabel metal3 s 69200 193128 70000 193248 6 slave3_wb_adr_i[22]
port 632 nsew signal output
rlabel metal3 s 69200 196392 70000 196512 6 slave3_wb_adr_i[23]
port 633 nsew signal output
rlabel metal3 s 69200 125672 70000 125792 6 slave3_wb_adr_i[2]
port 634 nsew signal output
rlabel metal3 s 69200 130024 70000 130144 6 slave3_wb_adr_i[3]
port 635 nsew signal output
rlabel metal3 s 69200 134376 70000 134496 6 slave3_wb_adr_i[4]
port 636 nsew signal output
rlabel metal3 s 69200 137640 70000 137760 6 slave3_wb_adr_i[5]
port 637 nsew signal output
rlabel metal3 s 69200 140904 70000 141024 6 slave3_wb_adr_i[6]
port 638 nsew signal output
rlabel metal3 s 69200 144168 70000 144288 6 slave3_wb_adr_i[7]
port 639 nsew signal output
rlabel metal3 s 69200 147432 70000 147552 6 slave3_wb_adr_i[8]
port 640 nsew signal output
rlabel metal3 s 69200 150696 70000 150816 6 slave3_wb_adr_i[9]
port 641 nsew signal output
rlabel metal3 s 69200 111528 70000 111648 6 slave3_wb_cyc_i
port 642 nsew signal output
rlabel metal3 s 69200 118056 70000 118176 6 slave3_wb_data_i[0]
port 643 nsew signal output
rlabel metal3 s 69200 155048 70000 155168 6 slave3_wb_data_i[10]
port 644 nsew signal output
rlabel metal3 s 69200 158312 70000 158432 6 slave3_wb_data_i[11]
port 645 nsew signal output
rlabel metal3 s 69200 161576 70000 161696 6 slave3_wb_data_i[12]
port 646 nsew signal output
rlabel metal3 s 69200 164840 70000 164960 6 slave3_wb_data_i[13]
port 647 nsew signal output
rlabel metal3 s 69200 168104 70000 168224 6 slave3_wb_data_i[14]
port 648 nsew signal output
rlabel metal3 s 69200 171368 70000 171488 6 slave3_wb_data_i[15]
port 649 nsew signal output
rlabel metal3 s 69200 174632 70000 174752 6 slave3_wb_data_i[16]
port 650 nsew signal output
rlabel metal3 s 69200 177896 70000 178016 6 slave3_wb_data_i[17]
port 651 nsew signal output
rlabel metal3 s 69200 181160 70000 181280 6 slave3_wb_data_i[18]
port 652 nsew signal output
rlabel metal3 s 69200 184424 70000 184544 6 slave3_wb_data_i[19]
port 653 nsew signal output
rlabel metal3 s 69200 122408 70000 122528 6 slave3_wb_data_i[1]
port 654 nsew signal output
rlabel metal3 s 69200 187688 70000 187808 6 slave3_wb_data_i[20]
port 655 nsew signal output
rlabel metal3 s 69200 190952 70000 191072 6 slave3_wb_data_i[21]
port 656 nsew signal output
rlabel metal3 s 69200 194216 70000 194336 6 slave3_wb_data_i[22]
port 657 nsew signal output
rlabel metal3 s 69200 197480 70000 197600 6 slave3_wb_data_i[23]
port 658 nsew signal output
rlabel metal3 s 69200 199656 70000 199776 6 slave3_wb_data_i[24]
port 659 nsew signal output
rlabel metal3 s 69200 201832 70000 201952 6 slave3_wb_data_i[25]
port 660 nsew signal output
rlabel metal3 s 69200 204008 70000 204128 6 slave3_wb_data_i[26]
port 661 nsew signal output
rlabel metal3 s 69200 206184 70000 206304 6 slave3_wb_data_i[27]
port 662 nsew signal output
rlabel metal3 s 69200 208360 70000 208480 6 slave3_wb_data_i[28]
port 663 nsew signal output
rlabel metal3 s 69200 210536 70000 210656 6 slave3_wb_data_i[29]
port 664 nsew signal output
rlabel metal3 s 69200 126760 70000 126880 6 slave3_wb_data_i[2]
port 665 nsew signal output
rlabel metal3 s 69200 212712 70000 212832 6 slave3_wb_data_i[30]
port 666 nsew signal output
rlabel metal3 s 69200 214888 70000 215008 6 slave3_wb_data_i[31]
port 667 nsew signal output
rlabel metal3 s 69200 131112 70000 131232 6 slave3_wb_data_i[3]
port 668 nsew signal output
rlabel metal3 s 69200 135464 70000 135584 6 slave3_wb_data_i[4]
port 669 nsew signal output
rlabel metal3 s 69200 138728 70000 138848 6 slave3_wb_data_i[5]
port 670 nsew signal output
rlabel metal3 s 69200 141992 70000 142112 6 slave3_wb_data_i[6]
port 671 nsew signal output
rlabel metal3 s 69200 145256 70000 145376 6 slave3_wb_data_i[7]
port 672 nsew signal output
rlabel metal3 s 69200 148520 70000 148640 6 slave3_wb_data_i[8]
port 673 nsew signal output
rlabel metal3 s 69200 151784 70000 151904 6 slave3_wb_data_i[9]
port 674 nsew signal output
rlabel metal3 s 69200 119144 70000 119264 6 slave3_wb_data_o[0]
port 675 nsew signal input
rlabel metal3 s 69200 156136 70000 156256 6 slave3_wb_data_o[10]
port 676 nsew signal input
rlabel metal3 s 69200 159400 70000 159520 6 slave3_wb_data_o[11]
port 677 nsew signal input
rlabel metal3 s 69200 162664 70000 162784 6 slave3_wb_data_o[12]
port 678 nsew signal input
rlabel metal3 s 69200 165928 70000 166048 6 slave3_wb_data_o[13]
port 679 nsew signal input
rlabel metal3 s 69200 169192 70000 169312 6 slave3_wb_data_o[14]
port 680 nsew signal input
rlabel metal3 s 69200 172456 70000 172576 6 slave3_wb_data_o[15]
port 681 nsew signal input
rlabel metal3 s 69200 175720 70000 175840 6 slave3_wb_data_o[16]
port 682 nsew signal input
rlabel metal3 s 69200 178984 70000 179104 6 slave3_wb_data_o[17]
port 683 nsew signal input
rlabel metal3 s 69200 182248 70000 182368 6 slave3_wb_data_o[18]
port 684 nsew signal input
rlabel metal3 s 69200 185512 70000 185632 6 slave3_wb_data_o[19]
port 685 nsew signal input
rlabel metal3 s 69200 123496 70000 123616 6 slave3_wb_data_o[1]
port 686 nsew signal input
rlabel metal3 s 69200 188776 70000 188896 6 slave3_wb_data_o[20]
port 687 nsew signal input
rlabel metal3 s 69200 192040 70000 192160 6 slave3_wb_data_o[21]
port 688 nsew signal input
rlabel metal3 s 69200 195304 70000 195424 6 slave3_wb_data_o[22]
port 689 nsew signal input
rlabel metal3 s 69200 198568 70000 198688 6 slave3_wb_data_o[23]
port 690 nsew signal input
rlabel metal3 s 69200 200744 70000 200864 6 slave3_wb_data_o[24]
port 691 nsew signal input
rlabel metal3 s 69200 202920 70000 203040 6 slave3_wb_data_o[25]
port 692 nsew signal input
rlabel metal3 s 69200 205096 70000 205216 6 slave3_wb_data_o[26]
port 693 nsew signal input
rlabel metal3 s 69200 207272 70000 207392 6 slave3_wb_data_o[27]
port 694 nsew signal input
rlabel metal3 s 69200 209448 70000 209568 6 slave3_wb_data_o[28]
port 695 nsew signal input
rlabel metal3 s 69200 211624 70000 211744 6 slave3_wb_data_o[29]
port 696 nsew signal input
rlabel metal3 s 69200 127848 70000 127968 6 slave3_wb_data_o[2]
port 697 nsew signal input
rlabel metal3 s 69200 213800 70000 213920 6 slave3_wb_data_o[30]
port 698 nsew signal input
rlabel metal3 s 69200 215976 70000 216096 6 slave3_wb_data_o[31]
port 699 nsew signal input
rlabel metal3 s 69200 132200 70000 132320 6 slave3_wb_data_o[3]
port 700 nsew signal input
rlabel metal3 s 69200 136552 70000 136672 6 slave3_wb_data_o[4]
port 701 nsew signal input
rlabel metal3 s 69200 139816 70000 139936 6 slave3_wb_data_o[5]
port 702 nsew signal input
rlabel metal3 s 69200 143080 70000 143200 6 slave3_wb_data_o[6]
port 703 nsew signal input
rlabel metal3 s 69200 146344 70000 146464 6 slave3_wb_data_o[7]
port 704 nsew signal input
rlabel metal3 s 69200 149608 70000 149728 6 slave3_wb_data_o[8]
port 705 nsew signal input
rlabel metal3 s 69200 152872 70000 152992 6 slave3_wb_data_o[9]
port 706 nsew signal input
rlabel metal3 s 69200 112616 70000 112736 6 slave3_wb_error_o
port 707 nsew signal input
rlabel metal3 s 69200 120232 70000 120352 6 slave3_wb_sel_i[0]
port 708 nsew signal output
rlabel metal3 s 69200 124584 70000 124704 6 slave3_wb_sel_i[1]
port 709 nsew signal output
rlabel metal3 s 69200 128936 70000 129056 6 slave3_wb_sel_i[2]
port 710 nsew signal output
rlabel metal3 s 69200 133288 70000 133408 6 slave3_wb_sel_i[3]
port 711 nsew signal output
rlabel metal3 s 69200 113704 70000 113824 6 slave3_wb_stall_o
port 712 nsew signal input
rlabel metal3 s 69200 114792 70000 114912 6 slave3_wb_stb_i
port 713 nsew signal output
rlabel metal3 s 69200 115880 70000 116000 6 slave3_wb_we_i
port 714 nsew signal output
rlabel metal3 s 69200 3816 70000 3936 6 slave4_wb_ack_o
port 715 nsew signal input
rlabel metal3 s 69200 10344 70000 10464 6 slave4_wb_adr_i[0]
port 716 nsew signal output
rlabel metal3 s 69200 47336 70000 47456 6 slave4_wb_adr_i[10]
port 717 nsew signal output
rlabel metal3 s 69200 50600 70000 50720 6 slave4_wb_adr_i[11]
port 718 nsew signal output
rlabel metal3 s 69200 53864 70000 53984 6 slave4_wb_adr_i[12]
port 719 nsew signal output
rlabel metal3 s 69200 57128 70000 57248 6 slave4_wb_adr_i[13]
port 720 nsew signal output
rlabel metal3 s 69200 60392 70000 60512 6 slave4_wb_adr_i[14]
port 721 nsew signal output
rlabel metal3 s 69200 63656 70000 63776 6 slave4_wb_adr_i[15]
port 722 nsew signal output
rlabel metal3 s 69200 66920 70000 67040 6 slave4_wb_adr_i[16]
port 723 nsew signal output
rlabel metal3 s 69200 70184 70000 70304 6 slave4_wb_adr_i[17]
port 724 nsew signal output
rlabel metal3 s 69200 73448 70000 73568 6 slave4_wb_adr_i[18]
port 725 nsew signal output
rlabel metal3 s 69200 76712 70000 76832 6 slave4_wb_adr_i[19]
port 726 nsew signal output
rlabel metal3 s 69200 14696 70000 14816 6 slave4_wb_adr_i[1]
port 727 nsew signal output
rlabel metal3 s 69200 79976 70000 80096 6 slave4_wb_adr_i[20]
port 728 nsew signal output
rlabel metal3 s 69200 83240 70000 83360 6 slave4_wb_adr_i[21]
port 729 nsew signal output
rlabel metal3 s 69200 86504 70000 86624 6 slave4_wb_adr_i[22]
port 730 nsew signal output
rlabel metal3 s 69200 89768 70000 89888 6 slave4_wb_adr_i[23]
port 731 nsew signal output
rlabel metal3 s 69200 19048 70000 19168 6 slave4_wb_adr_i[2]
port 732 nsew signal output
rlabel metal3 s 69200 23400 70000 23520 6 slave4_wb_adr_i[3]
port 733 nsew signal output
rlabel metal3 s 69200 27752 70000 27872 6 slave4_wb_adr_i[4]
port 734 nsew signal output
rlabel metal3 s 69200 31016 70000 31136 6 slave4_wb_adr_i[5]
port 735 nsew signal output
rlabel metal3 s 69200 34280 70000 34400 6 slave4_wb_adr_i[6]
port 736 nsew signal output
rlabel metal3 s 69200 37544 70000 37664 6 slave4_wb_adr_i[7]
port 737 nsew signal output
rlabel metal3 s 69200 40808 70000 40928 6 slave4_wb_adr_i[8]
port 738 nsew signal output
rlabel metal3 s 69200 44072 70000 44192 6 slave4_wb_adr_i[9]
port 739 nsew signal output
rlabel metal3 s 69200 4904 70000 5024 6 slave4_wb_cyc_i
port 740 nsew signal output
rlabel metal3 s 69200 11432 70000 11552 6 slave4_wb_data_i[0]
port 741 nsew signal output
rlabel metal3 s 69200 48424 70000 48544 6 slave4_wb_data_i[10]
port 742 nsew signal output
rlabel metal3 s 69200 51688 70000 51808 6 slave4_wb_data_i[11]
port 743 nsew signal output
rlabel metal3 s 69200 54952 70000 55072 6 slave4_wb_data_i[12]
port 744 nsew signal output
rlabel metal3 s 69200 58216 70000 58336 6 slave4_wb_data_i[13]
port 745 nsew signal output
rlabel metal3 s 69200 61480 70000 61600 6 slave4_wb_data_i[14]
port 746 nsew signal output
rlabel metal3 s 69200 64744 70000 64864 6 slave4_wb_data_i[15]
port 747 nsew signal output
rlabel metal3 s 69200 68008 70000 68128 6 slave4_wb_data_i[16]
port 748 nsew signal output
rlabel metal3 s 69200 71272 70000 71392 6 slave4_wb_data_i[17]
port 749 nsew signal output
rlabel metal3 s 69200 74536 70000 74656 6 slave4_wb_data_i[18]
port 750 nsew signal output
rlabel metal3 s 69200 77800 70000 77920 6 slave4_wb_data_i[19]
port 751 nsew signal output
rlabel metal3 s 69200 15784 70000 15904 6 slave4_wb_data_i[1]
port 752 nsew signal output
rlabel metal3 s 69200 81064 70000 81184 6 slave4_wb_data_i[20]
port 753 nsew signal output
rlabel metal3 s 69200 84328 70000 84448 6 slave4_wb_data_i[21]
port 754 nsew signal output
rlabel metal3 s 69200 87592 70000 87712 6 slave4_wb_data_i[22]
port 755 nsew signal output
rlabel metal3 s 69200 90856 70000 90976 6 slave4_wb_data_i[23]
port 756 nsew signal output
rlabel metal3 s 69200 93032 70000 93152 6 slave4_wb_data_i[24]
port 757 nsew signal output
rlabel metal3 s 69200 95208 70000 95328 6 slave4_wb_data_i[25]
port 758 nsew signal output
rlabel metal3 s 69200 97384 70000 97504 6 slave4_wb_data_i[26]
port 759 nsew signal output
rlabel metal3 s 69200 99560 70000 99680 6 slave4_wb_data_i[27]
port 760 nsew signal output
rlabel metal3 s 69200 101736 70000 101856 6 slave4_wb_data_i[28]
port 761 nsew signal output
rlabel metal3 s 69200 103912 70000 104032 6 slave4_wb_data_i[29]
port 762 nsew signal output
rlabel metal3 s 69200 20136 70000 20256 6 slave4_wb_data_i[2]
port 763 nsew signal output
rlabel metal3 s 69200 106088 70000 106208 6 slave4_wb_data_i[30]
port 764 nsew signal output
rlabel metal3 s 69200 108264 70000 108384 6 slave4_wb_data_i[31]
port 765 nsew signal output
rlabel metal3 s 69200 24488 70000 24608 6 slave4_wb_data_i[3]
port 766 nsew signal output
rlabel metal3 s 69200 28840 70000 28960 6 slave4_wb_data_i[4]
port 767 nsew signal output
rlabel metal3 s 69200 32104 70000 32224 6 slave4_wb_data_i[5]
port 768 nsew signal output
rlabel metal3 s 69200 35368 70000 35488 6 slave4_wb_data_i[6]
port 769 nsew signal output
rlabel metal3 s 69200 38632 70000 38752 6 slave4_wb_data_i[7]
port 770 nsew signal output
rlabel metal3 s 69200 41896 70000 42016 6 slave4_wb_data_i[8]
port 771 nsew signal output
rlabel metal3 s 69200 45160 70000 45280 6 slave4_wb_data_i[9]
port 772 nsew signal output
rlabel metal3 s 69200 12520 70000 12640 6 slave4_wb_data_o[0]
port 773 nsew signal input
rlabel metal3 s 69200 49512 70000 49632 6 slave4_wb_data_o[10]
port 774 nsew signal input
rlabel metal3 s 69200 52776 70000 52896 6 slave4_wb_data_o[11]
port 775 nsew signal input
rlabel metal3 s 69200 56040 70000 56160 6 slave4_wb_data_o[12]
port 776 nsew signal input
rlabel metal3 s 69200 59304 70000 59424 6 slave4_wb_data_o[13]
port 777 nsew signal input
rlabel metal3 s 69200 62568 70000 62688 6 slave4_wb_data_o[14]
port 778 nsew signal input
rlabel metal3 s 69200 65832 70000 65952 6 slave4_wb_data_o[15]
port 779 nsew signal input
rlabel metal3 s 69200 69096 70000 69216 6 slave4_wb_data_o[16]
port 780 nsew signal input
rlabel metal3 s 69200 72360 70000 72480 6 slave4_wb_data_o[17]
port 781 nsew signal input
rlabel metal3 s 69200 75624 70000 75744 6 slave4_wb_data_o[18]
port 782 nsew signal input
rlabel metal3 s 69200 78888 70000 79008 6 slave4_wb_data_o[19]
port 783 nsew signal input
rlabel metal3 s 69200 16872 70000 16992 6 slave4_wb_data_o[1]
port 784 nsew signal input
rlabel metal3 s 69200 82152 70000 82272 6 slave4_wb_data_o[20]
port 785 nsew signal input
rlabel metal3 s 69200 85416 70000 85536 6 slave4_wb_data_o[21]
port 786 nsew signal input
rlabel metal3 s 69200 88680 70000 88800 6 slave4_wb_data_o[22]
port 787 nsew signal input
rlabel metal3 s 69200 91944 70000 92064 6 slave4_wb_data_o[23]
port 788 nsew signal input
rlabel metal3 s 69200 94120 70000 94240 6 slave4_wb_data_o[24]
port 789 nsew signal input
rlabel metal3 s 69200 96296 70000 96416 6 slave4_wb_data_o[25]
port 790 nsew signal input
rlabel metal3 s 69200 98472 70000 98592 6 slave4_wb_data_o[26]
port 791 nsew signal input
rlabel metal3 s 69200 100648 70000 100768 6 slave4_wb_data_o[27]
port 792 nsew signal input
rlabel metal3 s 69200 102824 70000 102944 6 slave4_wb_data_o[28]
port 793 nsew signal input
rlabel metal3 s 69200 105000 70000 105120 6 slave4_wb_data_o[29]
port 794 nsew signal input
rlabel metal3 s 69200 21224 70000 21344 6 slave4_wb_data_o[2]
port 795 nsew signal input
rlabel metal3 s 69200 107176 70000 107296 6 slave4_wb_data_o[30]
port 796 nsew signal input
rlabel metal3 s 69200 109352 70000 109472 6 slave4_wb_data_o[31]
port 797 nsew signal input
rlabel metal3 s 69200 25576 70000 25696 6 slave4_wb_data_o[3]
port 798 nsew signal input
rlabel metal3 s 69200 29928 70000 30048 6 slave4_wb_data_o[4]
port 799 nsew signal input
rlabel metal3 s 69200 33192 70000 33312 6 slave4_wb_data_o[5]
port 800 nsew signal input
rlabel metal3 s 69200 36456 70000 36576 6 slave4_wb_data_o[6]
port 801 nsew signal input
rlabel metal3 s 69200 39720 70000 39840 6 slave4_wb_data_o[7]
port 802 nsew signal input
rlabel metal3 s 69200 42984 70000 43104 6 slave4_wb_data_o[8]
port 803 nsew signal input
rlabel metal3 s 69200 46248 70000 46368 6 slave4_wb_data_o[9]
port 804 nsew signal input
rlabel metal3 s 69200 5992 70000 6112 6 slave4_wb_error_o
port 805 nsew signal input
rlabel metal3 s 69200 13608 70000 13728 6 slave4_wb_sel_i[0]
port 806 nsew signal output
rlabel metal3 s 69200 17960 70000 18080 6 slave4_wb_sel_i[1]
port 807 nsew signal output
rlabel metal3 s 69200 22312 70000 22432 6 slave4_wb_sel_i[2]
port 808 nsew signal output
rlabel metal3 s 69200 26664 70000 26784 6 slave4_wb_sel_i[3]
port 809 nsew signal output
rlabel metal3 s 69200 7080 70000 7200 6 slave4_wb_stall_o
port 810 nsew signal input
rlabel metal3 s 69200 8168 70000 8288 6 slave4_wb_stb_i
port 811 nsew signal output
rlabel metal3 s 69200 9256 70000 9376 6 slave4_wb_we_i
port 812 nsew signal output
rlabel metal4 s 4208 2128 4528 217648 6 vccd1
port 813 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 217648 6 vccd1
port 813 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 217648 6 vccd1
port 813 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 217648 6 vssd1
port 814 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 217648 6 vssd1
port 814 nsew ground bidirectional
rlabel metal2 s 2134 0 2190 800 6 wb_clk_i
port 815 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wb_rst_i
port 816 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 220000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10824174
string GDS_FILE /mnt/f/WSL/ASIC/ExperiarSoC/openlane/WishboneInterconnect/runs/23_05_11_15_09/results/signoff/WishboneInterconnect.magic.gds
string GDS_START 698268
<< end >>

