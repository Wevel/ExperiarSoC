VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Peripherals
  CLASS BLOCK ;
  FOREIGN Peripherals ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 700.000 ;
  PIN flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END flash_csb
  PIN flash_io0_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END flash_io0_read
  PIN flash_io0_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END flash_io0_we
  PIN flash_io0_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END flash_io0_write
  PIN flash_io1_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END flash_io1_read
  PIN flash_io1_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END flash_io1_we
  PIN flash_io1_write
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END flash_io1_write
  PIN flash_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END flash_sck
  PIN internal_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END internal_uart_rx
  PIN internal_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END internal_uart_tx
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 696.000 2.670 700.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 696.000 160.450 700.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 696.000 176.090 700.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 696.000 191.730 700.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 696.000 207.830 700.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 696.000 223.470 700.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 696.000 239.110 700.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 696.000 255.210 700.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 696.000 270.850 700.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 696.000 286.490 700.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 696.000 302.590 700.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 696.000 18.310 700.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 696.000 318.230 700.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 696.000 333.870 700.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 696.000 349.510 700.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 696.000 365.610 700.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 696.000 381.250 700.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 696.000 396.890 700.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 696.000 412.990 700.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 696.000 428.630 700.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 696.000 444.270 700.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 696.000 460.370 700.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 696.000 33.950 700.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 696.000 476.010 700.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 696.000 491.650 700.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 696.000 507.750 700.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 696.000 523.390 700.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 696.000 539.030 700.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 696.000 555.130 700.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 696.000 570.770 700.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 696.000 586.410 700.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 696.000 49.590 700.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 696.000 65.690 700.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 696.000 81.330 700.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 696.000 96.970 700.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 696.000 113.070 700.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 696.000 128.710 700.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 696.000 144.350 700.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 696.000 7.730 700.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 696.000 165.510 700.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 696.000 181.150 700.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 696.000 197.250 700.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 696.000 212.890 700.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 696.000 228.530 700.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 696.000 244.630 700.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 696.000 260.270 700.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 696.000 275.910 700.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 696.000 292.010 700.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 696.000 307.650 700.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 696.000 23.370 700.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 696.000 323.290 700.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 696.000 339.390 700.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 696.000 355.030 700.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 696.000 370.670 700.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 696.000 386.770 700.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 696.000 402.410 700.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 696.000 418.050 700.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 696.000 433.690 700.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 696.000 449.790 700.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 696.000 465.430 700.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 696.000 39.470 700.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 696.000 481.070 700.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 696.000 497.170 700.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 696.000 512.810 700.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 696.000 528.450 700.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 696.000 544.550 700.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 696.000 560.190 700.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 696.000 575.830 700.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 696.000 591.930 700.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 696.000 55.110 700.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 696.000 70.750 700.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 696.000 86.850 700.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 696.000 102.490 700.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 696.000 118.130 700.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 696.000 133.770 700.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 696.000 149.870 700.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 696.000 12.790 700.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 696.000 171.030 700.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 696.000 186.670 700.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 696.000 202.310 700.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 696.000 217.950 700.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 696.000 234.050 700.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 696.000 249.690 700.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 696.000 265.330 700.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 696.000 281.430 700.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 696.000 297.070 700.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 696.000 312.710 700.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 696.000 28.890 700.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 696.000 328.810 700.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 696.000 344.450 700.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 696.000 360.090 700.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 696.000 376.190 700.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 696.000 391.830 700.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 696.000 407.470 700.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 696.000 423.570 700.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 696.000 439.210 700.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 696.000 454.850 700.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 696.000 470.950 700.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 696.000 44.530 700.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 696.000 486.590 700.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 696.000 502.230 700.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 696.000 517.870 700.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 696.000 533.970 700.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 696.000 549.610 700.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 696.000 565.250 700.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 696.000 581.350 700.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 696.000 596.990 700.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 696.000 60.170 700.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 696.000 76.270 700.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 696.000 91.910 700.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 696.000 107.550 700.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 696.000 123.650 700.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 696.000 139.290 700.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 696.000 154.930 700.000 ;
    END
  END io_out[9]
  PIN jtag_tck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 291.080 600.000 291.680 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 407.360 600.000 407.960 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 524.320 600.000 524.920 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 640.600 600.000 641.200 ;
    END
  END jtag_tms
  PIN probe_blink[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 57.840 600.000 58.440 ;
    END
  END probe_blink[0]
  PIN probe_blink[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 174.120 600.000 174.720 ;
    END
  END probe_blink[1]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 688.400 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.880 4.000 451.480 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.120 4.000 633.720 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.160 4.000 584.760 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 653.520 4.000 654.120 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.080 4.000 682.680 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.680 4.000 696.280 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 688.245 ;
      LAYER met1 ;
        RECT 5.520 10.640 597.010 689.480 ;
      LAYER met2 ;
        RECT 6.600 695.720 7.170 696.730 ;
        RECT 8.010 695.720 12.230 696.730 ;
        RECT 13.070 695.720 17.750 696.730 ;
        RECT 18.590 695.720 22.810 696.730 ;
        RECT 23.650 695.720 28.330 696.730 ;
        RECT 29.170 695.720 33.390 696.730 ;
        RECT 34.230 695.720 38.910 696.730 ;
        RECT 39.750 695.720 43.970 696.730 ;
        RECT 44.810 695.720 49.030 696.730 ;
        RECT 49.870 695.720 54.550 696.730 ;
        RECT 55.390 695.720 59.610 696.730 ;
        RECT 60.450 695.720 65.130 696.730 ;
        RECT 65.970 695.720 70.190 696.730 ;
        RECT 71.030 695.720 75.710 696.730 ;
        RECT 76.550 695.720 80.770 696.730 ;
        RECT 81.610 695.720 86.290 696.730 ;
        RECT 87.130 695.720 91.350 696.730 ;
        RECT 92.190 695.720 96.410 696.730 ;
        RECT 97.250 695.720 101.930 696.730 ;
        RECT 102.770 695.720 106.990 696.730 ;
        RECT 107.830 695.720 112.510 696.730 ;
        RECT 113.350 695.720 117.570 696.730 ;
        RECT 118.410 695.720 123.090 696.730 ;
        RECT 123.930 695.720 128.150 696.730 ;
        RECT 128.990 695.720 133.210 696.730 ;
        RECT 134.050 695.720 138.730 696.730 ;
        RECT 139.570 695.720 143.790 696.730 ;
        RECT 144.630 695.720 149.310 696.730 ;
        RECT 150.150 695.720 154.370 696.730 ;
        RECT 155.210 695.720 159.890 696.730 ;
        RECT 160.730 695.720 164.950 696.730 ;
        RECT 165.790 695.720 170.470 696.730 ;
        RECT 171.310 695.720 175.530 696.730 ;
        RECT 176.370 695.720 180.590 696.730 ;
        RECT 181.430 695.720 186.110 696.730 ;
        RECT 186.950 695.720 191.170 696.730 ;
        RECT 192.010 695.720 196.690 696.730 ;
        RECT 197.530 695.720 201.750 696.730 ;
        RECT 202.590 695.720 207.270 696.730 ;
        RECT 208.110 695.720 212.330 696.730 ;
        RECT 213.170 695.720 217.390 696.730 ;
        RECT 218.230 695.720 222.910 696.730 ;
        RECT 223.750 695.720 227.970 696.730 ;
        RECT 228.810 695.720 233.490 696.730 ;
        RECT 234.330 695.720 238.550 696.730 ;
        RECT 239.390 695.720 244.070 696.730 ;
        RECT 244.910 695.720 249.130 696.730 ;
        RECT 249.970 695.720 254.650 696.730 ;
        RECT 255.490 695.720 259.710 696.730 ;
        RECT 260.550 695.720 264.770 696.730 ;
        RECT 265.610 695.720 270.290 696.730 ;
        RECT 271.130 695.720 275.350 696.730 ;
        RECT 276.190 695.720 280.870 696.730 ;
        RECT 281.710 695.720 285.930 696.730 ;
        RECT 286.770 695.720 291.450 696.730 ;
        RECT 292.290 695.720 296.510 696.730 ;
        RECT 297.350 695.720 302.030 696.730 ;
        RECT 302.870 695.720 307.090 696.730 ;
        RECT 307.930 695.720 312.150 696.730 ;
        RECT 312.990 695.720 317.670 696.730 ;
        RECT 318.510 695.720 322.730 696.730 ;
        RECT 323.570 695.720 328.250 696.730 ;
        RECT 329.090 695.720 333.310 696.730 ;
        RECT 334.150 695.720 338.830 696.730 ;
        RECT 339.670 695.720 343.890 696.730 ;
        RECT 344.730 695.720 348.950 696.730 ;
        RECT 349.790 695.720 354.470 696.730 ;
        RECT 355.310 695.720 359.530 696.730 ;
        RECT 360.370 695.720 365.050 696.730 ;
        RECT 365.890 695.720 370.110 696.730 ;
        RECT 370.950 695.720 375.630 696.730 ;
        RECT 376.470 695.720 380.690 696.730 ;
        RECT 381.530 695.720 386.210 696.730 ;
        RECT 387.050 695.720 391.270 696.730 ;
        RECT 392.110 695.720 396.330 696.730 ;
        RECT 397.170 695.720 401.850 696.730 ;
        RECT 402.690 695.720 406.910 696.730 ;
        RECT 407.750 695.720 412.430 696.730 ;
        RECT 413.270 695.720 417.490 696.730 ;
        RECT 418.330 695.720 423.010 696.730 ;
        RECT 423.850 695.720 428.070 696.730 ;
        RECT 428.910 695.720 433.130 696.730 ;
        RECT 433.970 695.720 438.650 696.730 ;
        RECT 439.490 695.720 443.710 696.730 ;
        RECT 444.550 695.720 449.230 696.730 ;
        RECT 450.070 695.720 454.290 696.730 ;
        RECT 455.130 695.720 459.810 696.730 ;
        RECT 460.650 695.720 464.870 696.730 ;
        RECT 465.710 695.720 470.390 696.730 ;
        RECT 471.230 695.720 475.450 696.730 ;
        RECT 476.290 695.720 480.510 696.730 ;
        RECT 481.350 695.720 486.030 696.730 ;
        RECT 486.870 695.720 491.090 696.730 ;
        RECT 491.930 695.720 496.610 696.730 ;
        RECT 497.450 695.720 501.670 696.730 ;
        RECT 502.510 695.720 507.190 696.730 ;
        RECT 508.030 695.720 512.250 696.730 ;
        RECT 513.090 695.720 517.310 696.730 ;
        RECT 518.150 695.720 522.830 696.730 ;
        RECT 523.670 695.720 527.890 696.730 ;
        RECT 528.730 695.720 533.410 696.730 ;
        RECT 534.250 695.720 538.470 696.730 ;
        RECT 539.310 695.720 543.990 696.730 ;
        RECT 544.830 695.720 549.050 696.730 ;
        RECT 549.890 695.720 554.570 696.730 ;
        RECT 555.410 695.720 559.630 696.730 ;
        RECT 560.470 695.720 564.690 696.730 ;
        RECT 565.530 695.720 570.210 696.730 ;
        RECT 571.050 695.720 575.270 696.730 ;
        RECT 576.110 695.720 580.790 696.730 ;
        RECT 581.630 695.720 585.850 696.730 ;
        RECT 586.690 695.720 591.370 696.730 ;
        RECT 592.210 695.720 596.430 696.730 ;
        RECT 6.600 4.280 596.980 695.720 ;
        RECT 6.600 3.555 16.370 4.280 ;
        RECT 17.210 3.555 49.490 4.280 ;
        RECT 50.330 3.555 82.610 4.280 ;
        RECT 83.450 3.555 116.190 4.280 ;
        RECT 117.030 3.555 149.310 4.280 ;
        RECT 150.150 3.555 182.890 4.280 ;
        RECT 183.730 3.555 216.010 4.280 ;
        RECT 216.850 3.555 249.590 4.280 ;
        RECT 250.430 3.555 282.710 4.280 ;
        RECT 283.550 3.555 316.290 4.280 ;
        RECT 317.130 3.555 349.410 4.280 ;
        RECT 350.250 3.555 382.530 4.280 ;
        RECT 383.370 3.555 416.110 4.280 ;
        RECT 416.950 3.555 449.230 4.280 ;
        RECT 450.070 3.555 482.810 4.280 ;
        RECT 483.650 3.555 515.930 4.280 ;
        RECT 516.770 3.555 549.510 4.280 ;
        RECT 550.350 3.555 582.630 4.280 ;
        RECT 583.470 3.555 596.980 4.280 ;
      LAYER met3 ;
        RECT 4.400 695.280 596.000 696.145 ;
        RECT 4.000 689.880 596.000 695.280 ;
        RECT 4.400 688.480 596.000 689.880 ;
        RECT 4.000 683.080 596.000 688.480 ;
        RECT 4.400 681.680 596.000 683.080 ;
        RECT 4.000 675.600 596.000 681.680 ;
        RECT 4.400 674.200 596.000 675.600 ;
        RECT 4.000 668.800 596.000 674.200 ;
        RECT 4.400 667.400 596.000 668.800 ;
        RECT 4.000 662.000 596.000 667.400 ;
        RECT 4.400 660.600 596.000 662.000 ;
        RECT 4.000 654.520 596.000 660.600 ;
        RECT 4.400 653.120 596.000 654.520 ;
        RECT 4.000 647.720 596.000 653.120 ;
        RECT 4.400 646.320 596.000 647.720 ;
        RECT 4.000 641.600 596.000 646.320 ;
        RECT 4.000 640.920 595.600 641.600 ;
        RECT 4.400 640.200 595.600 640.920 ;
        RECT 4.400 639.520 596.000 640.200 ;
        RECT 4.000 634.120 596.000 639.520 ;
        RECT 4.400 632.720 596.000 634.120 ;
        RECT 4.000 626.640 596.000 632.720 ;
        RECT 4.400 625.240 596.000 626.640 ;
        RECT 4.000 619.840 596.000 625.240 ;
        RECT 4.400 618.440 596.000 619.840 ;
        RECT 4.000 613.040 596.000 618.440 ;
        RECT 4.400 611.640 596.000 613.040 ;
        RECT 4.000 605.560 596.000 611.640 ;
        RECT 4.400 604.160 596.000 605.560 ;
        RECT 4.000 598.760 596.000 604.160 ;
        RECT 4.400 597.360 596.000 598.760 ;
        RECT 4.000 591.960 596.000 597.360 ;
        RECT 4.400 590.560 596.000 591.960 ;
        RECT 4.000 585.160 596.000 590.560 ;
        RECT 4.400 583.760 596.000 585.160 ;
        RECT 4.000 577.680 596.000 583.760 ;
        RECT 4.400 576.280 596.000 577.680 ;
        RECT 4.000 570.880 596.000 576.280 ;
        RECT 4.400 569.480 596.000 570.880 ;
        RECT 4.000 564.080 596.000 569.480 ;
        RECT 4.400 562.680 596.000 564.080 ;
        RECT 4.000 556.600 596.000 562.680 ;
        RECT 4.400 555.200 596.000 556.600 ;
        RECT 4.000 549.800 596.000 555.200 ;
        RECT 4.400 548.400 596.000 549.800 ;
        RECT 4.000 543.000 596.000 548.400 ;
        RECT 4.400 541.600 596.000 543.000 ;
        RECT 4.000 536.200 596.000 541.600 ;
        RECT 4.400 534.800 596.000 536.200 ;
        RECT 4.000 528.720 596.000 534.800 ;
        RECT 4.400 527.320 596.000 528.720 ;
        RECT 4.000 525.320 596.000 527.320 ;
        RECT 4.000 523.920 595.600 525.320 ;
        RECT 4.000 521.920 596.000 523.920 ;
        RECT 4.400 520.520 596.000 521.920 ;
        RECT 4.000 515.120 596.000 520.520 ;
        RECT 4.400 513.720 596.000 515.120 ;
        RECT 4.000 507.640 596.000 513.720 ;
        RECT 4.400 506.240 596.000 507.640 ;
        RECT 4.000 500.840 596.000 506.240 ;
        RECT 4.400 499.440 596.000 500.840 ;
        RECT 4.000 494.040 596.000 499.440 ;
        RECT 4.400 492.640 596.000 494.040 ;
        RECT 4.000 487.240 596.000 492.640 ;
        RECT 4.400 485.840 596.000 487.240 ;
        RECT 4.000 479.760 596.000 485.840 ;
        RECT 4.400 478.360 596.000 479.760 ;
        RECT 4.000 472.960 596.000 478.360 ;
        RECT 4.400 471.560 596.000 472.960 ;
        RECT 4.000 466.160 596.000 471.560 ;
        RECT 4.400 464.760 596.000 466.160 ;
        RECT 4.000 458.680 596.000 464.760 ;
        RECT 4.400 457.280 596.000 458.680 ;
        RECT 4.000 451.880 596.000 457.280 ;
        RECT 4.400 450.480 596.000 451.880 ;
        RECT 4.000 445.080 596.000 450.480 ;
        RECT 4.400 443.680 596.000 445.080 ;
        RECT 4.000 437.600 596.000 443.680 ;
        RECT 4.400 436.200 596.000 437.600 ;
        RECT 4.000 430.800 596.000 436.200 ;
        RECT 4.400 429.400 596.000 430.800 ;
        RECT 4.000 424.000 596.000 429.400 ;
        RECT 4.400 422.600 596.000 424.000 ;
        RECT 4.000 417.200 596.000 422.600 ;
        RECT 4.400 415.800 596.000 417.200 ;
        RECT 4.000 409.720 596.000 415.800 ;
        RECT 4.400 408.360 596.000 409.720 ;
        RECT 4.400 408.320 595.600 408.360 ;
        RECT 4.000 406.960 595.600 408.320 ;
        RECT 4.000 402.920 596.000 406.960 ;
        RECT 4.400 401.520 596.000 402.920 ;
        RECT 4.000 396.120 596.000 401.520 ;
        RECT 4.400 394.720 596.000 396.120 ;
        RECT 4.000 388.640 596.000 394.720 ;
        RECT 4.400 387.240 596.000 388.640 ;
        RECT 4.000 381.840 596.000 387.240 ;
        RECT 4.400 380.440 596.000 381.840 ;
        RECT 4.000 375.040 596.000 380.440 ;
        RECT 4.400 373.640 596.000 375.040 ;
        RECT 4.000 368.240 596.000 373.640 ;
        RECT 4.400 366.840 596.000 368.240 ;
        RECT 4.000 360.760 596.000 366.840 ;
        RECT 4.400 359.360 596.000 360.760 ;
        RECT 4.000 353.960 596.000 359.360 ;
        RECT 4.400 352.560 596.000 353.960 ;
        RECT 4.000 347.160 596.000 352.560 ;
        RECT 4.400 345.760 596.000 347.160 ;
        RECT 4.000 339.680 596.000 345.760 ;
        RECT 4.400 338.280 596.000 339.680 ;
        RECT 4.000 332.880 596.000 338.280 ;
        RECT 4.400 331.480 596.000 332.880 ;
        RECT 4.000 326.080 596.000 331.480 ;
        RECT 4.400 324.680 596.000 326.080 ;
        RECT 4.000 319.280 596.000 324.680 ;
        RECT 4.400 317.880 596.000 319.280 ;
        RECT 4.000 311.800 596.000 317.880 ;
        RECT 4.400 310.400 596.000 311.800 ;
        RECT 4.000 305.000 596.000 310.400 ;
        RECT 4.400 303.600 596.000 305.000 ;
        RECT 4.000 298.200 596.000 303.600 ;
        RECT 4.400 296.800 596.000 298.200 ;
        RECT 4.000 292.080 596.000 296.800 ;
        RECT 4.000 290.720 595.600 292.080 ;
        RECT 4.400 290.680 595.600 290.720 ;
        RECT 4.400 289.320 596.000 290.680 ;
        RECT 4.000 283.920 596.000 289.320 ;
        RECT 4.400 282.520 596.000 283.920 ;
        RECT 4.000 277.120 596.000 282.520 ;
        RECT 4.400 275.720 596.000 277.120 ;
        RECT 4.000 270.320 596.000 275.720 ;
        RECT 4.400 268.920 596.000 270.320 ;
        RECT 4.000 262.840 596.000 268.920 ;
        RECT 4.400 261.440 596.000 262.840 ;
        RECT 4.000 256.040 596.000 261.440 ;
        RECT 4.400 254.640 596.000 256.040 ;
        RECT 4.000 249.240 596.000 254.640 ;
        RECT 4.400 247.840 596.000 249.240 ;
        RECT 4.000 241.760 596.000 247.840 ;
        RECT 4.400 240.360 596.000 241.760 ;
        RECT 4.000 234.960 596.000 240.360 ;
        RECT 4.400 233.560 596.000 234.960 ;
        RECT 4.000 228.160 596.000 233.560 ;
        RECT 4.400 226.760 596.000 228.160 ;
        RECT 4.000 220.680 596.000 226.760 ;
        RECT 4.400 219.280 596.000 220.680 ;
        RECT 4.000 213.880 596.000 219.280 ;
        RECT 4.400 212.480 596.000 213.880 ;
        RECT 4.000 207.080 596.000 212.480 ;
        RECT 4.400 205.680 596.000 207.080 ;
        RECT 4.000 200.280 596.000 205.680 ;
        RECT 4.400 198.880 596.000 200.280 ;
        RECT 4.000 192.800 596.000 198.880 ;
        RECT 4.400 191.400 596.000 192.800 ;
        RECT 4.000 186.000 596.000 191.400 ;
        RECT 4.400 184.600 596.000 186.000 ;
        RECT 4.000 179.200 596.000 184.600 ;
        RECT 4.400 177.800 596.000 179.200 ;
        RECT 4.000 175.120 596.000 177.800 ;
        RECT 4.000 173.720 595.600 175.120 ;
        RECT 4.000 171.720 596.000 173.720 ;
        RECT 4.400 170.320 596.000 171.720 ;
        RECT 4.000 164.920 596.000 170.320 ;
        RECT 4.400 163.520 596.000 164.920 ;
        RECT 4.000 158.120 596.000 163.520 ;
        RECT 4.400 156.720 596.000 158.120 ;
        RECT 4.000 151.320 596.000 156.720 ;
        RECT 4.400 149.920 596.000 151.320 ;
        RECT 4.000 143.840 596.000 149.920 ;
        RECT 4.400 142.440 596.000 143.840 ;
        RECT 4.000 137.040 596.000 142.440 ;
        RECT 4.400 135.640 596.000 137.040 ;
        RECT 4.000 130.240 596.000 135.640 ;
        RECT 4.400 128.840 596.000 130.240 ;
        RECT 4.000 122.760 596.000 128.840 ;
        RECT 4.400 121.360 596.000 122.760 ;
        RECT 4.000 115.960 596.000 121.360 ;
        RECT 4.400 114.560 596.000 115.960 ;
        RECT 4.000 109.160 596.000 114.560 ;
        RECT 4.400 107.760 596.000 109.160 ;
        RECT 4.000 102.360 596.000 107.760 ;
        RECT 4.400 100.960 596.000 102.360 ;
        RECT 4.000 94.880 596.000 100.960 ;
        RECT 4.400 93.480 596.000 94.880 ;
        RECT 4.000 88.080 596.000 93.480 ;
        RECT 4.400 86.680 596.000 88.080 ;
        RECT 4.000 81.280 596.000 86.680 ;
        RECT 4.400 79.880 596.000 81.280 ;
        RECT 4.000 73.800 596.000 79.880 ;
        RECT 4.400 72.400 596.000 73.800 ;
        RECT 4.000 67.000 596.000 72.400 ;
        RECT 4.400 65.600 596.000 67.000 ;
        RECT 4.000 60.200 596.000 65.600 ;
        RECT 4.400 58.840 596.000 60.200 ;
        RECT 4.400 58.800 595.600 58.840 ;
        RECT 4.000 57.440 595.600 58.800 ;
        RECT 4.000 53.400 596.000 57.440 ;
        RECT 4.400 52.000 596.000 53.400 ;
        RECT 4.000 45.920 596.000 52.000 ;
        RECT 4.400 44.520 596.000 45.920 ;
        RECT 4.000 39.120 596.000 44.520 ;
        RECT 4.400 37.720 596.000 39.120 ;
        RECT 4.000 32.320 596.000 37.720 ;
        RECT 4.400 30.920 596.000 32.320 ;
        RECT 4.000 24.840 596.000 30.920 ;
        RECT 4.400 23.440 596.000 24.840 ;
        RECT 4.000 18.040 596.000 23.440 ;
        RECT 4.400 16.640 596.000 18.040 ;
        RECT 4.000 11.240 596.000 16.640 ;
        RECT 4.400 9.840 596.000 11.240 ;
        RECT 4.000 4.440 596.000 9.840 ;
        RECT 4.400 3.575 596.000 4.440 ;
      LAYER met4 ;
        RECT 24.215 34.175 97.440 611.145 ;
        RECT 99.840 34.175 174.240 611.145 ;
        RECT 176.640 34.175 251.040 611.145 ;
        RECT 253.440 34.175 327.840 611.145 ;
        RECT 330.240 34.175 404.640 611.145 ;
        RECT 407.040 34.175 481.440 611.145 ;
        RECT 483.840 34.175 543.425 611.145 ;
  END
END Peripherals
END LIBRARY

