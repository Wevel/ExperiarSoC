magic
tech sky130A
magscale 1 2
timestamp 1652641936
<< obsli1 >>
rect 1104 2159 68816 197489
<< obsm1 >>
rect 290 1912 69722 197520
<< metal2 >>
rect 294 199200 350 200000
rect 938 199200 994 200000
rect 1674 199200 1730 200000
rect 2410 199200 2466 200000
rect 3146 199200 3202 200000
rect 3790 199200 3846 200000
rect 4526 199200 4582 200000
rect 5262 199200 5318 200000
rect 5998 199200 6054 200000
rect 6642 199200 6698 200000
rect 7378 199200 7434 200000
rect 8114 199200 8170 200000
rect 8850 199200 8906 200000
rect 9494 199200 9550 200000
rect 10230 199200 10286 200000
rect 10966 199200 11022 200000
rect 11702 199200 11758 200000
rect 12438 199200 12494 200000
rect 13082 199200 13138 200000
rect 13818 199200 13874 200000
rect 14554 199200 14610 200000
rect 15290 199200 15346 200000
rect 15934 199200 15990 200000
rect 16670 199200 16726 200000
rect 17406 199200 17462 200000
rect 18142 199200 18198 200000
rect 18786 199200 18842 200000
rect 19522 199200 19578 200000
rect 20258 199200 20314 200000
rect 20994 199200 21050 200000
rect 21638 199200 21694 200000
rect 22374 199200 22430 200000
rect 23110 199200 23166 200000
rect 23846 199200 23902 200000
rect 24582 199200 24638 200000
rect 25226 199200 25282 200000
rect 25962 199200 26018 200000
rect 26698 199200 26754 200000
rect 27434 199200 27490 200000
rect 28078 199200 28134 200000
rect 28814 199200 28870 200000
rect 29550 199200 29606 200000
rect 30286 199200 30342 200000
rect 30930 199200 30986 200000
rect 31666 199200 31722 200000
rect 32402 199200 32458 200000
rect 33138 199200 33194 200000
rect 33782 199200 33838 200000
rect 34518 199200 34574 200000
rect 35254 199200 35310 200000
rect 35990 199200 36046 200000
rect 36726 199200 36782 200000
rect 37370 199200 37426 200000
rect 38106 199200 38162 200000
rect 38842 199200 38898 200000
rect 39578 199200 39634 200000
rect 40222 199200 40278 200000
rect 40958 199200 41014 200000
rect 41694 199200 41750 200000
rect 42430 199200 42486 200000
rect 43074 199200 43130 200000
rect 43810 199200 43866 200000
rect 44546 199200 44602 200000
rect 45282 199200 45338 200000
rect 45926 199200 45982 200000
rect 46662 199200 46718 200000
rect 47398 199200 47454 200000
rect 48134 199200 48190 200000
rect 48870 199200 48926 200000
rect 49514 199200 49570 200000
rect 50250 199200 50306 200000
rect 50986 199200 51042 200000
rect 51722 199200 51778 200000
rect 52366 199200 52422 200000
rect 53102 199200 53158 200000
rect 53838 199200 53894 200000
rect 54574 199200 54630 200000
rect 55218 199200 55274 200000
rect 55954 199200 56010 200000
rect 56690 199200 56746 200000
rect 57426 199200 57482 200000
rect 58070 199200 58126 200000
rect 58806 199200 58862 200000
rect 59542 199200 59598 200000
rect 60278 199200 60334 200000
rect 61014 199200 61070 200000
rect 61658 199200 61714 200000
rect 62394 199200 62450 200000
rect 63130 199200 63186 200000
rect 63866 199200 63922 200000
rect 64510 199200 64566 200000
rect 65246 199200 65302 200000
rect 65982 199200 66038 200000
rect 66718 199200 66774 200000
rect 67362 199200 67418 200000
rect 68098 199200 68154 200000
rect 68834 199200 68890 200000
rect 69570 199200 69626 200000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3790 0 3846 800
rect 4342 0 4398 800
rect 4894 0 4950 800
rect 5538 0 5594 800
rect 6090 0 6146 800
rect 6642 0 6698 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9586 0 9642 800
rect 10138 0 10194 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 16026 0 16082 800
rect 16578 0 16634 800
rect 17130 0 17186 800
rect 17774 0 17830 800
rect 18326 0 18382 800
rect 18878 0 18934 800
rect 19522 0 19578 800
rect 20074 0 20130 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21822 0 21878 800
rect 22374 0 22430 800
rect 23018 0 23074 800
rect 23570 0 23626 800
rect 24214 0 24270 800
rect 24766 0 24822 800
rect 25318 0 25374 800
rect 25962 0 26018 800
rect 26514 0 26570 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29458 0 29514 800
rect 30010 0 30066 800
rect 30562 0 30618 800
rect 31206 0 31262 800
rect 31758 0 31814 800
rect 32310 0 32366 800
rect 32954 0 33010 800
rect 33506 0 33562 800
rect 34058 0 34114 800
rect 34702 0 34758 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36450 0 36506 800
rect 37002 0 37058 800
rect 37554 0 37610 800
rect 38198 0 38254 800
rect 38750 0 38806 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 41050 0 41106 800
rect 41694 0 41750 800
rect 42246 0 42302 800
rect 42798 0 42854 800
rect 43442 0 43498 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 45190 0 45246 800
rect 45742 0 45798 800
rect 46294 0 46350 800
rect 46938 0 46994 800
rect 47490 0 47546 800
rect 48134 0 48190 800
rect 48686 0 48742 800
rect 49238 0 49294 800
rect 49882 0 49938 800
rect 50434 0 50490 800
rect 50986 0 51042 800
rect 51630 0 51686 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53378 0 53434 800
rect 53930 0 53986 800
rect 54482 0 54538 800
rect 55126 0 55182 800
rect 55678 0 55734 800
rect 56230 0 56286 800
rect 56874 0 56930 800
rect 57426 0 57482 800
rect 57978 0 58034 800
rect 58622 0 58678 800
rect 59174 0 59230 800
rect 59726 0 59782 800
rect 60370 0 60426 800
rect 60922 0 60978 800
rect 61474 0 61530 800
rect 62118 0 62174 800
rect 62670 0 62726 800
rect 63222 0 63278 800
rect 63866 0 63922 800
rect 64418 0 64474 800
rect 64970 0 65026 800
rect 65614 0 65670 800
rect 66166 0 66222 800
rect 66718 0 66774 800
rect 67362 0 67418 800
rect 67914 0 67970 800
rect 68466 0 68522 800
rect 69110 0 69166 800
rect 69662 0 69718 800
<< obsm2 >>
rect 406 199144 882 199753
rect 1050 199144 1618 199753
rect 1786 199144 2354 199753
rect 2522 199144 3090 199753
rect 3258 199144 3734 199753
rect 3902 199144 4470 199753
rect 4638 199144 5206 199753
rect 5374 199144 5942 199753
rect 6110 199144 6586 199753
rect 6754 199144 7322 199753
rect 7490 199144 8058 199753
rect 8226 199144 8794 199753
rect 8962 199144 9438 199753
rect 9606 199144 10174 199753
rect 10342 199144 10910 199753
rect 11078 199144 11646 199753
rect 11814 199144 12382 199753
rect 12550 199144 13026 199753
rect 13194 199144 13762 199753
rect 13930 199144 14498 199753
rect 14666 199144 15234 199753
rect 15402 199144 15878 199753
rect 16046 199144 16614 199753
rect 16782 199144 17350 199753
rect 17518 199144 18086 199753
rect 18254 199144 18730 199753
rect 18898 199144 19466 199753
rect 19634 199144 20202 199753
rect 20370 199144 20938 199753
rect 21106 199144 21582 199753
rect 21750 199144 22318 199753
rect 22486 199144 23054 199753
rect 23222 199144 23790 199753
rect 23958 199144 24526 199753
rect 24694 199144 25170 199753
rect 25338 199144 25906 199753
rect 26074 199144 26642 199753
rect 26810 199144 27378 199753
rect 27546 199144 28022 199753
rect 28190 199144 28758 199753
rect 28926 199144 29494 199753
rect 29662 199144 30230 199753
rect 30398 199144 30874 199753
rect 31042 199144 31610 199753
rect 31778 199144 32346 199753
rect 32514 199144 33082 199753
rect 33250 199144 33726 199753
rect 33894 199144 34462 199753
rect 34630 199144 35198 199753
rect 35366 199144 35934 199753
rect 36102 199144 36670 199753
rect 36838 199144 37314 199753
rect 37482 199144 38050 199753
rect 38218 199144 38786 199753
rect 38954 199144 39522 199753
rect 39690 199144 40166 199753
rect 40334 199144 40902 199753
rect 41070 199144 41638 199753
rect 41806 199144 42374 199753
rect 42542 199144 43018 199753
rect 43186 199144 43754 199753
rect 43922 199144 44490 199753
rect 44658 199144 45226 199753
rect 45394 199144 45870 199753
rect 46038 199144 46606 199753
rect 46774 199144 47342 199753
rect 47510 199144 48078 199753
rect 48246 199144 48814 199753
rect 48982 199144 49458 199753
rect 49626 199144 50194 199753
rect 50362 199144 50930 199753
rect 51098 199144 51666 199753
rect 51834 199144 52310 199753
rect 52478 199144 53046 199753
rect 53214 199144 53782 199753
rect 53950 199144 54518 199753
rect 54686 199144 55162 199753
rect 55330 199144 55898 199753
rect 56066 199144 56634 199753
rect 56802 199144 57370 199753
rect 57538 199144 58014 199753
rect 58182 199144 58750 199753
rect 58918 199144 59486 199753
rect 59654 199144 60222 199753
rect 60390 199144 60958 199753
rect 61126 199144 61602 199753
rect 61770 199144 62338 199753
rect 62506 199144 63074 199753
rect 63242 199144 63810 199753
rect 63978 199144 64454 199753
rect 64622 199144 65190 199753
rect 65358 199144 65926 199753
rect 66094 199144 66662 199753
rect 66830 199144 67306 199753
rect 67474 199144 68042 199753
rect 68210 199144 68778 199753
rect 68946 199144 69514 199753
rect 69682 199144 69716 199753
rect 296 856 69716 199144
rect 406 167 790 856
rect 958 167 1342 856
rect 1510 167 1986 856
rect 2154 167 2538 856
rect 2706 167 3090 856
rect 3258 167 3734 856
rect 3902 167 4286 856
rect 4454 167 4838 856
rect 5006 167 5482 856
rect 5650 167 6034 856
rect 6202 167 6586 856
rect 6754 167 7230 856
rect 7398 167 7782 856
rect 7950 167 8334 856
rect 8502 167 8978 856
rect 9146 167 9530 856
rect 9698 167 10082 856
rect 10250 167 10726 856
rect 10894 167 11278 856
rect 11446 167 11830 856
rect 11998 167 12474 856
rect 12642 167 13026 856
rect 13194 167 13578 856
rect 13746 167 14222 856
rect 14390 167 14774 856
rect 14942 167 15326 856
rect 15494 167 15970 856
rect 16138 167 16522 856
rect 16690 167 17074 856
rect 17242 167 17718 856
rect 17886 167 18270 856
rect 18438 167 18822 856
rect 18990 167 19466 856
rect 19634 167 20018 856
rect 20186 167 20570 856
rect 20738 167 21214 856
rect 21382 167 21766 856
rect 21934 167 22318 856
rect 22486 167 22962 856
rect 23130 167 23514 856
rect 23682 167 24158 856
rect 24326 167 24710 856
rect 24878 167 25262 856
rect 25430 167 25906 856
rect 26074 167 26458 856
rect 26626 167 27010 856
rect 27178 167 27654 856
rect 27822 167 28206 856
rect 28374 167 28758 856
rect 28926 167 29402 856
rect 29570 167 29954 856
rect 30122 167 30506 856
rect 30674 167 31150 856
rect 31318 167 31702 856
rect 31870 167 32254 856
rect 32422 167 32898 856
rect 33066 167 33450 856
rect 33618 167 34002 856
rect 34170 167 34646 856
rect 34814 167 35198 856
rect 35366 167 35750 856
rect 35918 167 36394 856
rect 36562 167 36946 856
rect 37114 167 37498 856
rect 37666 167 38142 856
rect 38310 167 38694 856
rect 38862 167 39246 856
rect 39414 167 39890 856
rect 40058 167 40442 856
rect 40610 167 40994 856
rect 41162 167 41638 856
rect 41806 167 42190 856
rect 42358 167 42742 856
rect 42910 167 43386 856
rect 43554 167 43938 856
rect 44106 167 44490 856
rect 44658 167 45134 856
rect 45302 167 45686 856
rect 45854 167 46238 856
rect 46406 167 46882 856
rect 47050 167 47434 856
rect 47602 167 48078 856
rect 48246 167 48630 856
rect 48798 167 49182 856
rect 49350 167 49826 856
rect 49994 167 50378 856
rect 50546 167 50930 856
rect 51098 167 51574 856
rect 51742 167 52126 856
rect 52294 167 52678 856
rect 52846 167 53322 856
rect 53490 167 53874 856
rect 54042 167 54426 856
rect 54594 167 55070 856
rect 55238 167 55622 856
rect 55790 167 56174 856
rect 56342 167 56818 856
rect 56986 167 57370 856
rect 57538 167 57922 856
rect 58090 167 58566 856
rect 58734 167 59118 856
rect 59286 167 59670 856
rect 59838 167 60314 856
rect 60482 167 60866 856
rect 61034 167 61418 856
rect 61586 167 62062 856
rect 62230 167 62614 856
rect 62782 167 63166 856
rect 63334 167 63810 856
rect 63978 167 64362 856
rect 64530 167 64914 856
rect 65082 167 65558 856
rect 65726 167 66110 856
rect 66278 167 66662 856
rect 66830 167 67306 856
rect 67474 167 67858 856
rect 68026 167 68410 856
rect 68578 167 69054 856
rect 69222 167 69606 856
<< metal3 >>
rect 0 199656 800 199776
rect 0 199112 800 199232
rect 69200 198840 70000 198960
rect 0 198568 800 198688
rect 0 198160 800 198280
rect 0 197616 800 197736
rect 0 197072 800 197192
rect 0 196664 800 196784
rect 69200 196800 70000 196920
rect 0 196120 800 196240
rect 0 195576 800 195696
rect 0 195168 800 195288
rect 0 194624 800 194744
rect 69200 194760 70000 194880
rect 0 194080 800 194200
rect 0 193672 800 193792
rect 0 193128 800 193248
rect 0 192584 800 192704
rect 69200 192720 70000 192840
rect 0 192176 800 192296
rect 0 191632 800 191752
rect 0 191088 800 191208
rect 0 190680 800 190800
rect 69200 190680 70000 190800
rect 0 190136 800 190256
rect 0 189592 800 189712
rect 0 189184 800 189304
rect 0 188640 800 188760
rect 69200 188640 70000 188760
rect 0 188096 800 188216
rect 0 187688 800 187808
rect 0 187144 800 187264
rect 0 186600 800 186720
rect 69200 186600 70000 186720
rect 0 186192 800 186312
rect 0 185648 800 185768
rect 0 185104 800 185224
rect 0 184560 800 184680
rect 69200 184560 70000 184680
rect 0 184152 800 184272
rect 0 183608 800 183728
rect 0 183064 800 183184
rect 0 182656 800 182776
rect 69200 182520 70000 182640
rect 0 182112 800 182232
rect 0 181568 800 181688
rect 0 181160 800 181280
rect 0 180616 800 180736
rect 69200 180480 70000 180600
rect 0 180072 800 180192
rect 0 179664 800 179784
rect 0 179120 800 179240
rect 0 178576 800 178696
rect 69200 178440 70000 178560
rect 0 178168 800 178288
rect 0 177624 800 177744
rect 0 177080 800 177200
rect 0 176672 800 176792
rect 69200 176400 70000 176520
rect 0 176128 800 176248
rect 0 175584 800 175704
rect 0 175176 800 175296
rect 0 174632 800 174752
rect 69200 174360 70000 174480
rect 0 174088 800 174208
rect 0 173680 800 173800
rect 0 173136 800 173256
rect 0 172592 800 172712
rect 0 172184 800 172304
rect 69200 172320 70000 172440
rect 0 171640 800 171760
rect 0 171096 800 171216
rect 0 170688 800 170808
rect 0 170144 800 170264
rect 69200 170280 70000 170400
rect 0 169600 800 169720
rect 0 169056 800 169176
rect 0 168648 800 168768
rect 0 168104 800 168224
rect 69200 168240 70000 168360
rect 0 167560 800 167680
rect 0 167152 800 167272
rect 0 166608 800 166728
rect 0 166064 800 166184
rect 69200 166200 70000 166320
rect 0 165656 800 165776
rect 0 165112 800 165232
rect 0 164568 800 164688
rect 0 164160 800 164280
rect 69200 164160 70000 164280
rect 0 163616 800 163736
rect 0 163072 800 163192
rect 0 162664 800 162784
rect 0 162120 800 162240
rect 69200 162120 70000 162240
rect 0 161576 800 161696
rect 0 161168 800 161288
rect 0 160624 800 160744
rect 0 160080 800 160200
rect 69200 160080 70000 160200
rect 0 159672 800 159792
rect 0 159128 800 159248
rect 0 158584 800 158704
rect 0 158176 800 158296
rect 69200 158040 70000 158160
rect 0 157632 800 157752
rect 0 157088 800 157208
rect 0 156680 800 156800
rect 0 156136 800 156256
rect 69200 156000 70000 156120
rect 0 155592 800 155712
rect 0 155184 800 155304
rect 0 154640 800 154760
rect 0 154096 800 154216
rect 69200 153960 70000 154080
rect 0 153552 800 153672
rect 0 153144 800 153264
rect 0 152600 800 152720
rect 0 152056 800 152176
rect 69200 151920 70000 152040
rect 0 151648 800 151768
rect 0 151104 800 151224
rect 0 150560 800 150680
rect 0 150152 800 150272
rect 69200 149880 70000 150000
rect 0 149608 800 149728
rect 0 149064 800 149184
rect 0 148656 800 148776
rect 0 148112 800 148232
rect 69200 147840 70000 147960
rect 0 147568 800 147688
rect 0 147160 800 147280
rect 0 146616 800 146736
rect 0 146072 800 146192
rect 0 145664 800 145784
rect 69200 145800 70000 145920
rect 0 145120 800 145240
rect 0 144576 800 144696
rect 0 144168 800 144288
rect 0 143624 800 143744
rect 69200 143760 70000 143880
rect 0 143080 800 143200
rect 0 142672 800 142792
rect 0 142128 800 142248
rect 0 141584 800 141704
rect 69200 141720 70000 141840
rect 0 141176 800 141296
rect 0 140632 800 140752
rect 0 140088 800 140208
rect 0 139680 800 139800
rect 69200 139680 70000 139800
rect 0 139136 800 139256
rect 0 138592 800 138712
rect 0 138048 800 138168
rect 0 137640 800 137760
rect 69200 137640 70000 137760
rect 0 137096 800 137216
rect 0 136552 800 136672
rect 0 136144 800 136264
rect 0 135600 800 135720
rect 69200 135600 70000 135720
rect 0 135056 800 135176
rect 0 134648 800 134768
rect 0 134104 800 134224
rect 0 133560 800 133680
rect 69200 133560 70000 133680
rect 0 133152 800 133272
rect 0 132608 800 132728
rect 0 132064 800 132184
rect 0 131656 800 131776
rect 69200 131520 70000 131640
rect 0 131112 800 131232
rect 0 130568 800 130688
rect 0 130160 800 130280
rect 0 129616 800 129736
rect 69200 129480 70000 129600
rect 0 129072 800 129192
rect 0 128664 800 128784
rect 0 128120 800 128240
rect 0 127576 800 127696
rect 69200 127440 70000 127560
rect 0 127168 800 127288
rect 0 126624 800 126744
rect 0 126080 800 126200
rect 0 125672 800 125792
rect 69200 125400 70000 125520
rect 0 125128 800 125248
rect 0 124584 800 124704
rect 0 124176 800 124296
rect 0 123632 800 123752
rect 69200 123360 70000 123480
rect 0 123088 800 123208
rect 0 122544 800 122664
rect 0 122136 800 122256
rect 0 121592 800 121712
rect 69200 121320 70000 121440
rect 0 121048 800 121168
rect 0 120640 800 120760
rect 0 120096 800 120216
rect 0 119552 800 119672
rect 0 119144 800 119264
rect 69200 119280 70000 119400
rect 0 118600 800 118720
rect 0 118056 800 118176
rect 0 117648 800 117768
rect 0 117104 800 117224
rect 69200 117240 70000 117360
rect 0 116560 800 116680
rect 0 116152 800 116272
rect 0 115608 800 115728
rect 0 115064 800 115184
rect 69200 115200 70000 115320
rect 0 114656 800 114776
rect 0 114112 800 114232
rect 0 113568 800 113688
rect 0 113160 800 113280
rect 69200 113160 70000 113280
rect 0 112616 800 112736
rect 0 112072 800 112192
rect 0 111664 800 111784
rect 0 111120 800 111240
rect 69200 111120 70000 111240
rect 0 110576 800 110696
rect 0 110168 800 110288
rect 0 109624 800 109744
rect 0 109080 800 109200
rect 69200 109080 70000 109200
rect 0 108672 800 108792
rect 0 108128 800 108248
rect 0 107584 800 107704
rect 0 107040 800 107160
rect 69200 107040 70000 107160
rect 0 106632 800 106752
rect 0 106088 800 106208
rect 0 105544 800 105664
rect 0 105136 800 105256
rect 69200 105000 70000 105120
rect 0 104592 800 104712
rect 0 104048 800 104168
rect 0 103640 800 103760
rect 0 103096 800 103216
rect 69200 102960 70000 103080
rect 0 102552 800 102672
rect 0 102144 800 102264
rect 0 101600 800 101720
rect 0 101056 800 101176
rect 69200 100920 70000 101040
rect 0 100648 800 100768
rect 0 100104 800 100224
rect 0 99560 800 99680
rect 0 99152 800 99272
rect 69200 98880 70000 99000
rect 0 98608 800 98728
rect 0 98064 800 98184
rect 0 97656 800 97776
rect 0 97112 800 97232
rect 69200 96840 70000 96960
rect 0 96568 800 96688
rect 0 96160 800 96280
rect 0 95616 800 95736
rect 0 95072 800 95192
rect 0 94664 800 94784
rect 69200 94800 70000 94920
rect 0 94120 800 94240
rect 0 93576 800 93696
rect 0 93168 800 93288
rect 0 92624 800 92744
rect 69200 92760 70000 92880
rect 0 92080 800 92200
rect 0 91536 800 91656
rect 0 91128 800 91248
rect 0 90584 800 90704
rect 69200 90720 70000 90840
rect 0 90040 800 90160
rect 0 89632 800 89752
rect 0 89088 800 89208
rect 0 88544 800 88664
rect 69200 88680 70000 88800
rect 0 88136 800 88256
rect 0 87592 800 87712
rect 0 87048 800 87168
rect 0 86640 800 86760
rect 69200 86640 70000 86760
rect 0 86096 800 86216
rect 0 85552 800 85672
rect 0 85144 800 85264
rect 0 84600 800 84720
rect 69200 84600 70000 84720
rect 0 84056 800 84176
rect 0 83648 800 83768
rect 0 83104 800 83224
rect 0 82560 800 82680
rect 69200 82560 70000 82680
rect 0 82152 800 82272
rect 0 81608 800 81728
rect 0 81064 800 81184
rect 0 80656 800 80776
rect 69200 80520 70000 80640
rect 0 80112 800 80232
rect 0 79568 800 79688
rect 0 79160 800 79280
rect 0 78616 800 78736
rect 69200 78480 70000 78600
rect 0 78072 800 78192
rect 0 77664 800 77784
rect 0 77120 800 77240
rect 0 76576 800 76696
rect 69200 76440 70000 76560
rect 0 76032 800 76152
rect 0 75624 800 75744
rect 0 75080 800 75200
rect 0 74536 800 74656
rect 69200 74400 70000 74520
rect 0 74128 800 74248
rect 0 73584 800 73704
rect 0 73040 800 73160
rect 0 72632 800 72752
rect 69200 72360 70000 72480
rect 0 72088 800 72208
rect 0 71544 800 71664
rect 0 71136 800 71256
rect 0 70592 800 70712
rect 69200 70320 70000 70440
rect 0 70048 800 70168
rect 0 69640 800 69760
rect 0 69096 800 69216
rect 0 68552 800 68672
rect 0 68144 800 68264
rect 69200 68280 70000 68400
rect 0 67600 800 67720
rect 0 67056 800 67176
rect 0 66648 800 66768
rect 0 66104 800 66224
rect 69200 66240 70000 66360
rect 0 65560 800 65680
rect 0 65152 800 65272
rect 0 64608 800 64728
rect 0 64064 800 64184
rect 69200 64200 70000 64320
rect 0 63656 800 63776
rect 0 63112 800 63232
rect 0 62568 800 62688
rect 0 62160 800 62280
rect 69200 62160 70000 62280
rect 0 61616 800 61736
rect 0 61072 800 61192
rect 0 60528 800 60648
rect 0 60120 800 60240
rect 69200 60120 70000 60240
rect 0 59576 800 59696
rect 0 59032 800 59152
rect 0 58624 800 58744
rect 0 58080 800 58200
rect 69200 58080 70000 58200
rect 0 57536 800 57656
rect 0 57128 800 57248
rect 0 56584 800 56704
rect 0 56040 800 56160
rect 69200 56040 70000 56160
rect 0 55632 800 55752
rect 0 55088 800 55208
rect 0 54544 800 54664
rect 0 54136 800 54256
rect 69200 54000 70000 54120
rect 0 53592 800 53712
rect 0 53048 800 53168
rect 0 52640 800 52760
rect 0 52096 800 52216
rect 69200 51960 70000 52080
rect 0 51552 800 51672
rect 0 51144 800 51264
rect 0 50600 800 50720
rect 0 50056 800 50176
rect 69200 49920 70000 50040
rect 0 49648 800 49768
rect 0 49104 800 49224
rect 0 48560 800 48680
rect 0 48152 800 48272
rect 69200 47880 70000 48000
rect 0 47608 800 47728
rect 0 47064 800 47184
rect 0 46656 800 46776
rect 0 46112 800 46232
rect 69200 45840 70000 45960
rect 0 45568 800 45688
rect 0 45024 800 45144
rect 0 44616 800 44736
rect 0 44072 800 44192
rect 69200 43800 70000 43920
rect 0 43528 800 43648
rect 0 43120 800 43240
rect 0 42576 800 42696
rect 0 42032 800 42152
rect 0 41624 800 41744
rect 69200 41760 70000 41880
rect 0 41080 800 41200
rect 0 40536 800 40656
rect 0 40128 800 40248
rect 0 39584 800 39704
rect 69200 39720 70000 39840
rect 0 39040 800 39160
rect 0 38632 800 38752
rect 0 38088 800 38208
rect 0 37544 800 37664
rect 69200 37680 70000 37800
rect 0 37136 800 37256
rect 0 36592 800 36712
rect 0 36048 800 36168
rect 0 35640 800 35760
rect 69200 35640 70000 35760
rect 0 35096 800 35216
rect 0 34552 800 34672
rect 0 34144 800 34264
rect 0 33600 800 33720
rect 69200 33600 70000 33720
rect 0 33056 800 33176
rect 0 32648 800 32768
rect 0 32104 800 32224
rect 0 31560 800 31680
rect 69200 31560 70000 31680
rect 0 31152 800 31272
rect 0 30608 800 30728
rect 0 30064 800 30184
rect 0 29520 800 29640
rect 69200 29520 70000 29640
rect 0 29112 800 29232
rect 0 28568 800 28688
rect 0 28024 800 28144
rect 0 27616 800 27736
rect 69200 27480 70000 27600
rect 0 27072 800 27192
rect 0 26528 800 26648
rect 0 26120 800 26240
rect 0 25576 800 25696
rect 69200 25440 70000 25560
rect 0 25032 800 25152
rect 0 24624 800 24744
rect 0 24080 800 24200
rect 0 23536 800 23656
rect 69200 23400 70000 23520
rect 0 23128 800 23248
rect 0 22584 800 22704
rect 0 22040 800 22160
rect 0 21632 800 21752
rect 69200 21360 70000 21480
rect 0 21088 800 21208
rect 0 20544 800 20664
rect 0 20136 800 20256
rect 0 19592 800 19712
rect 69200 19320 70000 19440
rect 0 19048 800 19168
rect 0 18640 800 18760
rect 0 18096 800 18216
rect 0 17552 800 17672
rect 0 17144 800 17264
rect 69200 17280 70000 17400
rect 0 16600 800 16720
rect 0 16056 800 16176
rect 0 15648 800 15768
rect 0 15104 800 15224
rect 69200 15240 70000 15360
rect 0 14560 800 14680
rect 0 14016 800 14136
rect 0 13608 800 13728
rect 0 13064 800 13184
rect 69200 13200 70000 13320
rect 0 12520 800 12640
rect 0 12112 800 12232
rect 0 11568 800 11688
rect 0 11024 800 11144
rect 69200 11160 70000 11280
rect 0 10616 800 10736
rect 0 10072 800 10192
rect 0 9528 800 9648
rect 0 9120 800 9240
rect 69200 9120 70000 9240
rect 0 8576 800 8696
rect 0 8032 800 8152
rect 0 7624 800 7744
rect 0 7080 800 7200
rect 69200 7080 70000 7200
rect 0 6536 800 6656
rect 0 6128 800 6248
rect 0 5584 800 5704
rect 0 5040 800 5160
rect 69200 5040 70000 5160
rect 0 4632 800 4752
rect 0 4088 800 4208
rect 0 3544 800 3664
rect 0 3136 800 3256
rect 69200 3000 70000 3120
rect 0 2592 800 2712
rect 0 2048 800 2168
rect 0 1640 800 1760
rect 0 1096 800 1216
rect 69200 960 70000 1080
rect 0 552 800 672
rect 0 144 800 264
<< obsm3 >>
rect 880 199576 69200 199749
rect 381 199312 69200 199576
rect 880 199040 69200 199312
rect 880 199032 69120 199040
rect 381 198768 69120 199032
rect 880 198760 69120 198768
rect 880 198488 69200 198760
rect 381 198360 69200 198488
rect 880 198080 69200 198360
rect 381 197816 69200 198080
rect 880 197536 69200 197816
rect 381 197272 69200 197536
rect 880 197000 69200 197272
rect 880 196992 69120 197000
rect 381 196864 69120 196992
rect 880 196720 69120 196864
rect 880 196584 69200 196720
rect 381 196320 69200 196584
rect 880 196040 69200 196320
rect 381 195776 69200 196040
rect 880 195496 69200 195776
rect 381 195368 69200 195496
rect 880 195088 69200 195368
rect 381 194960 69200 195088
rect 381 194824 69120 194960
rect 880 194680 69120 194824
rect 880 194544 69200 194680
rect 381 194280 69200 194544
rect 880 194000 69200 194280
rect 381 193872 69200 194000
rect 880 193592 69200 193872
rect 381 193328 69200 193592
rect 880 193048 69200 193328
rect 381 192920 69200 193048
rect 381 192784 69120 192920
rect 880 192640 69120 192784
rect 880 192504 69200 192640
rect 381 192376 69200 192504
rect 880 192096 69200 192376
rect 381 191832 69200 192096
rect 880 191552 69200 191832
rect 381 191288 69200 191552
rect 880 191008 69200 191288
rect 381 190880 69200 191008
rect 880 190600 69120 190880
rect 381 190336 69200 190600
rect 880 190056 69200 190336
rect 381 189792 69200 190056
rect 880 189512 69200 189792
rect 381 189384 69200 189512
rect 880 189104 69200 189384
rect 381 188840 69200 189104
rect 880 188560 69120 188840
rect 381 188296 69200 188560
rect 880 188016 69200 188296
rect 381 187888 69200 188016
rect 880 187608 69200 187888
rect 381 187344 69200 187608
rect 880 187064 69200 187344
rect 381 186800 69200 187064
rect 880 186520 69120 186800
rect 381 186392 69200 186520
rect 880 186112 69200 186392
rect 381 185848 69200 186112
rect 880 185568 69200 185848
rect 381 185304 69200 185568
rect 880 185024 69200 185304
rect 381 184760 69200 185024
rect 880 184480 69120 184760
rect 381 184352 69200 184480
rect 880 184072 69200 184352
rect 381 183808 69200 184072
rect 880 183528 69200 183808
rect 381 183264 69200 183528
rect 880 182984 69200 183264
rect 381 182856 69200 182984
rect 880 182720 69200 182856
rect 880 182576 69120 182720
rect 381 182440 69120 182576
rect 381 182312 69200 182440
rect 880 182032 69200 182312
rect 381 181768 69200 182032
rect 880 181488 69200 181768
rect 381 181360 69200 181488
rect 880 181080 69200 181360
rect 381 180816 69200 181080
rect 880 180680 69200 180816
rect 880 180536 69120 180680
rect 381 180400 69120 180536
rect 381 180272 69200 180400
rect 880 179992 69200 180272
rect 381 179864 69200 179992
rect 880 179584 69200 179864
rect 381 179320 69200 179584
rect 880 179040 69200 179320
rect 381 178776 69200 179040
rect 880 178640 69200 178776
rect 880 178496 69120 178640
rect 381 178368 69120 178496
rect 880 178360 69120 178368
rect 880 178088 69200 178360
rect 381 177824 69200 178088
rect 880 177544 69200 177824
rect 381 177280 69200 177544
rect 880 177000 69200 177280
rect 381 176872 69200 177000
rect 880 176600 69200 176872
rect 880 176592 69120 176600
rect 381 176328 69120 176592
rect 880 176320 69120 176328
rect 880 176048 69200 176320
rect 381 175784 69200 176048
rect 880 175504 69200 175784
rect 381 175376 69200 175504
rect 880 175096 69200 175376
rect 381 174832 69200 175096
rect 880 174560 69200 174832
rect 880 174552 69120 174560
rect 381 174288 69120 174552
rect 880 174280 69120 174288
rect 880 174008 69200 174280
rect 381 173880 69200 174008
rect 880 173600 69200 173880
rect 381 173336 69200 173600
rect 880 173056 69200 173336
rect 381 172792 69200 173056
rect 880 172520 69200 172792
rect 880 172512 69120 172520
rect 381 172384 69120 172512
rect 880 172240 69120 172384
rect 880 172104 69200 172240
rect 381 171840 69200 172104
rect 880 171560 69200 171840
rect 381 171296 69200 171560
rect 880 171016 69200 171296
rect 381 170888 69200 171016
rect 880 170608 69200 170888
rect 381 170480 69200 170608
rect 381 170344 69120 170480
rect 880 170200 69120 170344
rect 880 170064 69200 170200
rect 381 169800 69200 170064
rect 880 169520 69200 169800
rect 381 169256 69200 169520
rect 880 168976 69200 169256
rect 381 168848 69200 168976
rect 880 168568 69200 168848
rect 381 168440 69200 168568
rect 381 168304 69120 168440
rect 880 168160 69120 168304
rect 880 168024 69200 168160
rect 381 167760 69200 168024
rect 880 167480 69200 167760
rect 381 167352 69200 167480
rect 880 167072 69200 167352
rect 381 166808 69200 167072
rect 880 166528 69200 166808
rect 381 166400 69200 166528
rect 381 166264 69120 166400
rect 880 166120 69120 166264
rect 880 165984 69200 166120
rect 381 165856 69200 165984
rect 880 165576 69200 165856
rect 381 165312 69200 165576
rect 880 165032 69200 165312
rect 381 164768 69200 165032
rect 880 164488 69200 164768
rect 381 164360 69200 164488
rect 880 164080 69120 164360
rect 381 163816 69200 164080
rect 880 163536 69200 163816
rect 381 163272 69200 163536
rect 880 162992 69200 163272
rect 381 162864 69200 162992
rect 880 162584 69200 162864
rect 381 162320 69200 162584
rect 880 162040 69120 162320
rect 381 161776 69200 162040
rect 880 161496 69200 161776
rect 381 161368 69200 161496
rect 880 161088 69200 161368
rect 381 160824 69200 161088
rect 880 160544 69200 160824
rect 381 160280 69200 160544
rect 880 160000 69120 160280
rect 381 159872 69200 160000
rect 880 159592 69200 159872
rect 381 159328 69200 159592
rect 880 159048 69200 159328
rect 381 158784 69200 159048
rect 880 158504 69200 158784
rect 381 158376 69200 158504
rect 880 158240 69200 158376
rect 880 158096 69120 158240
rect 381 157960 69120 158096
rect 381 157832 69200 157960
rect 880 157552 69200 157832
rect 381 157288 69200 157552
rect 880 157008 69200 157288
rect 381 156880 69200 157008
rect 880 156600 69200 156880
rect 381 156336 69200 156600
rect 880 156200 69200 156336
rect 880 156056 69120 156200
rect 381 155920 69120 156056
rect 381 155792 69200 155920
rect 880 155512 69200 155792
rect 381 155384 69200 155512
rect 880 155104 69200 155384
rect 381 154840 69200 155104
rect 880 154560 69200 154840
rect 381 154296 69200 154560
rect 880 154160 69200 154296
rect 880 154016 69120 154160
rect 381 153880 69120 154016
rect 381 153752 69200 153880
rect 880 153472 69200 153752
rect 381 153344 69200 153472
rect 880 153064 69200 153344
rect 381 152800 69200 153064
rect 880 152520 69200 152800
rect 381 152256 69200 152520
rect 880 152120 69200 152256
rect 880 151976 69120 152120
rect 381 151848 69120 151976
rect 880 151840 69120 151848
rect 880 151568 69200 151840
rect 381 151304 69200 151568
rect 880 151024 69200 151304
rect 381 150760 69200 151024
rect 880 150480 69200 150760
rect 381 150352 69200 150480
rect 880 150080 69200 150352
rect 880 150072 69120 150080
rect 381 149808 69120 150072
rect 880 149800 69120 149808
rect 880 149528 69200 149800
rect 381 149264 69200 149528
rect 880 148984 69200 149264
rect 381 148856 69200 148984
rect 880 148576 69200 148856
rect 381 148312 69200 148576
rect 880 148040 69200 148312
rect 880 148032 69120 148040
rect 381 147768 69120 148032
rect 880 147760 69120 147768
rect 880 147488 69200 147760
rect 381 147360 69200 147488
rect 880 147080 69200 147360
rect 381 146816 69200 147080
rect 880 146536 69200 146816
rect 381 146272 69200 146536
rect 880 146000 69200 146272
rect 880 145992 69120 146000
rect 381 145864 69120 145992
rect 880 145720 69120 145864
rect 880 145584 69200 145720
rect 381 145320 69200 145584
rect 880 145040 69200 145320
rect 381 144776 69200 145040
rect 880 144496 69200 144776
rect 381 144368 69200 144496
rect 880 144088 69200 144368
rect 381 143960 69200 144088
rect 381 143824 69120 143960
rect 880 143680 69120 143824
rect 880 143544 69200 143680
rect 381 143280 69200 143544
rect 880 143000 69200 143280
rect 381 142872 69200 143000
rect 880 142592 69200 142872
rect 381 142328 69200 142592
rect 880 142048 69200 142328
rect 381 141920 69200 142048
rect 381 141784 69120 141920
rect 880 141640 69120 141784
rect 880 141504 69200 141640
rect 381 141376 69200 141504
rect 880 141096 69200 141376
rect 381 140832 69200 141096
rect 880 140552 69200 140832
rect 381 140288 69200 140552
rect 880 140008 69200 140288
rect 381 139880 69200 140008
rect 880 139600 69120 139880
rect 381 139336 69200 139600
rect 880 139056 69200 139336
rect 381 138792 69200 139056
rect 880 138512 69200 138792
rect 381 138248 69200 138512
rect 880 137968 69200 138248
rect 381 137840 69200 137968
rect 880 137560 69120 137840
rect 381 137296 69200 137560
rect 880 137016 69200 137296
rect 381 136752 69200 137016
rect 880 136472 69200 136752
rect 381 136344 69200 136472
rect 880 136064 69200 136344
rect 381 135800 69200 136064
rect 880 135520 69120 135800
rect 381 135256 69200 135520
rect 880 134976 69200 135256
rect 381 134848 69200 134976
rect 880 134568 69200 134848
rect 381 134304 69200 134568
rect 880 134024 69200 134304
rect 381 133760 69200 134024
rect 880 133480 69120 133760
rect 381 133352 69200 133480
rect 880 133072 69200 133352
rect 381 132808 69200 133072
rect 880 132528 69200 132808
rect 381 132264 69200 132528
rect 880 131984 69200 132264
rect 381 131856 69200 131984
rect 880 131720 69200 131856
rect 880 131576 69120 131720
rect 381 131440 69120 131576
rect 381 131312 69200 131440
rect 880 131032 69200 131312
rect 381 130768 69200 131032
rect 880 130488 69200 130768
rect 381 130360 69200 130488
rect 880 130080 69200 130360
rect 381 129816 69200 130080
rect 880 129680 69200 129816
rect 880 129536 69120 129680
rect 381 129400 69120 129536
rect 381 129272 69200 129400
rect 880 128992 69200 129272
rect 381 128864 69200 128992
rect 880 128584 69200 128864
rect 381 128320 69200 128584
rect 880 128040 69200 128320
rect 381 127776 69200 128040
rect 880 127640 69200 127776
rect 880 127496 69120 127640
rect 381 127368 69120 127496
rect 880 127360 69120 127368
rect 880 127088 69200 127360
rect 381 126824 69200 127088
rect 880 126544 69200 126824
rect 381 126280 69200 126544
rect 880 126000 69200 126280
rect 381 125872 69200 126000
rect 880 125600 69200 125872
rect 880 125592 69120 125600
rect 381 125328 69120 125592
rect 880 125320 69120 125328
rect 880 125048 69200 125320
rect 381 124784 69200 125048
rect 880 124504 69200 124784
rect 381 124376 69200 124504
rect 880 124096 69200 124376
rect 381 123832 69200 124096
rect 880 123560 69200 123832
rect 880 123552 69120 123560
rect 381 123288 69120 123552
rect 880 123280 69120 123288
rect 880 123008 69200 123280
rect 381 122744 69200 123008
rect 880 122464 69200 122744
rect 381 122336 69200 122464
rect 880 122056 69200 122336
rect 381 121792 69200 122056
rect 880 121520 69200 121792
rect 880 121512 69120 121520
rect 381 121248 69120 121512
rect 880 121240 69120 121248
rect 880 120968 69200 121240
rect 381 120840 69200 120968
rect 880 120560 69200 120840
rect 381 120296 69200 120560
rect 880 120016 69200 120296
rect 381 119752 69200 120016
rect 880 119480 69200 119752
rect 880 119472 69120 119480
rect 381 119344 69120 119472
rect 880 119200 69120 119344
rect 880 119064 69200 119200
rect 381 118800 69200 119064
rect 880 118520 69200 118800
rect 381 118256 69200 118520
rect 880 117976 69200 118256
rect 381 117848 69200 117976
rect 880 117568 69200 117848
rect 381 117440 69200 117568
rect 381 117304 69120 117440
rect 880 117160 69120 117304
rect 880 117024 69200 117160
rect 381 116760 69200 117024
rect 880 116480 69200 116760
rect 381 116352 69200 116480
rect 880 116072 69200 116352
rect 381 115808 69200 116072
rect 880 115528 69200 115808
rect 381 115400 69200 115528
rect 381 115264 69120 115400
rect 880 115120 69120 115264
rect 880 114984 69200 115120
rect 381 114856 69200 114984
rect 880 114576 69200 114856
rect 381 114312 69200 114576
rect 880 114032 69200 114312
rect 381 113768 69200 114032
rect 880 113488 69200 113768
rect 381 113360 69200 113488
rect 880 113080 69120 113360
rect 381 112816 69200 113080
rect 880 112536 69200 112816
rect 381 112272 69200 112536
rect 880 111992 69200 112272
rect 381 111864 69200 111992
rect 880 111584 69200 111864
rect 381 111320 69200 111584
rect 880 111040 69120 111320
rect 381 110776 69200 111040
rect 880 110496 69200 110776
rect 381 110368 69200 110496
rect 880 110088 69200 110368
rect 381 109824 69200 110088
rect 880 109544 69200 109824
rect 381 109280 69200 109544
rect 880 109000 69120 109280
rect 381 108872 69200 109000
rect 880 108592 69200 108872
rect 381 108328 69200 108592
rect 880 108048 69200 108328
rect 381 107784 69200 108048
rect 880 107504 69200 107784
rect 381 107240 69200 107504
rect 880 106960 69120 107240
rect 381 106832 69200 106960
rect 880 106552 69200 106832
rect 381 106288 69200 106552
rect 880 106008 69200 106288
rect 381 105744 69200 106008
rect 880 105464 69200 105744
rect 381 105336 69200 105464
rect 880 105200 69200 105336
rect 880 105056 69120 105200
rect 381 104920 69120 105056
rect 381 104792 69200 104920
rect 880 104512 69200 104792
rect 381 104248 69200 104512
rect 880 103968 69200 104248
rect 381 103840 69200 103968
rect 880 103560 69200 103840
rect 381 103296 69200 103560
rect 880 103160 69200 103296
rect 880 103016 69120 103160
rect 381 102880 69120 103016
rect 381 102752 69200 102880
rect 880 102472 69200 102752
rect 381 102344 69200 102472
rect 880 102064 69200 102344
rect 381 101800 69200 102064
rect 880 101520 69200 101800
rect 381 101256 69200 101520
rect 880 101120 69200 101256
rect 880 100976 69120 101120
rect 381 100848 69120 100976
rect 880 100840 69120 100848
rect 880 100568 69200 100840
rect 381 100304 69200 100568
rect 880 100024 69200 100304
rect 381 99760 69200 100024
rect 880 99480 69200 99760
rect 381 99352 69200 99480
rect 880 99080 69200 99352
rect 880 99072 69120 99080
rect 381 98808 69120 99072
rect 880 98800 69120 98808
rect 880 98528 69200 98800
rect 381 98264 69200 98528
rect 880 97984 69200 98264
rect 381 97856 69200 97984
rect 880 97576 69200 97856
rect 381 97312 69200 97576
rect 880 97040 69200 97312
rect 880 97032 69120 97040
rect 381 96768 69120 97032
rect 880 96760 69120 96768
rect 880 96488 69200 96760
rect 381 96360 69200 96488
rect 880 96080 69200 96360
rect 381 95816 69200 96080
rect 880 95536 69200 95816
rect 381 95272 69200 95536
rect 880 95000 69200 95272
rect 880 94992 69120 95000
rect 381 94864 69120 94992
rect 880 94720 69120 94864
rect 880 94584 69200 94720
rect 381 94320 69200 94584
rect 880 94040 69200 94320
rect 381 93776 69200 94040
rect 880 93496 69200 93776
rect 381 93368 69200 93496
rect 880 93088 69200 93368
rect 381 92960 69200 93088
rect 381 92824 69120 92960
rect 880 92680 69120 92824
rect 880 92544 69200 92680
rect 381 92280 69200 92544
rect 880 92000 69200 92280
rect 381 91736 69200 92000
rect 880 91456 69200 91736
rect 381 91328 69200 91456
rect 880 91048 69200 91328
rect 381 90920 69200 91048
rect 381 90784 69120 90920
rect 880 90640 69120 90784
rect 880 90504 69200 90640
rect 381 90240 69200 90504
rect 880 89960 69200 90240
rect 381 89832 69200 89960
rect 880 89552 69200 89832
rect 381 89288 69200 89552
rect 880 89008 69200 89288
rect 381 88880 69200 89008
rect 381 88744 69120 88880
rect 880 88600 69120 88744
rect 880 88464 69200 88600
rect 381 88336 69200 88464
rect 880 88056 69200 88336
rect 381 87792 69200 88056
rect 880 87512 69200 87792
rect 381 87248 69200 87512
rect 880 86968 69200 87248
rect 381 86840 69200 86968
rect 880 86560 69120 86840
rect 381 86296 69200 86560
rect 880 86016 69200 86296
rect 381 85752 69200 86016
rect 880 85472 69200 85752
rect 381 85344 69200 85472
rect 880 85064 69200 85344
rect 381 84800 69200 85064
rect 880 84520 69120 84800
rect 381 84256 69200 84520
rect 880 83976 69200 84256
rect 381 83848 69200 83976
rect 880 83568 69200 83848
rect 381 83304 69200 83568
rect 880 83024 69200 83304
rect 381 82760 69200 83024
rect 880 82480 69120 82760
rect 381 82352 69200 82480
rect 880 82072 69200 82352
rect 381 81808 69200 82072
rect 880 81528 69200 81808
rect 381 81264 69200 81528
rect 880 80984 69200 81264
rect 381 80856 69200 80984
rect 880 80720 69200 80856
rect 880 80576 69120 80720
rect 381 80440 69120 80576
rect 381 80312 69200 80440
rect 880 80032 69200 80312
rect 381 79768 69200 80032
rect 880 79488 69200 79768
rect 381 79360 69200 79488
rect 880 79080 69200 79360
rect 381 78816 69200 79080
rect 880 78680 69200 78816
rect 880 78536 69120 78680
rect 381 78400 69120 78536
rect 381 78272 69200 78400
rect 880 77992 69200 78272
rect 381 77864 69200 77992
rect 880 77584 69200 77864
rect 381 77320 69200 77584
rect 880 77040 69200 77320
rect 381 76776 69200 77040
rect 880 76640 69200 76776
rect 880 76496 69120 76640
rect 381 76360 69120 76496
rect 381 76232 69200 76360
rect 880 75952 69200 76232
rect 381 75824 69200 75952
rect 880 75544 69200 75824
rect 381 75280 69200 75544
rect 880 75000 69200 75280
rect 381 74736 69200 75000
rect 880 74600 69200 74736
rect 880 74456 69120 74600
rect 381 74328 69120 74456
rect 880 74320 69120 74328
rect 880 74048 69200 74320
rect 381 73784 69200 74048
rect 880 73504 69200 73784
rect 381 73240 69200 73504
rect 880 72960 69200 73240
rect 381 72832 69200 72960
rect 880 72560 69200 72832
rect 880 72552 69120 72560
rect 381 72288 69120 72552
rect 880 72280 69120 72288
rect 880 72008 69200 72280
rect 381 71744 69200 72008
rect 880 71464 69200 71744
rect 381 71336 69200 71464
rect 880 71056 69200 71336
rect 381 70792 69200 71056
rect 880 70520 69200 70792
rect 880 70512 69120 70520
rect 381 70248 69120 70512
rect 880 70240 69120 70248
rect 880 69968 69200 70240
rect 381 69840 69200 69968
rect 880 69560 69200 69840
rect 381 69296 69200 69560
rect 880 69016 69200 69296
rect 381 68752 69200 69016
rect 880 68480 69200 68752
rect 880 68472 69120 68480
rect 381 68344 69120 68472
rect 880 68200 69120 68344
rect 880 68064 69200 68200
rect 381 67800 69200 68064
rect 880 67520 69200 67800
rect 381 67256 69200 67520
rect 880 66976 69200 67256
rect 381 66848 69200 66976
rect 880 66568 69200 66848
rect 381 66440 69200 66568
rect 381 66304 69120 66440
rect 880 66160 69120 66304
rect 880 66024 69200 66160
rect 381 65760 69200 66024
rect 880 65480 69200 65760
rect 381 65352 69200 65480
rect 880 65072 69200 65352
rect 381 64808 69200 65072
rect 880 64528 69200 64808
rect 381 64400 69200 64528
rect 381 64264 69120 64400
rect 880 64120 69120 64264
rect 880 63984 69200 64120
rect 381 63856 69200 63984
rect 880 63576 69200 63856
rect 381 63312 69200 63576
rect 880 63032 69200 63312
rect 381 62768 69200 63032
rect 880 62488 69200 62768
rect 381 62360 69200 62488
rect 880 62080 69120 62360
rect 381 61816 69200 62080
rect 880 61536 69200 61816
rect 381 61272 69200 61536
rect 880 60992 69200 61272
rect 381 60728 69200 60992
rect 880 60448 69200 60728
rect 381 60320 69200 60448
rect 880 60040 69120 60320
rect 381 59776 69200 60040
rect 880 59496 69200 59776
rect 381 59232 69200 59496
rect 880 58952 69200 59232
rect 381 58824 69200 58952
rect 880 58544 69200 58824
rect 381 58280 69200 58544
rect 880 58000 69120 58280
rect 381 57736 69200 58000
rect 880 57456 69200 57736
rect 381 57328 69200 57456
rect 880 57048 69200 57328
rect 381 56784 69200 57048
rect 880 56504 69200 56784
rect 381 56240 69200 56504
rect 880 55960 69120 56240
rect 381 55832 69200 55960
rect 880 55552 69200 55832
rect 381 55288 69200 55552
rect 880 55008 69200 55288
rect 381 54744 69200 55008
rect 880 54464 69200 54744
rect 381 54336 69200 54464
rect 880 54200 69200 54336
rect 880 54056 69120 54200
rect 381 53920 69120 54056
rect 381 53792 69200 53920
rect 880 53512 69200 53792
rect 381 53248 69200 53512
rect 880 52968 69200 53248
rect 381 52840 69200 52968
rect 880 52560 69200 52840
rect 381 52296 69200 52560
rect 880 52160 69200 52296
rect 880 52016 69120 52160
rect 381 51880 69120 52016
rect 381 51752 69200 51880
rect 880 51472 69200 51752
rect 381 51344 69200 51472
rect 880 51064 69200 51344
rect 381 50800 69200 51064
rect 880 50520 69200 50800
rect 381 50256 69200 50520
rect 880 50120 69200 50256
rect 880 49976 69120 50120
rect 381 49848 69120 49976
rect 880 49840 69120 49848
rect 880 49568 69200 49840
rect 381 49304 69200 49568
rect 880 49024 69200 49304
rect 381 48760 69200 49024
rect 880 48480 69200 48760
rect 381 48352 69200 48480
rect 880 48080 69200 48352
rect 880 48072 69120 48080
rect 381 47808 69120 48072
rect 880 47800 69120 47808
rect 880 47528 69200 47800
rect 381 47264 69200 47528
rect 880 46984 69200 47264
rect 381 46856 69200 46984
rect 880 46576 69200 46856
rect 381 46312 69200 46576
rect 880 46040 69200 46312
rect 880 46032 69120 46040
rect 381 45768 69120 46032
rect 880 45760 69120 45768
rect 880 45488 69200 45760
rect 381 45224 69200 45488
rect 880 44944 69200 45224
rect 381 44816 69200 44944
rect 880 44536 69200 44816
rect 381 44272 69200 44536
rect 880 44000 69200 44272
rect 880 43992 69120 44000
rect 381 43728 69120 43992
rect 880 43720 69120 43728
rect 880 43448 69200 43720
rect 381 43320 69200 43448
rect 880 43040 69200 43320
rect 381 42776 69200 43040
rect 880 42496 69200 42776
rect 381 42232 69200 42496
rect 880 41960 69200 42232
rect 880 41952 69120 41960
rect 381 41824 69120 41952
rect 880 41680 69120 41824
rect 880 41544 69200 41680
rect 381 41280 69200 41544
rect 880 41000 69200 41280
rect 381 40736 69200 41000
rect 880 40456 69200 40736
rect 381 40328 69200 40456
rect 880 40048 69200 40328
rect 381 39920 69200 40048
rect 381 39784 69120 39920
rect 880 39640 69120 39784
rect 880 39504 69200 39640
rect 381 39240 69200 39504
rect 880 38960 69200 39240
rect 381 38832 69200 38960
rect 880 38552 69200 38832
rect 381 38288 69200 38552
rect 880 38008 69200 38288
rect 381 37880 69200 38008
rect 381 37744 69120 37880
rect 880 37600 69120 37744
rect 880 37464 69200 37600
rect 381 37336 69200 37464
rect 880 37056 69200 37336
rect 381 36792 69200 37056
rect 880 36512 69200 36792
rect 381 36248 69200 36512
rect 880 35968 69200 36248
rect 381 35840 69200 35968
rect 880 35560 69120 35840
rect 381 35296 69200 35560
rect 880 35016 69200 35296
rect 381 34752 69200 35016
rect 880 34472 69200 34752
rect 381 34344 69200 34472
rect 880 34064 69200 34344
rect 381 33800 69200 34064
rect 880 33520 69120 33800
rect 381 33256 69200 33520
rect 880 32976 69200 33256
rect 381 32848 69200 32976
rect 880 32568 69200 32848
rect 381 32304 69200 32568
rect 880 32024 69200 32304
rect 381 31760 69200 32024
rect 880 31480 69120 31760
rect 381 31352 69200 31480
rect 880 31072 69200 31352
rect 381 30808 69200 31072
rect 880 30528 69200 30808
rect 381 30264 69200 30528
rect 880 29984 69200 30264
rect 381 29720 69200 29984
rect 880 29440 69120 29720
rect 381 29312 69200 29440
rect 880 29032 69200 29312
rect 381 28768 69200 29032
rect 880 28488 69200 28768
rect 381 28224 69200 28488
rect 880 27944 69200 28224
rect 381 27816 69200 27944
rect 880 27680 69200 27816
rect 880 27536 69120 27680
rect 381 27400 69120 27536
rect 381 27272 69200 27400
rect 880 26992 69200 27272
rect 381 26728 69200 26992
rect 880 26448 69200 26728
rect 381 26320 69200 26448
rect 880 26040 69200 26320
rect 381 25776 69200 26040
rect 880 25640 69200 25776
rect 880 25496 69120 25640
rect 381 25360 69120 25496
rect 381 25232 69200 25360
rect 880 24952 69200 25232
rect 381 24824 69200 24952
rect 880 24544 69200 24824
rect 381 24280 69200 24544
rect 880 24000 69200 24280
rect 381 23736 69200 24000
rect 880 23600 69200 23736
rect 880 23456 69120 23600
rect 381 23328 69120 23456
rect 880 23320 69120 23328
rect 880 23048 69200 23320
rect 381 22784 69200 23048
rect 880 22504 69200 22784
rect 381 22240 69200 22504
rect 880 21960 69200 22240
rect 381 21832 69200 21960
rect 880 21560 69200 21832
rect 880 21552 69120 21560
rect 381 21288 69120 21552
rect 880 21280 69120 21288
rect 880 21008 69200 21280
rect 381 20744 69200 21008
rect 880 20464 69200 20744
rect 381 20336 69200 20464
rect 880 20056 69200 20336
rect 381 19792 69200 20056
rect 880 19520 69200 19792
rect 880 19512 69120 19520
rect 381 19248 69120 19512
rect 880 19240 69120 19248
rect 880 18968 69200 19240
rect 381 18840 69200 18968
rect 880 18560 69200 18840
rect 381 18296 69200 18560
rect 880 18016 69200 18296
rect 381 17752 69200 18016
rect 880 17480 69200 17752
rect 880 17472 69120 17480
rect 381 17344 69120 17472
rect 880 17200 69120 17344
rect 880 17064 69200 17200
rect 381 16800 69200 17064
rect 880 16520 69200 16800
rect 381 16256 69200 16520
rect 880 15976 69200 16256
rect 381 15848 69200 15976
rect 880 15568 69200 15848
rect 381 15440 69200 15568
rect 381 15304 69120 15440
rect 880 15160 69120 15304
rect 880 15024 69200 15160
rect 381 14760 69200 15024
rect 880 14480 69200 14760
rect 381 14216 69200 14480
rect 880 13936 69200 14216
rect 381 13808 69200 13936
rect 880 13528 69200 13808
rect 381 13400 69200 13528
rect 381 13264 69120 13400
rect 880 13120 69120 13264
rect 880 12984 69200 13120
rect 381 12720 69200 12984
rect 880 12440 69200 12720
rect 381 12312 69200 12440
rect 880 12032 69200 12312
rect 381 11768 69200 12032
rect 880 11488 69200 11768
rect 381 11360 69200 11488
rect 381 11224 69120 11360
rect 880 11080 69120 11224
rect 880 10944 69200 11080
rect 381 10816 69200 10944
rect 880 10536 69200 10816
rect 381 10272 69200 10536
rect 880 9992 69200 10272
rect 381 9728 69200 9992
rect 880 9448 69200 9728
rect 381 9320 69200 9448
rect 880 9040 69120 9320
rect 381 8776 69200 9040
rect 880 8496 69200 8776
rect 381 8232 69200 8496
rect 880 7952 69200 8232
rect 381 7824 69200 7952
rect 880 7544 69200 7824
rect 381 7280 69200 7544
rect 880 7000 69120 7280
rect 381 6736 69200 7000
rect 880 6456 69200 6736
rect 381 6328 69200 6456
rect 880 6048 69200 6328
rect 381 5784 69200 6048
rect 880 5504 69200 5784
rect 381 5240 69200 5504
rect 880 4960 69120 5240
rect 381 4832 69200 4960
rect 880 4552 69200 4832
rect 381 4288 69200 4552
rect 880 4008 69200 4288
rect 381 3744 69200 4008
rect 880 3464 69200 3744
rect 381 3336 69200 3464
rect 880 3200 69200 3336
rect 880 3056 69120 3200
rect 381 2920 69120 3056
rect 381 2792 69200 2920
rect 880 2512 69200 2792
rect 381 2248 69200 2512
rect 880 1968 69200 2248
rect 381 1840 69200 1968
rect 880 1560 69200 1840
rect 381 1296 69200 1560
rect 880 1160 69200 1296
rect 880 1016 69120 1160
rect 381 880 69120 1016
rect 381 752 69200 880
rect 880 472 69200 752
rect 381 344 69200 472
rect 880 171 69200 344
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
<< obsm4 >>
rect 614 3707 4128 197165
rect 4608 3707 19488 197165
rect 19968 3707 34848 197165
rect 35328 3707 45389 197165
<< labels >>
rlabel metal2 s 10782 0 10838 800 6 master0_wb_ack_i
port 1 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 master0_wb_adr_o[0]
port 2 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 master0_wb_adr_o[10]
port 3 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 master0_wb_adr_o[11]
port 4 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 master0_wb_adr_o[12]
port 5 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 master0_wb_adr_o[13]
port 6 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 master0_wb_adr_o[14]
port 7 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 master0_wb_adr_o[15]
port 8 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 master0_wb_adr_o[16]
port 9 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 master0_wb_adr_o[17]
port 10 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 master0_wb_adr_o[18]
port 11 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 master0_wb_adr_o[19]
port 12 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 master0_wb_adr_o[1]
port 13 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 master0_wb_adr_o[20]
port 14 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 master0_wb_adr_o[21]
port 15 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 master0_wb_adr_o[22]
port 16 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 master0_wb_adr_o[23]
port 17 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 master0_wb_adr_o[24]
port 18 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 master0_wb_adr_o[25]
port 19 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 master0_wb_adr_o[26]
port 20 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 master0_wb_adr_o[27]
port 21 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 master0_wb_adr_o[2]
port 22 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 master0_wb_adr_o[3]
port 23 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 master0_wb_adr_o[4]
port 24 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 master0_wb_adr_o[5]
port 25 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 master0_wb_adr_o[6]
port 26 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 master0_wb_adr_o[7]
port 27 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 master0_wb_adr_o[8]
port 28 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 master0_wb_adr_o[9]
port 29 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 master0_wb_cyc_o
port 30 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 master0_wb_data_i[0]
port 31 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 master0_wb_data_i[10]
port 32 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 master0_wb_data_i[11]
port 33 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 master0_wb_data_i[12]
port 34 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 master0_wb_data_i[13]
port 35 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 master0_wb_data_i[14]
port 36 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 master0_wb_data_i[15]
port 37 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 master0_wb_data_i[16]
port 38 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 master0_wb_data_i[17]
port 39 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 master0_wb_data_i[18]
port 40 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 master0_wb_data_i[19]
port 41 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 master0_wb_data_i[1]
port 42 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 master0_wb_data_i[20]
port 43 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 master0_wb_data_i[21]
port 44 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 master0_wb_data_i[22]
port 45 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 master0_wb_data_i[23]
port 46 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 master0_wb_data_i[24]
port 47 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 master0_wb_data_i[25]
port 48 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 master0_wb_data_i[26]
port 49 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 master0_wb_data_i[27]
port 50 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 master0_wb_data_i[28]
port 51 nsew signal output
rlabel metal2 s 66718 0 66774 800 6 master0_wb_data_i[29]
port 52 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 master0_wb_data_i[2]
port 53 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 master0_wb_data_i[30]
port 54 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 master0_wb_data_i[31]
port 55 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 master0_wb_data_i[3]
port 56 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 master0_wb_data_i[4]
port 57 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 master0_wb_data_i[5]
port 58 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 master0_wb_data_i[6]
port 59 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 master0_wb_data_i[7]
port 60 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 master0_wb_data_i[8]
port 61 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 master0_wb_data_i[9]
port 62 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 master0_wb_data_o[0]
port 63 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 master0_wb_data_o[10]
port 64 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 master0_wb_data_o[11]
port 65 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 master0_wb_data_o[12]
port 66 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 master0_wb_data_o[13]
port 67 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 master0_wb_data_o[14]
port 68 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 master0_wb_data_o[15]
port 69 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 master0_wb_data_o[16]
port 70 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 master0_wb_data_o[17]
port 71 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 master0_wb_data_o[18]
port 72 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 master0_wb_data_o[19]
port 73 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 master0_wb_data_o[1]
port 74 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 master0_wb_data_o[20]
port 75 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 master0_wb_data_o[21]
port 76 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 master0_wb_data_o[22]
port 77 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 master0_wb_data_o[23]
port 78 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 master0_wb_data_o[24]
port 79 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 master0_wb_data_o[25]
port 80 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 master0_wb_data_o[26]
port 81 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 master0_wb_data_o[27]
port 82 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 master0_wb_data_o[28]
port 83 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 master0_wb_data_o[29]
port 84 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 master0_wb_data_o[2]
port 85 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 master0_wb_data_o[30]
port 86 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 master0_wb_data_o[31]
port 87 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 master0_wb_data_o[3]
port 88 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 master0_wb_data_o[4]
port 89 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 master0_wb_data_o[5]
port 90 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 master0_wb_data_o[6]
port 91 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 master0_wb_data_o[7]
port 92 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 master0_wb_data_o[8]
port 93 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 master0_wb_data_o[9]
port 94 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 master0_wb_error_i
port 95 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 master0_wb_sel_o[0]
port 96 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 master0_wb_sel_o[1]
port 97 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 master0_wb_sel_o[2]
port 98 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 master0_wb_sel_o[3]
port 99 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 master0_wb_stall_i
port 100 nsew signal output
rlabel metal2 s 13082 0 13138 800 6 master0_wb_stb_o
port 101 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 master0_wb_we_o
port 102 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 master1_wb_ack_i
port 103 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 master1_wb_adr_o[0]
port 104 nsew signal input
rlabel metal3 s 0 120096 800 120216 6 master1_wb_adr_o[10]
port 105 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 master1_wb_adr_o[11]
port 106 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 master1_wb_adr_o[12]
port 107 nsew signal input
rlabel metal3 s 0 124584 800 124704 6 master1_wb_adr_o[13]
port 108 nsew signal input
rlabel metal3 s 0 126080 800 126200 6 master1_wb_adr_o[14]
port 109 nsew signal input
rlabel metal3 s 0 127576 800 127696 6 master1_wb_adr_o[15]
port 110 nsew signal input
rlabel metal3 s 0 129072 800 129192 6 master1_wb_adr_o[16]
port 111 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 master1_wb_adr_o[17]
port 112 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 master1_wb_adr_o[18]
port 113 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 master1_wb_adr_o[19]
port 114 nsew signal input
rlabel metal3 s 0 105136 800 105256 6 master1_wb_adr_o[1]
port 115 nsew signal input
rlabel metal3 s 0 135056 800 135176 6 master1_wb_adr_o[20]
port 116 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 master1_wb_adr_o[21]
port 117 nsew signal input
rlabel metal3 s 0 138048 800 138168 6 master1_wb_adr_o[22]
port 118 nsew signal input
rlabel metal3 s 0 139680 800 139800 6 master1_wb_adr_o[23]
port 119 nsew signal input
rlabel metal3 s 0 141176 800 141296 6 master1_wb_adr_o[24]
port 120 nsew signal input
rlabel metal3 s 0 142672 800 142792 6 master1_wb_adr_o[25]
port 121 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 master1_wb_adr_o[26]
port 122 nsew signal input
rlabel metal3 s 0 145664 800 145784 6 master1_wb_adr_o[27]
port 123 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 master1_wb_adr_o[2]
port 124 nsew signal input
rlabel metal3 s 0 109080 800 109200 6 master1_wb_adr_o[3]
port 125 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 master1_wb_adr_o[4]
port 126 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 master1_wb_adr_o[5]
port 127 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 master1_wb_adr_o[6]
port 128 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 master1_wb_adr_o[7]
port 129 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 master1_wb_adr_o[8]
port 130 nsew signal input
rlabel metal3 s 0 118600 800 118720 6 master1_wb_adr_o[9]
port 131 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 master1_wb_cyc_o
port 132 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 master1_wb_data_i[0]
port 133 nsew signal output
rlabel metal3 s 0 120640 800 120760 6 master1_wb_data_i[10]
port 134 nsew signal output
rlabel metal3 s 0 122136 800 122256 6 master1_wb_data_i[11]
port 135 nsew signal output
rlabel metal3 s 0 123632 800 123752 6 master1_wb_data_i[12]
port 136 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 master1_wb_data_i[13]
port 137 nsew signal output
rlabel metal3 s 0 126624 800 126744 6 master1_wb_data_i[14]
port 138 nsew signal output
rlabel metal3 s 0 128120 800 128240 6 master1_wb_data_i[15]
port 139 nsew signal output
rlabel metal3 s 0 129616 800 129736 6 master1_wb_data_i[16]
port 140 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 master1_wb_data_i[17]
port 141 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 master1_wb_data_i[18]
port 142 nsew signal output
rlabel metal3 s 0 134104 800 134224 6 master1_wb_data_i[19]
port 143 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 master1_wb_data_i[1]
port 144 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 master1_wb_data_i[20]
port 145 nsew signal output
rlabel metal3 s 0 137096 800 137216 6 master1_wb_data_i[21]
port 146 nsew signal output
rlabel metal3 s 0 138592 800 138712 6 master1_wb_data_i[22]
port 147 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 master1_wb_data_i[23]
port 148 nsew signal output
rlabel metal3 s 0 141584 800 141704 6 master1_wb_data_i[24]
port 149 nsew signal output
rlabel metal3 s 0 143080 800 143200 6 master1_wb_data_i[25]
port 150 nsew signal output
rlabel metal3 s 0 144576 800 144696 6 master1_wb_data_i[26]
port 151 nsew signal output
rlabel metal3 s 0 146072 800 146192 6 master1_wb_data_i[27]
port 152 nsew signal output
rlabel metal3 s 0 147160 800 147280 6 master1_wb_data_i[28]
port 153 nsew signal output
rlabel metal3 s 0 148112 800 148232 6 master1_wb_data_i[29]
port 154 nsew signal output
rlabel metal3 s 0 107584 800 107704 6 master1_wb_data_i[2]
port 155 nsew signal output
rlabel metal3 s 0 149064 800 149184 6 master1_wb_data_i[30]
port 156 nsew signal output
rlabel metal3 s 0 150152 800 150272 6 master1_wb_data_i[31]
port 157 nsew signal output
rlabel metal3 s 0 109624 800 109744 6 master1_wb_data_i[3]
port 158 nsew signal output
rlabel metal3 s 0 111664 800 111784 6 master1_wb_data_i[4]
port 159 nsew signal output
rlabel metal3 s 0 113160 800 113280 6 master1_wb_data_i[5]
port 160 nsew signal output
rlabel metal3 s 0 114656 800 114776 6 master1_wb_data_i[6]
port 161 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 master1_wb_data_i[7]
port 162 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 master1_wb_data_i[8]
port 163 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 master1_wb_data_i[9]
port 164 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 master1_wb_data_o[0]
port 165 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 master1_wb_data_o[10]
port 166 nsew signal input
rlabel metal3 s 0 122544 800 122664 6 master1_wb_data_o[11]
port 167 nsew signal input
rlabel metal3 s 0 124176 800 124296 6 master1_wb_data_o[12]
port 168 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 master1_wb_data_o[13]
port 169 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 master1_wb_data_o[14]
port 170 nsew signal input
rlabel metal3 s 0 128664 800 128784 6 master1_wb_data_o[15]
port 171 nsew signal input
rlabel metal3 s 0 130160 800 130280 6 master1_wb_data_o[16]
port 172 nsew signal input
rlabel metal3 s 0 131656 800 131776 6 master1_wb_data_o[17]
port 173 nsew signal input
rlabel metal3 s 0 133152 800 133272 6 master1_wb_data_o[18]
port 174 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 master1_wb_data_o[19]
port 175 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 master1_wb_data_o[1]
port 176 nsew signal input
rlabel metal3 s 0 136144 800 136264 6 master1_wb_data_o[20]
port 177 nsew signal input
rlabel metal3 s 0 137640 800 137760 6 master1_wb_data_o[21]
port 178 nsew signal input
rlabel metal3 s 0 139136 800 139256 6 master1_wb_data_o[22]
port 179 nsew signal input
rlabel metal3 s 0 140632 800 140752 6 master1_wb_data_o[23]
port 180 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 master1_wb_data_o[24]
port 181 nsew signal input
rlabel metal3 s 0 143624 800 143744 6 master1_wb_data_o[25]
port 182 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 master1_wb_data_o[26]
port 183 nsew signal input
rlabel metal3 s 0 146616 800 146736 6 master1_wb_data_o[27]
port 184 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 master1_wb_data_o[28]
port 185 nsew signal input
rlabel metal3 s 0 148656 800 148776 6 master1_wb_data_o[29]
port 186 nsew signal input
rlabel metal3 s 0 108128 800 108248 6 master1_wb_data_o[2]
port 187 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 master1_wb_data_o[30]
port 188 nsew signal input
rlabel metal3 s 0 150560 800 150680 6 master1_wb_data_o[31]
port 189 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 master1_wb_data_o[3]
port 190 nsew signal input
rlabel metal3 s 0 112072 800 112192 6 master1_wb_data_o[4]
port 191 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 master1_wb_data_o[5]
port 192 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 master1_wb_data_o[6]
port 193 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 master1_wb_data_o[7]
port 194 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 master1_wb_data_o[8]
port 195 nsew signal input
rlabel metal3 s 0 119552 800 119672 6 master1_wb_data_o[9]
port 196 nsew signal input
rlabel metal3 s 0 101056 800 101176 6 master1_wb_error_i
port 197 nsew signal output
rlabel metal3 s 0 104592 800 104712 6 master1_wb_sel_o[0]
port 198 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 master1_wb_sel_o[1]
port 199 nsew signal input
rlabel metal3 s 0 108672 800 108792 6 master1_wb_sel_o[2]
port 200 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 master1_wb_sel_o[3]
port 201 nsew signal input
rlabel metal3 s 0 101600 800 101720 6 master1_wb_stall_i
port 202 nsew signal output
rlabel metal3 s 0 102144 800 102264 6 master1_wb_stb_o
port 203 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 master1_wb_we_o
port 204 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 master2_wb_ack_i
port 205 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 master2_wb_adr_o[0]
port 206 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 master2_wb_adr_o[10]
port 207 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 master2_wb_adr_o[11]
port 208 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 master2_wb_adr_o[12]
port 209 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 master2_wb_adr_o[13]
port 210 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 master2_wb_adr_o[14]
port 211 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 master2_wb_adr_o[15]
port 212 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 master2_wb_adr_o[16]
port 213 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 master2_wb_adr_o[17]
port 214 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 master2_wb_adr_o[18]
port 215 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 master2_wb_adr_o[19]
port 216 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 master2_wb_adr_o[1]
port 217 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 master2_wb_adr_o[20]
port 218 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 master2_wb_adr_o[21]
port 219 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 master2_wb_adr_o[22]
port 220 nsew signal input
rlabel metal3 s 0 88544 800 88664 6 master2_wb_adr_o[23]
port 221 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 master2_wb_adr_o[24]
port 222 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 master2_wb_adr_o[25]
port 223 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 master2_wb_adr_o[26]
port 224 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 master2_wb_adr_o[27]
port 225 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 master2_wb_adr_o[2]
port 226 nsew signal input
rlabel metal3 s 0 58080 800 58200 6 master2_wb_adr_o[3]
port 227 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 master2_wb_adr_o[4]
port 228 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 master2_wb_adr_o[5]
port 229 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 master2_wb_adr_o[6]
port 230 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 master2_wb_adr_o[7]
port 231 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 master2_wb_adr_o[8]
port 232 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 master2_wb_adr_o[9]
port 233 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 master2_wb_cyc_o
port 234 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 master2_wb_data_i[0]
port 235 nsew signal output
rlabel metal3 s 0 69640 800 69760 6 master2_wb_data_i[10]
port 236 nsew signal output
rlabel metal3 s 0 71136 800 71256 6 master2_wb_data_i[11]
port 237 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 master2_wb_data_i[12]
port 238 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 master2_wb_data_i[13]
port 239 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 master2_wb_data_i[14]
port 240 nsew signal output
rlabel metal3 s 0 77120 800 77240 6 master2_wb_data_i[15]
port 241 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 master2_wb_data_i[16]
port 242 nsew signal output
rlabel metal3 s 0 80112 800 80232 6 master2_wb_data_i[17]
port 243 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 master2_wb_data_i[18]
port 244 nsew signal output
rlabel metal3 s 0 83104 800 83224 6 master2_wb_data_i[19]
port 245 nsew signal output
rlabel metal3 s 0 54544 800 54664 6 master2_wb_data_i[1]
port 246 nsew signal output
rlabel metal3 s 0 84600 800 84720 6 master2_wb_data_i[20]
port 247 nsew signal output
rlabel metal3 s 0 86096 800 86216 6 master2_wb_data_i[21]
port 248 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 master2_wb_data_i[22]
port 249 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 master2_wb_data_i[23]
port 250 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 master2_wb_data_i[24]
port 251 nsew signal output
rlabel metal3 s 0 92080 800 92200 6 master2_wb_data_i[25]
port 252 nsew signal output
rlabel metal3 s 0 93576 800 93696 6 master2_wb_data_i[26]
port 253 nsew signal output
rlabel metal3 s 0 95072 800 95192 6 master2_wb_data_i[27]
port 254 nsew signal output
rlabel metal3 s 0 96160 800 96280 6 master2_wb_data_i[28]
port 255 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 master2_wb_data_i[29]
port 256 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 master2_wb_data_i[2]
port 257 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 master2_wb_data_i[30]
port 258 nsew signal output
rlabel metal3 s 0 99152 800 99272 6 master2_wb_data_i[31]
port 259 nsew signal output
rlabel metal3 s 0 58624 800 58744 6 master2_wb_data_i[3]
port 260 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 master2_wb_data_i[4]
port 261 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 master2_wb_data_i[5]
port 262 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 master2_wb_data_i[6]
port 263 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 master2_wb_data_i[7]
port 264 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 master2_wb_data_i[8]
port 265 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 master2_wb_data_i[9]
port 266 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 master2_wb_data_o[0]
port 267 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 master2_wb_data_o[10]
port 268 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 master2_wb_data_o[11]
port 269 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 master2_wb_data_o[12]
port 270 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 master2_wb_data_o[13]
port 271 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 master2_wb_data_o[14]
port 272 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 master2_wb_data_o[15]
port 273 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 master2_wb_data_o[16]
port 274 nsew signal input
rlabel metal3 s 0 80656 800 80776 6 master2_wb_data_o[17]
port 275 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 master2_wb_data_o[18]
port 276 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 master2_wb_data_o[19]
port 277 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 master2_wb_data_o[1]
port 278 nsew signal input
rlabel metal3 s 0 85144 800 85264 6 master2_wb_data_o[20]
port 279 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 master2_wb_data_o[21]
port 280 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 master2_wb_data_o[22]
port 281 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 master2_wb_data_o[23]
port 282 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 master2_wb_data_o[24]
port 283 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 master2_wb_data_o[25]
port 284 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 master2_wb_data_o[26]
port 285 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 master2_wb_data_o[27]
port 286 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 master2_wb_data_o[28]
port 287 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 master2_wb_data_o[29]
port 288 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 master2_wb_data_o[2]
port 289 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 master2_wb_data_o[30]
port 290 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 master2_wb_data_o[31]
port 291 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 master2_wb_data_o[3]
port 292 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 master2_wb_data_o[4]
port 293 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 master2_wb_data_o[5]
port 294 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 master2_wb_data_o[6]
port 295 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 master2_wb_data_o[7]
port 296 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 master2_wb_data_o[8]
port 297 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 master2_wb_data_o[9]
port 298 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 master2_wb_error_i
port 299 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 master2_wb_sel_o[0]
port 300 nsew signal input
rlabel metal3 s 0 55632 800 55752 6 master2_wb_sel_o[1]
port 301 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 master2_wb_sel_o[2]
port 302 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 master2_wb_sel_o[3]
port 303 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 master2_wb_stall_i
port 304 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 master2_wb_stb_o
port 305 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 master2_wb_we_o
port 306 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 probe_master0_currentSlave[0]
port 307 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 probe_master0_currentSlave[1]
port 308 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 probe_master1_currentSlave[0]
port 309 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 probe_master1_currentSlave[1]
port 310 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 probe_master2_currentSlave[0]
port 311 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 probe_master2_currentSlave[1]
port 312 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 probe_master3_currentSlave[0]
port 313 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 probe_master3_currentSlave[1]
port 314 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 probe_slave0_currentMaster[0]
port 315 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 probe_slave0_currentMaster[1]
port 316 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 probe_slave1_currentMaster[0]
port 317 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 probe_slave1_currentMaster[1]
port 318 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 probe_slave2_currentMaster[0]
port 319 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 probe_slave2_currentMaster[1]
port 320 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 probe_slave3_currentMaster[0]
port 321 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 probe_slave3_currentMaster[1]
port 322 nsew signal output
rlabel metal3 s 0 151104 800 151224 6 slave0_wb_ack_o
port 323 nsew signal input
rlabel metal3 s 0 154096 800 154216 6 slave0_wb_adr_i[0]
port 324 nsew signal output
rlabel metal3 s 0 171096 800 171216 6 slave0_wb_adr_i[10]
port 325 nsew signal output
rlabel metal3 s 0 172592 800 172712 6 slave0_wb_adr_i[11]
port 326 nsew signal output
rlabel metal3 s 0 174088 800 174208 6 slave0_wb_adr_i[12]
port 327 nsew signal output
rlabel metal3 s 0 175584 800 175704 6 slave0_wb_adr_i[13]
port 328 nsew signal output
rlabel metal3 s 0 177080 800 177200 6 slave0_wb_adr_i[14]
port 329 nsew signal output
rlabel metal3 s 0 178576 800 178696 6 slave0_wb_adr_i[15]
port 330 nsew signal output
rlabel metal3 s 0 180072 800 180192 6 slave0_wb_adr_i[16]
port 331 nsew signal output
rlabel metal3 s 0 181568 800 181688 6 slave0_wb_adr_i[17]
port 332 nsew signal output
rlabel metal3 s 0 183064 800 183184 6 slave0_wb_adr_i[18]
port 333 nsew signal output
rlabel metal3 s 0 184560 800 184680 6 slave0_wb_adr_i[19]
port 334 nsew signal output
rlabel metal3 s 0 156136 800 156256 6 slave0_wb_adr_i[1]
port 335 nsew signal output
rlabel metal3 s 0 186192 800 186312 6 slave0_wb_adr_i[20]
port 336 nsew signal output
rlabel metal3 s 0 187688 800 187808 6 slave0_wb_adr_i[21]
port 337 nsew signal output
rlabel metal3 s 0 189184 800 189304 6 slave0_wb_adr_i[22]
port 338 nsew signal output
rlabel metal3 s 0 190680 800 190800 6 slave0_wb_adr_i[23]
port 339 nsew signal output
rlabel metal3 s 0 158176 800 158296 6 slave0_wb_adr_i[2]
port 340 nsew signal output
rlabel metal3 s 0 160080 800 160200 6 slave0_wb_adr_i[3]
port 341 nsew signal output
rlabel metal3 s 0 162120 800 162240 6 slave0_wb_adr_i[4]
port 342 nsew signal output
rlabel metal3 s 0 163616 800 163736 6 slave0_wb_adr_i[5]
port 343 nsew signal output
rlabel metal3 s 0 165112 800 165232 6 slave0_wb_adr_i[6]
port 344 nsew signal output
rlabel metal3 s 0 166608 800 166728 6 slave0_wb_adr_i[7]
port 345 nsew signal output
rlabel metal3 s 0 168104 800 168224 6 slave0_wb_adr_i[8]
port 346 nsew signal output
rlabel metal3 s 0 169600 800 169720 6 slave0_wb_adr_i[9]
port 347 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 slave0_wb_cyc_i
port 348 nsew signal output
rlabel metal3 s 0 154640 800 154760 6 slave0_wb_data_i[0]
port 349 nsew signal output
rlabel metal3 s 0 171640 800 171760 6 slave0_wb_data_i[10]
port 350 nsew signal output
rlabel metal3 s 0 173136 800 173256 6 slave0_wb_data_i[11]
port 351 nsew signal output
rlabel metal3 s 0 174632 800 174752 6 slave0_wb_data_i[12]
port 352 nsew signal output
rlabel metal3 s 0 176128 800 176248 6 slave0_wb_data_i[13]
port 353 nsew signal output
rlabel metal3 s 0 177624 800 177744 6 slave0_wb_data_i[14]
port 354 nsew signal output
rlabel metal3 s 0 179120 800 179240 6 slave0_wb_data_i[15]
port 355 nsew signal output
rlabel metal3 s 0 180616 800 180736 6 slave0_wb_data_i[16]
port 356 nsew signal output
rlabel metal3 s 0 182112 800 182232 6 slave0_wb_data_i[17]
port 357 nsew signal output
rlabel metal3 s 0 183608 800 183728 6 slave0_wb_data_i[18]
port 358 nsew signal output
rlabel metal3 s 0 185104 800 185224 6 slave0_wb_data_i[19]
port 359 nsew signal output
rlabel metal3 s 0 156680 800 156800 6 slave0_wb_data_i[1]
port 360 nsew signal output
rlabel metal3 s 0 186600 800 186720 6 slave0_wb_data_i[20]
port 361 nsew signal output
rlabel metal3 s 0 188096 800 188216 6 slave0_wb_data_i[21]
port 362 nsew signal output
rlabel metal3 s 0 189592 800 189712 6 slave0_wb_data_i[22]
port 363 nsew signal output
rlabel metal3 s 0 191088 800 191208 6 slave0_wb_data_i[23]
port 364 nsew signal output
rlabel metal3 s 0 192176 800 192296 6 slave0_wb_data_i[24]
port 365 nsew signal output
rlabel metal3 s 0 193128 800 193248 6 slave0_wb_data_i[25]
port 366 nsew signal output
rlabel metal3 s 0 194080 800 194200 6 slave0_wb_data_i[26]
port 367 nsew signal output
rlabel metal3 s 0 195168 800 195288 6 slave0_wb_data_i[27]
port 368 nsew signal output
rlabel metal3 s 0 196120 800 196240 6 slave0_wb_data_i[28]
port 369 nsew signal output
rlabel metal3 s 0 197072 800 197192 6 slave0_wb_data_i[29]
port 370 nsew signal output
rlabel metal3 s 0 158584 800 158704 6 slave0_wb_data_i[2]
port 371 nsew signal output
rlabel metal3 s 0 198160 800 198280 6 slave0_wb_data_i[30]
port 372 nsew signal output
rlabel metal3 s 0 199112 800 199232 6 slave0_wb_data_i[31]
port 373 nsew signal output
rlabel metal3 s 0 160624 800 160744 6 slave0_wb_data_i[3]
port 374 nsew signal output
rlabel metal3 s 0 162664 800 162784 6 slave0_wb_data_i[4]
port 375 nsew signal output
rlabel metal3 s 0 164160 800 164280 6 slave0_wb_data_i[5]
port 376 nsew signal output
rlabel metal3 s 0 165656 800 165776 6 slave0_wb_data_i[6]
port 377 nsew signal output
rlabel metal3 s 0 167152 800 167272 6 slave0_wb_data_i[7]
port 378 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 slave0_wb_data_i[8]
port 379 nsew signal output
rlabel metal3 s 0 170144 800 170264 6 slave0_wb_data_i[9]
port 380 nsew signal output
rlabel metal3 s 0 155184 800 155304 6 slave0_wb_data_o[0]
port 381 nsew signal input
rlabel metal3 s 0 172184 800 172304 6 slave0_wb_data_o[10]
port 382 nsew signal input
rlabel metal3 s 0 173680 800 173800 6 slave0_wb_data_o[11]
port 383 nsew signal input
rlabel metal3 s 0 175176 800 175296 6 slave0_wb_data_o[12]
port 384 nsew signal input
rlabel metal3 s 0 176672 800 176792 6 slave0_wb_data_o[13]
port 385 nsew signal input
rlabel metal3 s 0 178168 800 178288 6 slave0_wb_data_o[14]
port 386 nsew signal input
rlabel metal3 s 0 179664 800 179784 6 slave0_wb_data_o[15]
port 387 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 slave0_wb_data_o[16]
port 388 nsew signal input
rlabel metal3 s 0 182656 800 182776 6 slave0_wb_data_o[17]
port 389 nsew signal input
rlabel metal3 s 0 184152 800 184272 6 slave0_wb_data_o[18]
port 390 nsew signal input
rlabel metal3 s 0 185648 800 185768 6 slave0_wb_data_o[19]
port 391 nsew signal input
rlabel metal3 s 0 157088 800 157208 6 slave0_wb_data_o[1]
port 392 nsew signal input
rlabel metal3 s 0 187144 800 187264 6 slave0_wb_data_o[20]
port 393 nsew signal input
rlabel metal3 s 0 188640 800 188760 6 slave0_wb_data_o[21]
port 394 nsew signal input
rlabel metal3 s 0 190136 800 190256 6 slave0_wb_data_o[22]
port 395 nsew signal input
rlabel metal3 s 0 191632 800 191752 6 slave0_wb_data_o[23]
port 396 nsew signal input
rlabel metal3 s 0 192584 800 192704 6 slave0_wb_data_o[24]
port 397 nsew signal input
rlabel metal3 s 0 193672 800 193792 6 slave0_wb_data_o[25]
port 398 nsew signal input
rlabel metal3 s 0 194624 800 194744 6 slave0_wb_data_o[26]
port 399 nsew signal input
rlabel metal3 s 0 195576 800 195696 6 slave0_wb_data_o[27]
port 400 nsew signal input
rlabel metal3 s 0 196664 800 196784 6 slave0_wb_data_o[28]
port 401 nsew signal input
rlabel metal3 s 0 197616 800 197736 6 slave0_wb_data_o[29]
port 402 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 slave0_wb_data_o[2]
port 403 nsew signal input
rlabel metal3 s 0 198568 800 198688 6 slave0_wb_data_o[30]
port 404 nsew signal input
rlabel metal3 s 0 199656 800 199776 6 slave0_wb_data_o[31]
port 405 nsew signal input
rlabel metal3 s 0 161168 800 161288 6 slave0_wb_data_o[3]
port 406 nsew signal input
rlabel metal3 s 0 163072 800 163192 6 slave0_wb_data_o[4]
port 407 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 slave0_wb_data_o[5]
port 408 nsew signal input
rlabel metal3 s 0 166064 800 166184 6 slave0_wb_data_o[6]
port 409 nsew signal input
rlabel metal3 s 0 167560 800 167680 6 slave0_wb_data_o[7]
port 410 nsew signal input
rlabel metal3 s 0 169056 800 169176 6 slave0_wb_data_o[8]
port 411 nsew signal input
rlabel metal3 s 0 170688 800 170808 6 slave0_wb_data_o[9]
port 412 nsew signal input
rlabel metal3 s 0 152056 800 152176 6 slave0_wb_error_o
port 413 nsew signal input
rlabel metal3 s 0 155592 800 155712 6 slave0_wb_sel_i[0]
port 414 nsew signal output
rlabel metal3 s 0 157632 800 157752 6 slave0_wb_sel_i[1]
port 415 nsew signal output
rlabel metal3 s 0 159672 800 159792 6 slave0_wb_sel_i[2]
port 416 nsew signal output
rlabel metal3 s 0 161576 800 161696 6 slave0_wb_sel_i[3]
port 417 nsew signal output
rlabel metal3 s 0 152600 800 152720 6 slave0_wb_stall_o
port 418 nsew signal input
rlabel metal3 s 0 153144 800 153264 6 slave0_wb_stb_i
port 419 nsew signal output
rlabel metal3 s 0 153552 800 153672 6 slave0_wb_we_i
port 420 nsew signal output
rlabel metal3 s 0 144 800 264 6 slave1_wb_ack_o
port 421 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 slave1_wb_adr_i[0]
port 422 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 slave1_wb_adr_i[10]
port 423 nsew signal output
rlabel metal3 s 0 21632 800 21752 6 slave1_wb_adr_i[11]
port 424 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 slave1_wb_adr_i[12]
port 425 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 slave1_wb_adr_i[13]
port 426 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 slave1_wb_adr_i[14]
port 427 nsew signal output
rlabel metal3 s 0 27616 800 27736 6 slave1_wb_adr_i[15]
port 428 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 slave1_wb_adr_i[16]
port 429 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 slave1_wb_adr_i[17]
port 430 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 slave1_wb_adr_i[18]
port 431 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 slave1_wb_adr_i[19]
port 432 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 slave1_wb_adr_i[1]
port 433 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 slave1_wb_adr_i[20]
port 434 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 slave1_wb_adr_i[21]
port 435 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 slave1_wb_adr_i[22]
port 436 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 slave1_wb_adr_i[23]
port 437 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 slave1_wb_adr_i[2]
port 438 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 slave1_wb_adr_i[3]
port 439 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 slave1_wb_adr_i[4]
port 440 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 slave1_wb_adr_i[5]
port 441 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 slave1_wb_adr_i[6]
port 442 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 slave1_wb_adr_i[7]
port 443 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 slave1_wb_adr_i[8]
port 444 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 slave1_wb_adr_i[9]
port 445 nsew signal output
rlabel metal3 s 0 552 800 672 6 slave1_wb_cyc_i
port 446 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 slave1_wb_data_i[0]
port 447 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 slave1_wb_data_i[10]
port 448 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 slave1_wb_data_i[11]
port 449 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 slave1_wb_data_i[12]
port 450 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 slave1_wb_data_i[13]
port 451 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 slave1_wb_data_i[14]
port 452 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 slave1_wb_data_i[15]
port 453 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 slave1_wb_data_i[16]
port 454 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 slave1_wb_data_i[17]
port 455 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 slave1_wb_data_i[18]
port 456 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 slave1_wb_data_i[19]
port 457 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 slave1_wb_data_i[1]
port 458 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 slave1_wb_data_i[20]
port 459 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 slave1_wb_data_i[21]
port 460 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 slave1_wb_data_i[22]
port 461 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 slave1_wb_data_i[23]
port 462 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 slave1_wb_data_i[24]
port 463 nsew signal output
rlabel metal3 s 0 42032 800 42152 6 slave1_wb_data_i[25]
port 464 nsew signal output
rlabel metal3 s 0 43120 800 43240 6 slave1_wb_data_i[26]
port 465 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 slave1_wb_data_i[27]
port 466 nsew signal output
rlabel metal3 s 0 45024 800 45144 6 slave1_wb_data_i[28]
port 467 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 slave1_wb_data_i[29]
port 468 nsew signal output
rlabel metal3 s 0 7624 800 7744 6 slave1_wb_data_i[2]
port 469 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 slave1_wb_data_i[30]
port 470 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 slave1_wb_data_i[31]
port 471 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 slave1_wb_data_i[3]
port 472 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 slave1_wb_data_i[4]
port 473 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 slave1_wb_data_i[5]
port 474 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 slave1_wb_data_i[6]
port 475 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 slave1_wb_data_i[7]
port 476 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 slave1_wb_data_i[8]
port 477 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 slave1_wb_data_i[9]
port 478 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 slave1_wb_data_o[0]
port 479 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 slave1_wb_data_o[10]
port 480 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 slave1_wb_data_o[11]
port 481 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 slave1_wb_data_o[12]
port 482 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 slave1_wb_data_o[13]
port 483 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 slave1_wb_data_o[14]
port 484 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 slave1_wb_data_o[15]
port 485 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 slave1_wb_data_o[16]
port 486 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 slave1_wb_data_o[17]
port 487 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 slave1_wb_data_o[18]
port 488 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 slave1_wb_data_o[19]
port 489 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 slave1_wb_data_o[1]
port 490 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 slave1_wb_data_o[20]
port 491 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 slave1_wb_data_o[21]
port 492 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 slave1_wb_data_o[22]
port 493 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 slave1_wb_data_o[23]
port 494 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 slave1_wb_data_o[24]
port 495 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 slave1_wb_data_o[25]
port 496 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 slave1_wb_data_o[26]
port 497 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 slave1_wb_data_o[27]
port 498 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 slave1_wb_data_o[28]
port 499 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 slave1_wb_data_o[29]
port 500 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 slave1_wb_data_o[2]
port 501 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 slave1_wb_data_o[30]
port 502 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 slave1_wb_data_o[31]
port 503 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 slave1_wb_data_o[3]
port 504 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 slave1_wb_data_o[4]
port 505 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 slave1_wb_data_o[5]
port 506 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 slave1_wb_data_o[6]
port 507 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 slave1_wb_data_o[7]
port 508 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 slave1_wb_data_o[8]
port 509 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 slave1_wb_data_o[9]
port 510 nsew signal input
rlabel metal3 s 0 1096 800 1216 6 slave1_wb_error_o
port 511 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 slave1_wb_sel_i[0]
port 512 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 slave1_wb_sel_i[1]
port 513 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 slave1_wb_sel_i[2]
port 514 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 slave1_wb_sel_i[3]
port 515 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 slave1_wb_stall_o
port 516 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 slave1_wb_stb_i
port 517 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 slave1_wb_we_i
port 518 nsew signal output
rlabel metal2 s 294 199200 350 200000 6 slave2_wb_ack_o
port 519 nsew signal input
rlabel metal2 s 4526 199200 4582 200000 6 slave2_wb_adr_i[0]
port 520 nsew signal output
rlabel metal2 s 28814 199200 28870 200000 6 slave2_wb_adr_i[10]
port 521 nsew signal output
rlabel metal2 s 30930 199200 30986 200000 6 slave2_wb_adr_i[11]
port 522 nsew signal output
rlabel metal2 s 33138 199200 33194 200000 6 slave2_wb_adr_i[12]
port 523 nsew signal output
rlabel metal2 s 35254 199200 35310 200000 6 slave2_wb_adr_i[13]
port 524 nsew signal output
rlabel metal2 s 37370 199200 37426 200000 6 slave2_wb_adr_i[14]
port 525 nsew signal output
rlabel metal2 s 39578 199200 39634 200000 6 slave2_wb_adr_i[15]
port 526 nsew signal output
rlabel metal2 s 41694 199200 41750 200000 6 slave2_wb_adr_i[16]
port 527 nsew signal output
rlabel metal2 s 43810 199200 43866 200000 6 slave2_wb_adr_i[17]
port 528 nsew signal output
rlabel metal2 s 45926 199200 45982 200000 6 slave2_wb_adr_i[18]
port 529 nsew signal output
rlabel metal2 s 48134 199200 48190 200000 6 slave2_wb_adr_i[19]
port 530 nsew signal output
rlabel metal2 s 7378 199200 7434 200000 6 slave2_wb_adr_i[1]
port 531 nsew signal output
rlabel metal2 s 50250 199200 50306 200000 6 slave2_wb_adr_i[20]
port 532 nsew signal output
rlabel metal2 s 52366 199200 52422 200000 6 slave2_wb_adr_i[21]
port 533 nsew signal output
rlabel metal2 s 54574 199200 54630 200000 6 slave2_wb_adr_i[22]
port 534 nsew signal output
rlabel metal2 s 56690 199200 56746 200000 6 slave2_wb_adr_i[23]
port 535 nsew signal output
rlabel metal2 s 10230 199200 10286 200000 6 slave2_wb_adr_i[2]
port 536 nsew signal output
rlabel metal2 s 13082 199200 13138 200000 6 slave2_wb_adr_i[3]
port 537 nsew signal output
rlabel metal2 s 15934 199200 15990 200000 6 slave2_wb_adr_i[4]
port 538 nsew signal output
rlabel metal2 s 18142 199200 18198 200000 6 slave2_wb_adr_i[5]
port 539 nsew signal output
rlabel metal2 s 20258 199200 20314 200000 6 slave2_wb_adr_i[6]
port 540 nsew signal output
rlabel metal2 s 22374 199200 22430 200000 6 slave2_wb_adr_i[7]
port 541 nsew signal output
rlabel metal2 s 24582 199200 24638 200000 6 slave2_wb_adr_i[8]
port 542 nsew signal output
rlabel metal2 s 26698 199200 26754 200000 6 slave2_wb_adr_i[9]
port 543 nsew signal output
rlabel metal2 s 938 199200 994 200000 6 slave2_wb_cyc_i
port 544 nsew signal output
rlabel metal2 s 5262 199200 5318 200000 6 slave2_wb_data_i[0]
port 545 nsew signal output
rlabel metal2 s 29550 199200 29606 200000 6 slave2_wb_data_i[10]
port 546 nsew signal output
rlabel metal2 s 31666 199200 31722 200000 6 slave2_wb_data_i[11]
port 547 nsew signal output
rlabel metal2 s 33782 199200 33838 200000 6 slave2_wb_data_i[12]
port 548 nsew signal output
rlabel metal2 s 35990 199200 36046 200000 6 slave2_wb_data_i[13]
port 549 nsew signal output
rlabel metal2 s 38106 199200 38162 200000 6 slave2_wb_data_i[14]
port 550 nsew signal output
rlabel metal2 s 40222 199200 40278 200000 6 slave2_wb_data_i[15]
port 551 nsew signal output
rlabel metal2 s 42430 199200 42486 200000 6 slave2_wb_data_i[16]
port 552 nsew signal output
rlabel metal2 s 44546 199200 44602 200000 6 slave2_wb_data_i[17]
port 553 nsew signal output
rlabel metal2 s 46662 199200 46718 200000 6 slave2_wb_data_i[18]
port 554 nsew signal output
rlabel metal2 s 48870 199200 48926 200000 6 slave2_wb_data_i[19]
port 555 nsew signal output
rlabel metal2 s 8114 199200 8170 200000 6 slave2_wb_data_i[1]
port 556 nsew signal output
rlabel metal2 s 50986 199200 51042 200000 6 slave2_wb_data_i[20]
port 557 nsew signal output
rlabel metal2 s 53102 199200 53158 200000 6 slave2_wb_data_i[21]
port 558 nsew signal output
rlabel metal2 s 55218 199200 55274 200000 6 slave2_wb_data_i[22]
port 559 nsew signal output
rlabel metal2 s 57426 199200 57482 200000 6 slave2_wb_data_i[23]
port 560 nsew signal output
rlabel metal2 s 58806 199200 58862 200000 6 slave2_wb_data_i[24]
port 561 nsew signal output
rlabel metal2 s 60278 199200 60334 200000 6 slave2_wb_data_i[25]
port 562 nsew signal output
rlabel metal2 s 61658 199200 61714 200000 6 slave2_wb_data_i[26]
port 563 nsew signal output
rlabel metal2 s 63130 199200 63186 200000 6 slave2_wb_data_i[27]
port 564 nsew signal output
rlabel metal2 s 64510 199200 64566 200000 6 slave2_wb_data_i[28]
port 565 nsew signal output
rlabel metal2 s 65982 199200 66038 200000 6 slave2_wb_data_i[29]
port 566 nsew signal output
rlabel metal2 s 10966 199200 11022 200000 6 slave2_wb_data_i[2]
port 567 nsew signal output
rlabel metal2 s 67362 199200 67418 200000 6 slave2_wb_data_i[30]
port 568 nsew signal output
rlabel metal2 s 68834 199200 68890 200000 6 slave2_wb_data_i[31]
port 569 nsew signal output
rlabel metal2 s 13818 199200 13874 200000 6 slave2_wb_data_i[3]
port 570 nsew signal output
rlabel metal2 s 16670 199200 16726 200000 6 slave2_wb_data_i[4]
port 571 nsew signal output
rlabel metal2 s 18786 199200 18842 200000 6 slave2_wb_data_i[5]
port 572 nsew signal output
rlabel metal2 s 20994 199200 21050 200000 6 slave2_wb_data_i[6]
port 573 nsew signal output
rlabel metal2 s 23110 199200 23166 200000 6 slave2_wb_data_i[7]
port 574 nsew signal output
rlabel metal2 s 25226 199200 25282 200000 6 slave2_wb_data_i[8]
port 575 nsew signal output
rlabel metal2 s 27434 199200 27490 200000 6 slave2_wb_data_i[9]
port 576 nsew signal output
rlabel metal2 s 5998 199200 6054 200000 6 slave2_wb_data_o[0]
port 577 nsew signal input
rlabel metal2 s 30286 199200 30342 200000 6 slave2_wb_data_o[10]
port 578 nsew signal input
rlabel metal2 s 32402 199200 32458 200000 6 slave2_wb_data_o[11]
port 579 nsew signal input
rlabel metal2 s 34518 199200 34574 200000 6 slave2_wb_data_o[12]
port 580 nsew signal input
rlabel metal2 s 36726 199200 36782 200000 6 slave2_wb_data_o[13]
port 581 nsew signal input
rlabel metal2 s 38842 199200 38898 200000 6 slave2_wb_data_o[14]
port 582 nsew signal input
rlabel metal2 s 40958 199200 41014 200000 6 slave2_wb_data_o[15]
port 583 nsew signal input
rlabel metal2 s 43074 199200 43130 200000 6 slave2_wb_data_o[16]
port 584 nsew signal input
rlabel metal2 s 45282 199200 45338 200000 6 slave2_wb_data_o[17]
port 585 nsew signal input
rlabel metal2 s 47398 199200 47454 200000 6 slave2_wb_data_o[18]
port 586 nsew signal input
rlabel metal2 s 49514 199200 49570 200000 6 slave2_wb_data_o[19]
port 587 nsew signal input
rlabel metal2 s 8850 199200 8906 200000 6 slave2_wb_data_o[1]
port 588 nsew signal input
rlabel metal2 s 51722 199200 51778 200000 6 slave2_wb_data_o[20]
port 589 nsew signal input
rlabel metal2 s 53838 199200 53894 200000 6 slave2_wb_data_o[21]
port 590 nsew signal input
rlabel metal2 s 55954 199200 56010 200000 6 slave2_wb_data_o[22]
port 591 nsew signal input
rlabel metal2 s 58070 199200 58126 200000 6 slave2_wb_data_o[23]
port 592 nsew signal input
rlabel metal2 s 59542 199200 59598 200000 6 slave2_wb_data_o[24]
port 593 nsew signal input
rlabel metal2 s 61014 199200 61070 200000 6 slave2_wb_data_o[25]
port 594 nsew signal input
rlabel metal2 s 62394 199200 62450 200000 6 slave2_wb_data_o[26]
port 595 nsew signal input
rlabel metal2 s 63866 199200 63922 200000 6 slave2_wb_data_o[27]
port 596 nsew signal input
rlabel metal2 s 65246 199200 65302 200000 6 slave2_wb_data_o[28]
port 597 nsew signal input
rlabel metal2 s 66718 199200 66774 200000 6 slave2_wb_data_o[29]
port 598 nsew signal input
rlabel metal2 s 11702 199200 11758 200000 6 slave2_wb_data_o[2]
port 599 nsew signal input
rlabel metal2 s 68098 199200 68154 200000 6 slave2_wb_data_o[30]
port 600 nsew signal input
rlabel metal2 s 69570 199200 69626 200000 6 slave2_wb_data_o[31]
port 601 nsew signal input
rlabel metal2 s 14554 199200 14610 200000 6 slave2_wb_data_o[3]
port 602 nsew signal input
rlabel metal2 s 17406 199200 17462 200000 6 slave2_wb_data_o[4]
port 603 nsew signal input
rlabel metal2 s 19522 199200 19578 200000 6 slave2_wb_data_o[5]
port 604 nsew signal input
rlabel metal2 s 21638 199200 21694 200000 6 slave2_wb_data_o[6]
port 605 nsew signal input
rlabel metal2 s 23846 199200 23902 200000 6 slave2_wb_data_o[7]
port 606 nsew signal input
rlabel metal2 s 25962 199200 26018 200000 6 slave2_wb_data_o[8]
port 607 nsew signal input
rlabel metal2 s 28078 199200 28134 200000 6 slave2_wb_data_o[9]
port 608 nsew signal input
rlabel metal2 s 1674 199200 1730 200000 6 slave2_wb_error_o
port 609 nsew signal input
rlabel metal2 s 6642 199200 6698 200000 6 slave2_wb_sel_i[0]
port 610 nsew signal output
rlabel metal2 s 9494 199200 9550 200000 6 slave2_wb_sel_i[1]
port 611 nsew signal output
rlabel metal2 s 12438 199200 12494 200000 6 slave2_wb_sel_i[2]
port 612 nsew signal output
rlabel metal2 s 15290 199200 15346 200000 6 slave2_wb_sel_i[3]
port 613 nsew signal output
rlabel metal2 s 2410 199200 2466 200000 6 slave2_wb_stall_o
port 614 nsew signal input
rlabel metal2 s 3146 199200 3202 200000 6 slave2_wb_stb_i
port 615 nsew signal output
rlabel metal2 s 3790 199200 3846 200000 6 slave2_wb_we_i
port 616 nsew signal output
rlabel metal3 s 69200 960 70000 1080 6 slave3_wb_ack_o
port 617 nsew signal input
rlabel metal3 s 69200 13200 70000 13320 6 slave3_wb_adr_i[0]
port 618 nsew signal output
rlabel metal3 s 69200 82560 70000 82680 6 slave3_wb_adr_i[10]
port 619 nsew signal output
rlabel metal3 s 69200 88680 70000 88800 6 slave3_wb_adr_i[11]
port 620 nsew signal output
rlabel metal3 s 69200 94800 70000 94920 6 slave3_wb_adr_i[12]
port 621 nsew signal output
rlabel metal3 s 69200 100920 70000 101040 6 slave3_wb_adr_i[13]
port 622 nsew signal output
rlabel metal3 s 69200 107040 70000 107160 6 slave3_wb_adr_i[14]
port 623 nsew signal output
rlabel metal3 s 69200 113160 70000 113280 6 slave3_wb_adr_i[15]
port 624 nsew signal output
rlabel metal3 s 69200 119280 70000 119400 6 slave3_wb_adr_i[16]
port 625 nsew signal output
rlabel metal3 s 69200 125400 70000 125520 6 slave3_wb_adr_i[17]
port 626 nsew signal output
rlabel metal3 s 69200 131520 70000 131640 6 slave3_wb_adr_i[18]
port 627 nsew signal output
rlabel metal3 s 69200 137640 70000 137760 6 slave3_wb_adr_i[19]
port 628 nsew signal output
rlabel metal3 s 69200 21360 70000 21480 6 slave3_wb_adr_i[1]
port 629 nsew signal output
rlabel metal3 s 69200 143760 70000 143880 6 slave3_wb_adr_i[20]
port 630 nsew signal output
rlabel metal3 s 69200 149880 70000 150000 6 slave3_wb_adr_i[21]
port 631 nsew signal output
rlabel metal3 s 69200 156000 70000 156120 6 slave3_wb_adr_i[22]
port 632 nsew signal output
rlabel metal3 s 69200 162120 70000 162240 6 slave3_wb_adr_i[23]
port 633 nsew signal output
rlabel metal3 s 69200 29520 70000 29640 6 slave3_wb_adr_i[2]
port 634 nsew signal output
rlabel metal3 s 69200 37680 70000 37800 6 slave3_wb_adr_i[3]
port 635 nsew signal output
rlabel metal3 s 69200 45840 70000 45960 6 slave3_wb_adr_i[4]
port 636 nsew signal output
rlabel metal3 s 69200 51960 70000 52080 6 slave3_wb_adr_i[5]
port 637 nsew signal output
rlabel metal3 s 69200 58080 70000 58200 6 slave3_wb_adr_i[6]
port 638 nsew signal output
rlabel metal3 s 69200 64200 70000 64320 6 slave3_wb_adr_i[7]
port 639 nsew signal output
rlabel metal3 s 69200 70320 70000 70440 6 slave3_wb_adr_i[8]
port 640 nsew signal output
rlabel metal3 s 69200 76440 70000 76560 6 slave3_wb_adr_i[9]
port 641 nsew signal output
rlabel metal3 s 69200 3000 70000 3120 6 slave3_wb_cyc_i
port 642 nsew signal output
rlabel metal3 s 69200 15240 70000 15360 6 slave3_wb_data_i[0]
port 643 nsew signal output
rlabel metal3 s 69200 84600 70000 84720 6 slave3_wb_data_i[10]
port 644 nsew signal output
rlabel metal3 s 69200 90720 70000 90840 6 slave3_wb_data_i[11]
port 645 nsew signal output
rlabel metal3 s 69200 96840 70000 96960 6 slave3_wb_data_i[12]
port 646 nsew signal output
rlabel metal3 s 69200 102960 70000 103080 6 slave3_wb_data_i[13]
port 647 nsew signal output
rlabel metal3 s 69200 109080 70000 109200 6 slave3_wb_data_i[14]
port 648 nsew signal output
rlabel metal3 s 69200 115200 70000 115320 6 slave3_wb_data_i[15]
port 649 nsew signal output
rlabel metal3 s 69200 121320 70000 121440 6 slave3_wb_data_i[16]
port 650 nsew signal output
rlabel metal3 s 69200 127440 70000 127560 6 slave3_wb_data_i[17]
port 651 nsew signal output
rlabel metal3 s 69200 133560 70000 133680 6 slave3_wb_data_i[18]
port 652 nsew signal output
rlabel metal3 s 69200 139680 70000 139800 6 slave3_wb_data_i[19]
port 653 nsew signal output
rlabel metal3 s 69200 23400 70000 23520 6 slave3_wb_data_i[1]
port 654 nsew signal output
rlabel metal3 s 69200 145800 70000 145920 6 slave3_wb_data_i[20]
port 655 nsew signal output
rlabel metal3 s 69200 151920 70000 152040 6 slave3_wb_data_i[21]
port 656 nsew signal output
rlabel metal3 s 69200 158040 70000 158160 6 slave3_wb_data_i[22]
port 657 nsew signal output
rlabel metal3 s 69200 164160 70000 164280 6 slave3_wb_data_i[23]
port 658 nsew signal output
rlabel metal3 s 69200 168240 70000 168360 6 slave3_wb_data_i[24]
port 659 nsew signal output
rlabel metal3 s 69200 172320 70000 172440 6 slave3_wb_data_i[25]
port 660 nsew signal output
rlabel metal3 s 69200 176400 70000 176520 6 slave3_wb_data_i[26]
port 661 nsew signal output
rlabel metal3 s 69200 180480 70000 180600 6 slave3_wb_data_i[27]
port 662 nsew signal output
rlabel metal3 s 69200 184560 70000 184680 6 slave3_wb_data_i[28]
port 663 nsew signal output
rlabel metal3 s 69200 188640 70000 188760 6 slave3_wb_data_i[29]
port 664 nsew signal output
rlabel metal3 s 69200 31560 70000 31680 6 slave3_wb_data_i[2]
port 665 nsew signal output
rlabel metal3 s 69200 192720 70000 192840 6 slave3_wb_data_i[30]
port 666 nsew signal output
rlabel metal3 s 69200 196800 70000 196920 6 slave3_wb_data_i[31]
port 667 nsew signal output
rlabel metal3 s 69200 39720 70000 39840 6 slave3_wb_data_i[3]
port 668 nsew signal output
rlabel metal3 s 69200 47880 70000 48000 6 slave3_wb_data_i[4]
port 669 nsew signal output
rlabel metal3 s 69200 54000 70000 54120 6 slave3_wb_data_i[5]
port 670 nsew signal output
rlabel metal3 s 69200 60120 70000 60240 6 slave3_wb_data_i[6]
port 671 nsew signal output
rlabel metal3 s 69200 66240 70000 66360 6 slave3_wb_data_i[7]
port 672 nsew signal output
rlabel metal3 s 69200 72360 70000 72480 6 slave3_wb_data_i[8]
port 673 nsew signal output
rlabel metal3 s 69200 78480 70000 78600 6 slave3_wb_data_i[9]
port 674 nsew signal output
rlabel metal3 s 69200 17280 70000 17400 6 slave3_wb_data_o[0]
port 675 nsew signal input
rlabel metal3 s 69200 86640 70000 86760 6 slave3_wb_data_o[10]
port 676 nsew signal input
rlabel metal3 s 69200 92760 70000 92880 6 slave3_wb_data_o[11]
port 677 nsew signal input
rlabel metal3 s 69200 98880 70000 99000 6 slave3_wb_data_o[12]
port 678 nsew signal input
rlabel metal3 s 69200 105000 70000 105120 6 slave3_wb_data_o[13]
port 679 nsew signal input
rlabel metal3 s 69200 111120 70000 111240 6 slave3_wb_data_o[14]
port 680 nsew signal input
rlabel metal3 s 69200 117240 70000 117360 6 slave3_wb_data_o[15]
port 681 nsew signal input
rlabel metal3 s 69200 123360 70000 123480 6 slave3_wb_data_o[16]
port 682 nsew signal input
rlabel metal3 s 69200 129480 70000 129600 6 slave3_wb_data_o[17]
port 683 nsew signal input
rlabel metal3 s 69200 135600 70000 135720 6 slave3_wb_data_o[18]
port 684 nsew signal input
rlabel metal3 s 69200 141720 70000 141840 6 slave3_wb_data_o[19]
port 685 nsew signal input
rlabel metal3 s 69200 25440 70000 25560 6 slave3_wb_data_o[1]
port 686 nsew signal input
rlabel metal3 s 69200 147840 70000 147960 6 slave3_wb_data_o[20]
port 687 nsew signal input
rlabel metal3 s 69200 153960 70000 154080 6 slave3_wb_data_o[21]
port 688 nsew signal input
rlabel metal3 s 69200 160080 70000 160200 6 slave3_wb_data_o[22]
port 689 nsew signal input
rlabel metal3 s 69200 166200 70000 166320 6 slave3_wb_data_o[23]
port 690 nsew signal input
rlabel metal3 s 69200 170280 70000 170400 6 slave3_wb_data_o[24]
port 691 nsew signal input
rlabel metal3 s 69200 174360 70000 174480 6 slave3_wb_data_o[25]
port 692 nsew signal input
rlabel metal3 s 69200 178440 70000 178560 6 slave3_wb_data_o[26]
port 693 nsew signal input
rlabel metal3 s 69200 182520 70000 182640 6 slave3_wb_data_o[27]
port 694 nsew signal input
rlabel metal3 s 69200 186600 70000 186720 6 slave3_wb_data_o[28]
port 695 nsew signal input
rlabel metal3 s 69200 190680 70000 190800 6 slave3_wb_data_o[29]
port 696 nsew signal input
rlabel metal3 s 69200 33600 70000 33720 6 slave3_wb_data_o[2]
port 697 nsew signal input
rlabel metal3 s 69200 194760 70000 194880 6 slave3_wb_data_o[30]
port 698 nsew signal input
rlabel metal3 s 69200 198840 70000 198960 6 slave3_wb_data_o[31]
port 699 nsew signal input
rlabel metal3 s 69200 41760 70000 41880 6 slave3_wb_data_o[3]
port 700 nsew signal input
rlabel metal3 s 69200 49920 70000 50040 6 slave3_wb_data_o[4]
port 701 nsew signal input
rlabel metal3 s 69200 56040 70000 56160 6 slave3_wb_data_o[5]
port 702 nsew signal input
rlabel metal3 s 69200 62160 70000 62280 6 slave3_wb_data_o[6]
port 703 nsew signal input
rlabel metal3 s 69200 68280 70000 68400 6 slave3_wb_data_o[7]
port 704 nsew signal input
rlabel metal3 s 69200 74400 70000 74520 6 slave3_wb_data_o[8]
port 705 nsew signal input
rlabel metal3 s 69200 80520 70000 80640 6 slave3_wb_data_o[9]
port 706 nsew signal input
rlabel metal3 s 69200 5040 70000 5160 6 slave3_wb_error_o
port 707 nsew signal input
rlabel metal3 s 69200 19320 70000 19440 6 slave3_wb_sel_i[0]
port 708 nsew signal output
rlabel metal3 s 69200 27480 70000 27600 6 slave3_wb_sel_i[1]
port 709 nsew signal output
rlabel metal3 s 69200 35640 70000 35760 6 slave3_wb_sel_i[2]
port 710 nsew signal output
rlabel metal3 s 69200 43800 70000 43920 6 slave3_wb_sel_i[3]
port 711 nsew signal output
rlabel metal3 s 69200 7080 70000 7200 6 slave3_wb_stall_o
port 712 nsew signal input
rlabel metal3 s 69200 9120 70000 9240 6 slave3_wb_stb_i
port 713 nsew signal output
rlabel metal3 s 69200 11160 70000 11280 6 slave3_wb_we_i
port 714 nsew signal output
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 715 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 715 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 715 nsew power input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 716 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 716 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 717 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_rst_i
port 718 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11035876
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/WishboneInterconnect/runs/WishboneInterconnect/results/finishing/WishboneInterconnect.magic.gds
string GDS_START 609466
<< end >>

