* NGSPICE file created from CaravelHost.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

.subckt CaravelHost caravel_uart_rx caravel_uart_tx caravel_wb_ack_i caravel_wb_adr_o[0]
+ caravel_wb_adr_o[10] caravel_wb_adr_o[11] caravel_wb_adr_o[12] caravel_wb_adr_o[13]
+ caravel_wb_adr_o[14] caravel_wb_adr_o[15] caravel_wb_adr_o[16] caravel_wb_adr_o[17]
+ caravel_wb_adr_o[18] caravel_wb_adr_o[19] caravel_wb_adr_o[1] caravel_wb_adr_o[20]
+ caravel_wb_adr_o[21] caravel_wb_adr_o[22] caravel_wb_adr_o[23] caravel_wb_adr_o[24]
+ caravel_wb_adr_o[25] caravel_wb_adr_o[26] caravel_wb_adr_o[27] caravel_wb_adr_o[2]
+ caravel_wb_adr_o[3] caravel_wb_adr_o[4] caravel_wb_adr_o[5] caravel_wb_adr_o[6]
+ caravel_wb_adr_o[7] caravel_wb_adr_o[8] caravel_wb_adr_o[9] caravel_wb_cyc_o caravel_wb_data_i[0]
+ caravel_wb_data_i[10] caravel_wb_data_i[11] caravel_wb_data_i[12] caravel_wb_data_i[13]
+ caravel_wb_data_i[14] caravel_wb_data_i[15] caravel_wb_data_i[16] caravel_wb_data_i[17]
+ caravel_wb_data_i[18] caravel_wb_data_i[19] caravel_wb_data_i[1] caravel_wb_data_i[20]
+ caravel_wb_data_i[21] caravel_wb_data_i[22] caravel_wb_data_i[23] caravel_wb_data_i[24]
+ caravel_wb_data_i[25] caravel_wb_data_i[26] caravel_wb_data_i[27] caravel_wb_data_i[28]
+ caravel_wb_data_i[29] caravel_wb_data_i[2] caravel_wb_data_i[30] caravel_wb_data_i[31]
+ caravel_wb_data_i[3] caravel_wb_data_i[4] caravel_wb_data_i[5] caravel_wb_data_i[6]
+ caravel_wb_data_i[7] caravel_wb_data_i[8] caravel_wb_data_i[9] caravel_wb_data_o[0]
+ caravel_wb_data_o[10] caravel_wb_data_o[11] caravel_wb_data_o[12] caravel_wb_data_o[13]
+ caravel_wb_data_o[14] caravel_wb_data_o[15] caravel_wb_data_o[16] caravel_wb_data_o[17]
+ caravel_wb_data_o[18] caravel_wb_data_o[19] caravel_wb_data_o[1] caravel_wb_data_o[20]
+ caravel_wb_data_o[21] caravel_wb_data_o[22] caravel_wb_data_o[23] caravel_wb_data_o[24]
+ caravel_wb_data_o[25] caravel_wb_data_o[26] caravel_wb_data_o[27] caravel_wb_data_o[28]
+ caravel_wb_data_o[29] caravel_wb_data_o[2] caravel_wb_data_o[30] caravel_wb_data_o[31]
+ caravel_wb_data_o[3] caravel_wb_data_o[4] caravel_wb_data_o[5] caravel_wb_data_o[6]
+ caravel_wb_data_o[7] caravel_wb_data_o[8] caravel_wb_data_o[9] caravel_wb_error_i
+ caravel_wb_sel_o[0] caravel_wb_sel_o[1] caravel_wb_sel_o[2] caravel_wb_sel_o[3]
+ caravel_wb_stall_i caravel_wb_stb_o caravel_wb_we_o vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_data_i[0] wbs_data_i[10] wbs_data_i[11] wbs_data_i[12]
+ wbs_data_i[13] wbs_data_i[14] wbs_data_i[15] wbs_data_i[16] wbs_data_i[17] wbs_data_i[18]
+ wbs_data_i[19] wbs_data_i[1] wbs_data_i[20] wbs_data_i[21] wbs_data_i[22] wbs_data_i[23]
+ wbs_data_i[24] wbs_data_i[25] wbs_data_i[26] wbs_data_i[27] wbs_data_i[28] wbs_data_i[29]
+ wbs_data_i[2] wbs_data_i[30] wbs_data_i[31] wbs_data_i[3] wbs_data_i[4] wbs_data_i[5]
+ wbs_data_i[6] wbs_data_i[7] wbs_data_i[8] wbs_data_i[9] wbs_data_o[0] wbs_data_o[10]
+ wbs_data_o[11] wbs_data_o[12] wbs_data_o[13] wbs_data_o[14] wbs_data_o[15] wbs_data_o[16]
+ wbs_data_o[17] wbs_data_o[18] wbs_data_o[19] wbs_data_o[1] wbs_data_o[20] wbs_data_o[21]
+ wbs_data_o[22] wbs_data_o[23] wbs_data_o[24] wbs_data_o[25] wbs_data_o[26] wbs_data_o[27]
+ wbs_data_o[28] wbs_data_o[29] wbs_data_o[2] wbs_data_o[30] wbs_data_o[31] wbs_data_o[3]
+ wbs_data_o[4] wbs_data_o[5] wbs_data_o[6] wbs_data_o[7] wbs_data_o[8] wbs_data_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6914_ _6914_/CLK _6914_/D vssd1 vssd1 vccd1 vccd1 _6914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6845_ _6845_/CLK _6845_/D vssd1 vssd1 vccd1 vccd1 _6845_/Q sky130_fd_sc_hd__dfxtp_1
X_6776_ _6776_/CLK _6776_/D vssd1 vssd1 vccd1 vccd1 _6776_/Q sky130_fd_sc_hd__dfxtp_1
X_3988_ _3977_/B _3988_/B _5774_/C vssd1 vssd1 vccd1 vccd1 _3989_/A sky130_fd_sc_hd__and3b_1
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5727_ _5727_/A vssd1 vssd1 vccd1 vccd1 _6744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5658_ _7005_/Q _5623_/X _5626_/Y _5642_/X _5657_/X vssd1 vssd1 vccd1 vccd1 _5669_/B
+ sky130_fd_sc_hd__a2111o_1
X_4609_ _4624_/S vssd1 vssd1 vccd1 vccd1 _4618_/S sky130_fd_sc_hd__buf_2
X_5589_ _5589_/A vssd1 vssd1 vccd1 vccd1 _6696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5524__355 _5528__359/A vssd1 vssd1 vccd1 vccd1 _6645_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4960_ _3968_/A _4955_/X _4959_/X _3974_/A vssd1 vssd1 vccd1 vccd1 _4960_/X sky130_fd_sc_hd__o211a_1
XFILLER_83_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4891_ _7044_/Q _4891_/B vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__or2_1
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3911_ _3911_/A vssd1 vssd1 vccd1 vccd1 _6790_/D sky130_fd_sc_hd__clkbuf_1
X_6630_ _6630_/CLK _6630_/D vssd1 vssd1 vccd1 vccd1 _6630_/Q sky130_fd_sc_hd__dfxtp_1
X_3842_ _3842_/A vssd1 vssd1 vccd1 vccd1 _6813_/D sky130_fd_sc_hd__clkbuf_1
X_6561_ _6561_/CLK _6561_/D vssd1 vssd1 vccd1 vccd1 _6561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3773_ _3773_/A vssd1 vssd1 vccd1 vccd1 _3773_/X sky130_fd_sc_hd__buf_2
X_6492_ _6492_/CLK _6492_/D vssd1 vssd1 vccd1 vccd1 _6492_/Q sky130_fd_sc_hd__dfxtp_1
X_5443_ _5324_/A _5442_/X _5321_/A vssd1 vssd1 vccd1 vccd1 _5443_/Y sky130_fd_sc_hd__o21ai_1
X_5374_ _5372_/X _5373_/X _5429_/S vssd1 vssd1 vccd1 vccd1 _5374_/X sky130_fd_sc_hd__mux2_1
X_7113_ _7113_/A vssd1 vssd1 vccd1 vccd1 _7113_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4325_ _4325_/A vssd1 vssd1 vccd1 vccd1 _6625_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7044_ _7044_/CLK _7044_/D vssd1 vssd1 vccd1 vccd1 _7044_/Q sky130_fd_sc_hd__dfxtp_1
X_4256_ _4256_/A vssd1 vssd1 vccd1 vccd1 _6655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5816__505 _5816__505/A vssd1 vssd1 vccd1 vccd1 _6811_/CLK sky130_fd_sc_hd__inv_2
X_4187_ _4202_/S vssd1 vssd1 vccd1 vccd1 _4196_/S sky130_fd_sc_hd__buf_2
X_3207_ _6731_/Q vssd1 vssd1 vccd1 vccd1 _5258_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6828_ _6828_/CLK _6828_/D vssd1 vssd1 vccd1 vccd1 _6828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6759_ _6759_/CLK _6759_/D vssd1 vssd1 vccd1 vccd1 _6759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5201__255 _5202__256/A vssd1 vssd1 vccd1 vccd1 _6537_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4110_/A vssd1 vssd1 vccd1 vccd1 _6720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5090_ _5090_/A vssd1 vssd1 vccd1 vccd1 _6461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4041_ _3623_/A _4040_/Y _4404_/B _4049_/B _4037_/X vssd1 vssd1 vccd1 vccd1 _6739_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5992_ _6002_/A _5992_/B vssd1 vssd1 vccd1 vccd1 _5993_/A sky130_fd_sc_hd__and2_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _6509_/Q _6443_/Q _6541_/Q _6693_/Q _4778_/X _4914_/X vssd1 vssd1 vccd1 vccd1
+ _4944_/B sky130_fd_sc_hd__mux4_2
XFILLER_24_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2741_ _5529_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2741_/X sky130_fd_sc_hd__clkbuf_16
X_4874_ _6482_/Q _6554_/Q _7043_/Q _6974_/Q _4957_/S _4914_/A vssd1 vssd1 vccd1 vccd1
+ _4874_/X sky130_fd_sc_hd__mux4_1
X_6613_ _6613_/CLK _6613_/D vssd1 vssd1 vccd1 vccd1 _6613_/Q sky130_fd_sc_hd__dfxtp_1
X_3825_ _6820_/Q _3620_/X _3825_/S vssd1 vssd1 vccd1 vccd1 _3826_/A sky130_fd_sc_hd__mux2_1
X_6544_ _6544_/CLK _6544_/D vssd1 vssd1 vccd1 vccd1 _6544_/Q sky130_fd_sc_hd__dfxtp_1
X_3756_ _6847_/Q _3611_/X _3756_/S vssd1 vssd1 vccd1 vccd1 _3757_/A sky130_fd_sc_hd__mux2_1
X_6475_ _6475_/CLK _6475_/D vssd1 vssd1 vccd1 vccd1 _6475_/Q sky130_fd_sc_hd__dfxtp_1
X_3687_ _4014_/A vssd1 vssd1 vccd1 vccd1 _3687_/X sky130_fd_sc_hd__clkbuf_4
X_5426_ _6580_/Q _5321_/X _5425_/X _5406_/X vssd1 vssd1 vccd1 vccd1 _6580_/D sky130_fd_sc_hd__o211a_1
XFILLER_99_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5357_ _5355_/B _5356_/X _5394_/S vssd1 vssd1 vccd1 vccd1 _5357_/Y sky130_fd_sc_hd__o21ai_1
XINSDIODE2_4 _5774_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3155_ _6343_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3155_/X sky130_fd_sc_hd__clkbuf_16
X_4308_ _3782_/X _6632_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__mux2_1
X_5288_ _5302_/A vssd1 vssd1 vccd1 vccd1 _5435_/B sky130_fd_sc_hd__clkbuf_1
X_7027_ _7030_/CLK _7027_/D vssd1 vssd1 vccd1 vccd1 _7027_/Q sky130_fd_sc_hd__dfxtp_1
X_4239_ _3788_/X _6662_/Q _4239_/S vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6371__53 _6372__54/A vssd1 vssd1 vccd1 vccd1 _7073_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5199__254 _5199__254/A vssd1 vssd1 vccd1 vccd1 _6536_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5537__365 _5538__366/A vssd1 vssd1 vccd1 vccd1 _6655_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4590_ _4590_/A _4590_/B vssd1 vssd1 vccd1 vccd1 _4606_/S sky130_fd_sc_hd__nor2_2
XFILLER_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3610_ _3610_/A vssd1 vssd1 vccd1 vccd1 _6926_/D sky130_fd_sc_hd__clkbuf_1
X_3541_ _3541_/A vssd1 vssd1 vccd1 vccd1 _6954_/D sky130_fd_sc_hd__clkbuf_1
X_6260_ _6260_/A vssd1 vssd1 vccd1 vccd1 _7008_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3472_ _3372_/X _6983_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3473_/A sky130_fd_sc_hd__mux2_1
X_6191_ _6290_/A vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5073_ _5588_/S vssd1 vssd1 vccd1 vccd1 _5082_/S sky130_fd_sc_hd__clkbuf_2
X_4024_ _4023_/X _6754_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4025_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__2756_ clkbuf_0__2756_/X vssd1 vssd1 vccd1 vccd1 _5756_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5975_ _6877_/Q _5944_/X _5974_/Y _5953_/B vssd1 vssd1 vccd1 vccd1 _5976_/B sky130_fd_sc_hd__o2bb2a_1
X_4926_ _6476_/Q _6628_/Q _7061_/Q _6786_/Q _4719_/X _4772_/S vssd1 vssd1 vccd1 vccd1
+ _4927_/B sky130_fd_sc_hd__mux4_1
X_4857_ _4883_/B vssd1 vssd1 vccd1 vccd1 _4857_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3808_ _3808_/A vssd1 vssd1 vccd1 vccd1 _6828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6527_ _6527_/CLK _6527_/D vssd1 vssd1 vccd1 vccd1 _6527_/Q sky130_fd_sc_hd__dfxtp_1
X_5746__451 _5747__452/A vssd1 vssd1 vccd1 vccd1 _6755_/CLK sky130_fd_sc_hd__inv_2
X_4788_ _4786_/X _4787_/X _4905_/A vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__mux2_1
X_3739_ _3739_/A vssd1 vssd1 vccd1 vccd1 _6855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6458_ _7079_/CLK _6458_/D vssd1 vssd1 vccd1 vccd1 _6458_/Q sky130_fd_sc_hd__dfxtp_1
X_6389_ _6389_/A _6389_/B vssd1 vssd1 vccd1 vccd1 _6390_/A sky130_fd_sc_hd__and2_1
X_5409_ _6676_/Q _6668_/Q _6660_/Q _6652_/Q _5263_/X _5264_/X vssd1 vssd1 vccd1 vccd1
+ _5409_/X sky130_fd_sc_hd__mux4_2
XFILLER_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5864__63 _5865__64/A vssd1 vssd1 vccd1 vccd1 _6849_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5829__515 _5831__517/A vssd1 vssd1 vccd1 vccd1 _6821_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6073__120 _6075__122/A vssd1 vssd1 vccd1 vccd1 _6928_/CLK sky130_fd_sc_hd__inv_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5691_ _5697_/A vssd1 vssd1 vccd1 vccd1 _5691_/X sky130_fd_sc_hd__buf_1
X_4711_ _6770_/Q vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4642_ _3868_/X _6478_/Q _4642_/S vssd1 vssd1 vccd1 vccd1 _4643_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5214__265 _5216__267/A vssd1 vssd1 vccd1 vccd1 _6547_/CLK sky130_fd_sc_hd__inv_2
X_4573_ _4588_/S vssd1 vssd1 vccd1 vccd1 _4582_/S sky130_fd_sc_hd__buf_2
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6312_ _7129_/A _6314_/B _6312_/C vssd1 vssd1 vccd1 vccd1 _6313_/A sky130_fd_sc_hd__and3_1
X_3524_ _4205_/A _3579_/A vssd1 vssd1 vccd1 vccd1 _3540_/S sky130_fd_sc_hd__nor2_2
X_6243_ _6250_/A _6249_/D vssd1 vssd1 vccd1 vccd1 _6243_/X sky130_fd_sc_hd__or2_1
X_3455_ _3455_/A vssd1 vssd1 vccd1 vccd1 _6989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6174_ _6174_/A _6174_/B vssd1 vssd1 vccd1 vccd1 _6175_/B sky130_fd_sc_hd__nand2_1
X_3386_ _3386_/A vssd1 vssd1 vccd1 vccd1 _7049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5056_ _5056_/A vssd1 vssd1 vccd1 vccd1 _6446_/D sky130_fd_sc_hd__clkbuf_1
X_4007_ _3705_/X _6759_/Q _4007_/S vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5958_ _6874_/Q _5944_/X _5957_/Y _5953_/B vssd1 vssd1 vccd1 vccd1 _5959_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__2739_ clkbuf_0__2739_/X vssd1 vssd1 vccd1 vccd1 _5519__351/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _4909_/A vssd1 vssd1 vccd1 vccd1 _4944_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5889_ _6883_/Q _5609_/Y _5610_/X _6885_/Q _5888_/X vssd1 vssd1 vccd1 vccd1 _5922_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6137__172 _6137__172/A vssd1 vssd1 vccd1 vccd1 _6980_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _6453_/Q _6454_/Q _3240_/C _4752_/B vssd1 vssd1 vccd1 vccd1 _5044_/B sky130_fd_sc_hd__nor4_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6930_ _6930_/CLK _6930_/D vssd1 vssd1 vccd1 vccd1 _6930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6861_ _6861_/CLK _6861_/D vssd1 vssd1 vccd1 vccd1 _6861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6792_ _6792_/CLK _6792_/D vssd1 vssd1 vccd1 vccd1 _6792_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__2524_ clkbuf_0__2524_/X vssd1 vssd1 vccd1 vccd1 _5199__254/A sky130_fd_sc_hd__clkbuf_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5674_ _6271_/A _6272_/B _6290_/A vssd1 vssd1 vccd1 vccd1 _5675_/A sky130_fd_sc_hd__and3b_1
Xclkbuf_1_1_0__2455_ clkbuf_0__2455_/X vssd1 vssd1 vccd1 vccd1 _5030_/A sky130_fd_sc_hd__clkbuf_4
X_4625_ _4625_/A vssd1 vssd1 vccd1 vccd1 _6486_/D sky130_fd_sc_hd__clkbuf_1
X_4556_ _6517_/Q _4009_/A _4562_/S vssd1 vssd1 vccd1 vccd1 _4557_/A sky130_fd_sc_hd__mux2_1
X_5034__183 _5035__184/A vssd1 vssd1 vccd1 vccd1 _6439_/CLK sky130_fd_sc_hd__inv_2
X_3507_ _3522_/S vssd1 vssd1 vccd1 vccd1 _3516_/S sky130_fd_sc_hd__buf_2
X_4487_ _6745_/Q vssd1 vssd1 vccd1 vccd1 _4487_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__3007_ clkbuf_0__3007_/X vssd1 vssd1 vccd1 vccd1 _6083__129/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0_0__2740_ clkbuf_0__2740_/X vssd1 vssd1 vccd1 vccd1 _5528__359/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6226_ _6226_/A vssd1 vssd1 vccd1 vccd1 _7001_/D sky130_fd_sc_hd__clkbuf_1
X_3438_ _4204_/A vssd1 vssd1 vccd1 vccd1 _4277_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6157_ _7009_/Q vssd1 vssd1 vccd1 vccd1 _6262_/A sky130_fd_sc_hd__inv_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3368_/X _7053_/Q _3381_/S vssd1 vssd1 vccd1 vccd1 _3370_/A sky130_fd_sc_hd__mux2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _6574_/Q _6575_/Q _6576_/Q _6577_/Q _6886_/Q _6887_/Q vssd1 vssd1 vccd1 vccd1
+ _5108_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5460__304 _5460__304/A vssd1 vssd1 vccd1 vccd1 _6594_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__2869_ clkbuf_0__2869_/X vssd1 vssd1 vccd1 vccd1 _5833__519/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5759__461 _5760__462/A vssd1 vssd1 vccd1 vccd1 _6765_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2532_ clkbuf_0__2532_/X vssd1 vssd1 vccd1 vccd1 _5560_/A sky130_fd_sc_hd__clkbuf_16
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4410_ _3254_/X _6587_/Q _4414_/S vssd1 vssd1 vccd1 vccd1 _4411_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5390_ _5388_/X _5389_/X _5410_/S vssd1 vssd1 vccd1 vccd1 _5390_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4341_ _4341_/A vssd1 vssd1 vccd1 vccd1 _6618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7060_ _7060_/CLK _7060_/D vssd1 vssd1 vccd1 vccd1 _7060_/Q sky130_fd_sc_hd__dfxtp_1
X_4272_ _4272_/A vssd1 vssd1 vccd1 vccd1 _6648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6011_ _5954_/B _6012_/B _6012_/D vssd1 vssd1 vccd1 vccd1 _6011_/X sky130_fd_sc_hd__and3b_1
X_3223_ _6736_/Q _6731_/Q vssd1 vssd1 vccd1 vccd1 _3223_/X sky130_fd_sc_hd__or2_1
XFILLER_94_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6913_ _6913_/CLK _6913_/D vssd1 vssd1 vccd1 vccd1 _6913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6086__130 _6088__132/A vssd1 vssd1 vccd1 vccd1 _6938_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6844_ _6844_/CLK _6844_/D vssd1 vssd1 vccd1 vccd1 _6844_/Q sky130_fd_sc_hd__dfxtp_1
X_3987_ _3982_/Y _4856_/A _3986_/X vssd1 vssd1 vccd1 vccd1 _3988_/B sky130_fd_sc_hd__o21ai_1
X_6775_ _6775_/CLK _6775_/D vssd1 vssd1 vccd1 vccd1 _6775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5726_ _7018_/Q _5734_/B vssd1 vssd1 vccd1 vccd1 _5727_/A sky130_fd_sc_hd__and2_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5657_ _5657_/A _5657_/B _5657_/C _5657_/D vssd1 vssd1 vccd1 vccd1 _5657_/X sky130_fd_sc_hd__or4_1
X_4608_ _4608_/A _4608_/B vssd1 vssd1 vccd1 vccd1 _4624_/S sky130_fd_sc_hd__or2_2
X_5588_ _6696_/Q _7159_/A _5588_/S vssd1 vssd1 vccd1 vccd1 _5589_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4539_ _4554_/S vssd1 vssd1 vccd1 vccd1 _4548_/S sky130_fd_sc_hd__buf_2
XFILLER_2_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6209_ _6216_/B _6216_/C _6249_/C _6217_/B vssd1 vssd1 vccd1 vccd1 _6210_/B sky130_fd_sc_hd__a31o_1
XFILLER_77_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5193__249 _5193__249/A vssd1 vssd1 vccd1 vccd1 _6531_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2867_ clkbuf_0__2867_/X vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4890_ _5918_/A _4763_/X _4695_/A vssd1 vssd1 vccd1 vccd1 _4890_/X sky130_fd_sc_hd__o21a_1
X_3910_ _6790_/Q _3614_/X _3914_/S vssd1 vssd1 vccd1 vccd1 _3911_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3841_ _6813_/Q _3617_/X _3843_/S vssd1 vssd1 vccd1 vccd1 _3842_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6560_ _6560_/CLK _6560_/D vssd1 vssd1 vccd1 vccd1 _6560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3772_ _3772_/A vssd1 vssd1 vccd1 vccd1 _6842_/D sky130_fd_sc_hd__clkbuf_1
X_5511_ _5523_/A vssd1 vssd1 vccd1 vccd1 _5511_/X sky130_fd_sc_hd__buf_1
X_6491_ _6491_/CLK _6491_/D vssd1 vssd1 vccd1 vccd1 _6491_/Q sky130_fd_sc_hd__dfxtp_1
X_5442_ _5334_/X _5435_/X _5437_/Y _5439_/X _5441_/Y vssd1 vssd1 vccd1 vccd1 _5442_/X
+ sky130_fd_sc_hd__o32a_2
X_5373_ _6602_/Q _6586_/Q _6840_/Q _6824_/Q _5329_/X _5330_/X vssd1 vssd1 vccd1 vccd1
+ _5373_/X sky130_fd_sc_hd__mux4_1
X_7112_ _7112_/A vssd1 vssd1 vccd1 vccd1 _7112_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4324_ _6625_/Q _3886_/X _4324_/S vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7043_ _7043_/CLK _7043_/D vssd1 vssd1 vccd1 vccd1 _7043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4255_ _3785_/X _6655_/Q _4257_/S vssd1 vssd1 vccd1 vccd1 _4256_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4186_ _4186_/A _4386_/B vssd1 vssd1 vccd1 vccd1 _4202_/S sky130_fd_sc_hd__nor2_2
X_3206_ _3361_/A vssd1 vssd1 vccd1 vccd1 _4048_/A sky130_fd_sc_hd__inv_2
XFILLER_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6827_ _6827_/CLK _6827_/D vssd1 vssd1 vccd1 vccd1 _6827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6758_ _6758_/CLK _6758_/D vssd1 vssd1 vccd1 vccd1 _6758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6689_ _6689_/CLK _6689_/D vssd1 vssd1 vccd1 vccd1 _6689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7011_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_4040_ _4040_/A _4049_/B vssd1 vssd1 vccd1 vccd1 _4040_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5991_ _5994_/B _5966_/X _5990_/X _5970_/X vssd1 vssd1 vccd1 vccd1 _5992_/B sky130_fd_sc_hd__a22o_1
X_5473__314 _5473__314/A vssd1 vssd1 vccd1 vccd1 _6604_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _4888_/X input31/X _4695_/X _4941_/X vssd1 vssd1 vccd1 vccd1 _4942_/X sky130_fd_sc_hd__a22o_2
XFILLER_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2740_ _5523_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2740_/X sky130_fd_sc_hd__clkbuf_16
X_4873_ _6902_/Q _6562_/Q _6910_/Q _6490_/Q _4906_/A _4898_/A vssd1 vssd1 vccd1 vccd1
+ _4873_/X sky130_fd_sc_hd__mux4_1
X_6612_ _6612_/CLK _6612_/D vssd1 vssd1 vccd1 vccd1 _6612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3824_ _3824_/A vssd1 vssd1 vccd1 vccd1 _6821_/D sky130_fd_sc_hd__clkbuf_1
X_6543_ _6543_/CLK _6543_/D vssd1 vssd1 vccd1 vccd1 _6543_/Q sky130_fd_sc_hd__dfxtp_1
X_3755_ _3755_/A vssd1 vssd1 vccd1 vccd1 _6848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3686_ _3686_/A vssd1 vssd1 vccd1 vccd1 _6896_/D sky130_fd_sc_hd__clkbuf_1
X_6474_ _6474_/CLK _6474_/D vssd1 vssd1 vccd1 vccd1 _6474_/Q sky130_fd_sc_hd__dfxtp_1
X_5425_ _5324_/X _5414_/X _5424_/Y vssd1 vssd1 vccd1 vccd1 _5425_/X sky130_fd_sc_hd__a21o_1
XFILLER_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5356_ _6957_/Q _6941_/Q _7066_/Q _6933_/Q _5282_/X _4083_/X vssd1 vssd1 vccd1 vccd1
+ _5356_/X sky130_fd_sc_hd__mux4_2
XINSDIODE2_5 _4009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5779__475 _5780__476/A vssd1 vssd1 vccd1 vccd1 _6781_/CLK sky130_fd_sc_hd__inv_2
X_4307_ _4307_/A vssd1 vssd1 vccd1 vccd1 _6633_/D sky130_fd_sc_hd__clkbuf_1
X_5287_ _5285_/X _5432_/S vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__and2b_1
Xclkbuf_0__3154_ _6342_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3154_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_101_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7026_ _7030_/CLK _7026_/D vssd1 vssd1 vccd1 vccd1 _7026_/Q sky130_fd_sc_hd__dfxtp_1
X_4238_ _4238_/A vssd1 vssd1 vccd1 vccd1 _6663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4169_ _4184_/S vssd1 vssd1 vccd1 vccd1 _4178_/S sky130_fd_sc_hd__buf_2
XFILLER_83_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6131__167 _6132__168/A vssd1 vssd1 vccd1 vccd1 _6975_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2869_ _5828_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2869_/X sky130_fd_sc_hd__clkbuf_16
X_6356__40 _6358__42/A vssd1 vssd1 vccd1 vccd1 _7060_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3540_ _6954_/Q _3462_/X _3540_/S vssd1 vssd1 vccd1 vccd1 _3541_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3471_ _3471_/A vssd1 vssd1 vccd1 vccd1 _6984_/D sky130_fd_sc_hd__clkbuf_1
X_6190_ _6245_/B _6187_/B _6187_/C _6245_/A vssd1 vssd1 vccd1 vccd1 _6190_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5072_ _5072_/A vssd1 vssd1 vccd1 vccd1 _6453_/D sky130_fd_sc_hd__clkbuf_1
X_4023_ _4023_/A vssd1 vssd1 vccd1 vccd1 _4023_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2755_ clkbuf_0__2755_/X vssd1 vssd1 vccd1 vccd1 _5596__409/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5974_ _6877_/Q _5978_/C vssd1 vssd1 vccd1 vccd1 _5974_/Y sky130_fd_sc_hd__xnor2_1
X_4925_ _4927_/A _4924_/X _4802_/X vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4856_ _4856_/A _4856_/B vssd1 vssd1 vccd1 vccd1 _4856_/Y sky130_fd_sc_hd__nor2_2
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3807_ _3705_/X _6828_/Q _3807_/S vssd1 vssd1 vccd1 vccd1 _3808_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6526_ _6526_/CLK _6526_/D vssd1 vssd1 vccd1 vccd1 _6526_/Q sky130_fd_sc_hd__dfxtp_1
X_4787_ _6503_/Q _6437_/Q _6535_/Q _6687_/Q _4900_/S _4728_/X vssd1 vssd1 vccd1 vccd1
+ _4787_/X sky130_fd_sc_hd__mux4_2
X_5150__214 _5150__214/A vssd1 vssd1 vccd1 vccd1 _6496_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3738_ _3696_/X _6855_/Q _3738_/S vssd1 vssd1 vccd1 vccd1 _3739_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3669_ _3669_/A vssd1 vssd1 vccd1 vccd1 _6903_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6457_ _7079_/CLK _6457_/D vssd1 vssd1 vccd1 vccd1 _6457_/Q sky130_fd_sc_hd__dfxtp_1
X_6388_ _7139_/A _6155_/A _6401_/S vssd1 vssd1 vccd1 vccd1 _6389_/B sky130_fd_sc_hd__mux2_1
X_5408_ _7077_/Q _6703_/Q _6572_/Q _6850_/Q _5257_/X _5254_/X vssd1 vssd1 vccd1 vccd1
+ _5408_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5339_ _6948_/Q _6680_/Q _6592_/Q _6814_/Q _5337_/X _5338_/X vssd1 vssd1 vccd1 vccd1
+ _5340_/B sky130_fd_sc_hd__mux4_1
XFILLER_48_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7009_ _7011_/CLK _7009_/D vssd1 vssd1 vccd1 vccd1 _7009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6026__83 _6027__84/A vssd1 vssd1 vccd1 vccd1 _6890_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5543__370 _5544__371/A vssd1 vssd1 vccd1 vccd1 _6660_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4710_ _6759_/Q _6751_/Q _6714_/Q _6706_/Q _4891_/B _4709_/X vssd1 vssd1 vccd1 vccd1
+ _4710_/X sky130_fd_sc_hd__mux4_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4641_ _4641_/A vssd1 vssd1 vccd1 vccd1 _6479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4572_ _4572_/A _4662_/B vssd1 vssd1 vccd1 vccd1 _4588_/S sky130_fd_sc_hd__or2_2
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6311_ _6311_/A vssd1 vssd1 vccd1 vccd1 _7026_/D sky130_fd_sc_hd__clkbuf_1
X_3523_ _3523_/A vssd1 vssd1 vccd1 vccd1 _6962_/D sky130_fd_sc_hd__clkbuf_1
X_6242_ _7001_/Q _6250_/C _6250_/D vssd1 vssd1 vccd1 vccd1 _6249_/D sky130_fd_sc_hd__and3_1
X_6350__35 _6352__37/A vssd1 vssd1 vccd1 vccd1 _7055_/CLK sky130_fd_sc_hd__inv_2
X_3454_ _6989_/Q _3453_/X _3454_/S vssd1 vssd1 vccd1 vccd1 _3455_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6173_ _6173_/A _6217_/B vssd1 vssd1 vccd1 vccd1 _6174_/B sky130_fd_sc_hd__xnor2_1
X_3385_ _3384_/X _7049_/Q _3393_/S vssd1 vssd1 vccd1 vccd1 _3386_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5055_ _4795_/A _7100_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5056_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4006_ _4006_/A vssd1 vssd1 vccd1 vccd1 _6760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _6874_/Q _5961_/C vssd1 vssd1 vccd1 vccd1 _5957_/Y sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1_0__2738_ clkbuf_0__2738_/X vssd1 vssd1 vccd1 vccd1 _5516__349/A sky130_fd_sc_hd__clkbuf_4
X_4908_ _4927_/A _4908_/B vssd1 vssd1 vccd1 vccd1 _4908_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5888_ _6885_/Q _6884_/Q _5888_/C vssd1 vssd1 vccd1 vccd1 _5888_/X sky130_fd_sc_hd__and3b_1
X_4839_ _6892_/Q _6521_/Q _4876_/A vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6509_ _6509_/CLK _6509_/D vssd1 vssd1 vccd1 vccd1 _6509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5835__520 _5836__521/A vssd1 vssd1 vccd1 vccd1 _6826_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5220__270 _5223__273/A vssd1 vssd1 vccd1 vccd1 _6552_/CLK sky130_fd_sc_hd__inv_2
X_6860_ _6860_/CLK _6860_/D vssd1 vssd1 vccd1 vccd1 _6860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6791_ _6791_/CLK _6791_/D vssd1 vssd1 vccd1 vccd1 _6791_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__2523_ clkbuf_0__2523_/X vssd1 vssd1 vccd1 vccd1 _5190__246/A sky130_fd_sc_hd__clkbuf_4
X_5673_ _7125_/A _3242_/X _6433_/A vssd1 vssd1 vccd1 vccd1 _6290_/A sky130_fd_sc_hd__a21oi_4
X_4624_ _3868_/X _6486_/Q _4624_/S vssd1 vssd1 vccd1 vccd1 _4625_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4555_ _4555_/A vssd1 vssd1 vccd1 vccd1 _6518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3506_ _3827_/A _3898_/B vssd1 vssd1 vccd1 vccd1 _3522_/S sky130_fd_sc_hd__nor2_2
X_4486_ _4486_/A vssd1 vssd1 vccd1 vccd1 _6547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__3006_ clkbuf_0__3006_/X vssd1 vssd1 vccd1 vccd1 _6077__124/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6225_ _6228_/B _6225_/B _6229_/C vssd1 vssd1 vccd1 vccd1 _6226_/A sky130_fd_sc_hd__and3b_1
X_3437_ _3764_/A vssd1 vssd1 vccd1 vccd1 _3437_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6156_ _6999_/Q vssd1 vssd1 vccd1 vccd1 _6156_/Y sky130_fd_sc_hd__inv_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3368_/X sky130_fd_sc_hd__buf_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5924_/D vssd1 vssd1 vccd1 vccd1 _5929_/A sky130_fd_sc_hd__inv_2
X_3299_ _6774_/Q vssd1 vssd1 vccd1 vccd1 _4167_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5121__190 _5125__194/A vssd1 vssd1 vccd1 vccd1 _6472_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3153_ clkbuf_0__3153_/X vssd1 vssd1 vccd1 vccd1 _6341__29/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6989_ _6989_/CLK _6989_/D vssd1 vssd1 vccd1 vccd1 _6989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2868_ clkbuf_0__2868_/X vssd1 vssd1 vccd1 vccd1 _5825__512/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4340_ _3776_/X _6618_/Q _4342_/S vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4271_ _6648_/Q _4158_/X _4275_/S vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6010_ _6012_/D _6005_/X _6009_/Y _5976_/A vssd1 vssd1 vccd1 vccd1 _6884_/D sky130_fd_sc_hd__a211oi_1
X_3222_ _6736_/Q _5258_/A vssd1 vssd1 vccd1 vccd1 _3222_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6912_ _6912_/CLK _6912_/D vssd1 vssd1 vccd1 vccd1 _6912_/Q sky130_fd_sc_hd__dfxtp_1
X_6843_ _6843_/CLK _6843_/D vssd1 vssd1 vccd1 vccd1 _6843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3986_ _3986_/A vssd1 vssd1 vccd1 vccd1 _3986_/X sky130_fd_sc_hd__buf_2
X_6774_ _6774_/CLK _6774_/D vssd1 vssd1 vccd1 vccd1 _6774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5725_ _5774_/C vssd1 vssd1 vccd1 vccd1 _5734_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5656_ _5890_/B _6178_/A vssd1 vssd1 vccd1 vccd1 _5657_/D sky130_fd_sc_hd__xor2_1
XFILLER_31_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4607_ _4607_/A vssd1 vssd1 vccd1 vccd1 _6494_/D sky130_fd_sc_hd__clkbuf_1
X_5587_ _5587_/A vssd1 vssd1 vccd1 vccd1 _6695_/D sky130_fd_sc_hd__clkbuf_1
X_4538_ _4662_/A _4590_/B vssd1 vssd1 vccd1 vccd1 _4554_/S sky130_fd_sc_hd__or2_2
XFILLER_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4469_ _4469_/A vssd1 vssd1 vccd1 vccd1 _6553_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6208_ _6254_/C vssd1 vssd1 vccd1 vccd1 _6249_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5227__276 _5230__279/A vssd1 vssd1 vccd1 vccd1 _6558_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2866_ clkbuf_0__2866_/X vssd1 vssd1 vccd1 vccd1 _5816__505/A sky130_fd_sc_hd__clkbuf_16
X_5128__196 _5130__198/A vssd1 vssd1 vccd1 vccd1 _6478_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3840_ _3840_/A vssd1 vssd1 vccd1 vccd1 _6814_/D sky130_fd_sc_hd__clkbuf_1
X_3771_ _3770_/X _6842_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3772_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6490_ _6490_/CLK _6490_/D vssd1 vssd1 vccd1 vccd1 _6490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5441_ _5351_/B _5440_/X _5334_/A vssd1 vssd1 vccd1 vccd1 _5441_/Y sky130_fd_sc_hd__o21ai_1
X_5372_ _6642_/Q _6634_/Q _6618_/Q _6610_/Q _4083_/A _5264_/X vssd1 vssd1 vccd1 vccd1
+ _5372_/X sky130_fd_sc_hd__mux4_1
X_7111_ _7111_/A vssd1 vssd1 vccd1 vccd1 _7111_/X sky130_fd_sc_hd__clkbuf_1
X_4323_ _4323_/A vssd1 vssd1 vccd1 vccd1 _6626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7042_ _7042_/CLK _7042_/D vssd1 vssd1 vccd1 vccd1 _7042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4254_ _4254_/A vssd1 vssd1 vccd1 vccd1 _6656_/D sky130_fd_sc_hd__clkbuf_1
X_4185_ _4185_/A vssd1 vssd1 vccd1 vccd1 _6686_/D sky130_fd_sc_hd__clkbuf_1
X_3205_ _6735_/Q vssd1 vssd1 vccd1 vccd1 _4051_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6826_ _6826_/CLK _6826_/D vssd1 vssd1 vccd1 vccd1 _6826_/Q sky130_fd_sc_hd__dfxtp_1
X_6757_ _6757_/CLK _6757_/D vssd1 vssd1 vccd1 vccd1 _6757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3969_ _3974_/A _3978_/B vssd1 vssd1 vccd1 vccd1 _3975_/B sky130_fd_sc_hd__nand2_1
X_6688_ _6688_/CLK _6688_/D vssd1 vssd1 vccd1 vccd1 _6688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5639_ _7091_/Q _7000_/Q vssd1 vssd1 vccd1 vccd1 _6178_/B sky130_fd_sc_hd__xor2_1
XFILLER_105_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5507__341 _5508__342/A vssd1 vssd1 vccd1 vccd1 _6631_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5990_ _5994_/B _5994_/C vssd1 vssd1 vccd1 vccd1 _5990_/X sky130_fd_sc_hd__xor2_1
X_4941_ _4856_/Y _4930_/X _4940_/X _4987_/C _7090_/Q vssd1 vssd1 vccd1 vccd1 _4941_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4872_ _4722_/X _4863_/X _4865_/X _4871_/X _3951_/Y vssd1 vssd1 vccd1 vccd1 _4872_/X
+ sky130_fd_sc_hd__a311o_2
X_6611_ _6611_/CLK _6611_/D vssd1 vssd1 vccd1 vccd1 _6611_/Q sky130_fd_sc_hd__dfxtp_1
X_3823_ _6821_/Q _3617_/X _3825_/S vssd1 vssd1 vccd1 vccd1 _3824_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6542_ _6542_/CLK _6542_/D vssd1 vssd1 vccd1 vccd1 _6542_/Q sky130_fd_sc_hd__dfxtp_1
X_3754_ _6848_/Q _3608_/X _3756_/S vssd1 vssd1 vccd1 vccd1 _3755_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3685_ _3680_/X _6896_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3686_/A sky130_fd_sc_hd__mux2_1
X_6473_ _6473_/CLK _6473_/D vssd1 vssd1 vccd1 vccd1 _6473_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput200 _5019_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[31] sky130_fd_sc_hd__buf_2
X_5424_ _5324_/A _5423_/X _5321_/A vssd1 vssd1 vccd1 vccd1 _5424_/Y sky130_fd_sc_hd__o21ai_1
X_5355_ _5354_/X _5355_/B vssd1 vssd1 vccd1 vccd1 _5355_/X sky130_fd_sc_hd__and2b_1
XINSDIODE2_6 _4014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5876__73 _5876__73/A vssd1 vssd1 vccd1 vccd1 _6859_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__3153_ _6336_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3153_/X sky130_fd_sc_hd__clkbuf_16
X_4306_ _3779_/X _6633_/Q _4306_/S vssd1 vssd1 vccd1 vccd1 _4307_/A sky130_fd_sc_hd__mux2_1
X_5286_ _5286_/A vssd1 vssd1 vccd1 vccd1 _5432_/S sky130_fd_sc_hd__buf_4
XFILLER_87_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7025_ _7030_/CLK _7025_/D vssd1 vssd1 vccd1 vccd1 _7025_/Q sky130_fd_sc_hd__dfxtp_1
X_4237_ _3785_/X _6663_/Q _4239_/S vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4168_ _4168_/A _4662_/B vssd1 vssd1 vccd1 vccd1 _4184_/S sky130_fd_sc_hd__or2_2
XFILLER_83_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4099_ _4026_/X _6724_/Q _4103_/S vssd1 vssd1 vccd1 vccd1 _4100_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6038__92 _6038__92/A vssd1 vssd1 vccd1 vccd1 _6900_/CLK sky130_fd_sc_hd__inv_2
X_6809_ _6809_/CLK _6809_/D vssd1 vssd1 vccd1 vccd1 _6809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2868_ _5822_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2868_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6099__141 _6099__141/A vssd1 vssd1 vccd1 vccd1 _6949_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3470_ _3368_/X _6984_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3471_/A sky130_fd_sc_hd__mux2_1
X_5698__430 _5702__434/A vssd1 vssd1 vccd1 vccd1 _6724_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5071_ _6453_/Q _7107_/A _5071_/S vssd1 vssd1 vccd1 vccd1 _5072_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4022_ _4022_/A vssd1 vssd1 vccd1 vccd1 _6755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5973_ _5973_/A vssd1 vssd1 vccd1 vccd1 _6876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4924_ _6858_/Q _6834_/Q _6810_/Q _6802_/Q _4923_/X _4892_/X vssd1 vssd1 vccd1 vccd1
+ _4924_/X sky130_fd_sc_hd__mux4_2
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4855_ _4722_/X _4848_/X _4854_/X _3951_/Y vssd1 vssd1 vccd1 vccd1 _4855_/X sky130_fd_sc_hd__a211o_1
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4786_ _6853_/Q _6829_/Q _6805_/Q _6797_/Q _4900_/S _4728_/X vssd1 vssd1 vccd1 vccd1
+ _4786_/X sky130_fd_sc_hd__mux4_1
X_3806_ _3806_/A vssd1 vssd1 vccd1 vccd1 _6829_/D sky130_fd_sc_hd__clkbuf_1
X_6525_ _6525_/CLK _6525_/D vssd1 vssd1 vccd1 vccd1 _6525_/Q sky130_fd_sc_hd__dfxtp_1
X_3737_ _3737_/A vssd1 vssd1 vccd1 vccd1 _6856_/D sky130_fd_sc_hd__clkbuf_1
X_5785__480 _5786__481/A vssd1 vssd1 vccd1 vccd1 _6786_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5707__437 _5709__439/A vssd1 vssd1 vccd1 vccd1 _6731_/CLK sky130_fd_sc_hd__inv_2
X_3668_ _3333_/X _6903_/Q _3672_/S vssd1 vssd1 vccd1 vccd1 _3669_/A sky130_fd_sc_hd__mux2_1
X_6456_ _7089_/CLK _6456_/D vssd1 vssd1 vccd1 vccd1 _6456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6387_ _6387_/A vssd1 vssd1 vccd1 vccd1 _7081_/D sky130_fd_sc_hd__clkbuf_1
X_3599_ _3621_/S vssd1 vssd1 vccd1 vccd1 _3612_/S sky130_fd_sc_hd__clkbuf_2
X_5407_ _6579_/Q _5321_/X _5405_/X _5406_/X vssd1 vssd1 vccd1 vccd1 _6579_/D sky130_fd_sc_hd__o211a_1
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5338_ _5338_/A vssd1 vssd1 vccd1 vccd1 _5338_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7008_ _7008_/CLK _7008_/D vssd1 vssd1 vccd1 vccd1 _7008_/Q sky130_fd_sc_hd__dfxtp_1
X_5269_ _6598_/Q _6582_/Q _6836_/Q _6820_/Q _5266_/X _5268_/X vssd1 vssd1 vccd1 vccd1
+ _5269_/X sky130_fd_sc_hd__mux4_2
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5753__457 _5755__459/A vssd1 vssd1 vccd1 vccd1 _6761_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5246__290 _5448__294/A vssd1 vssd1 vccd1 vccd1 _6572_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5870__68 _5870__68/A vssd1 vssd1 vccd1 vccd1 _6854_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6080__126 _6082__128/A vssd1 vssd1 vccd1 vccd1 _6934_/CLK sky130_fd_sc_hd__inv_2
X_4640_ _3865_/X _6479_/Q _4642_/S vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4571_ _4571_/A vssd1 vssd1 vccd1 vccd1 _6510_/D sky130_fd_sc_hd__clkbuf_1
X_6310_ _7128_/A _6314_/B _6312_/C vssd1 vssd1 vccd1 vccd1 _6311_/A sky130_fd_sc_hd__and3_1
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3522_ _6962_/Q _3462_/X _3522_/S vssd1 vssd1 vccd1 vccd1 _3523_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6241_ _7004_/Q _6241_/B _6241_/C vssd1 vssd1 vccd1 vccd1 _6250_/D sky130_fd_sc_hd__and3_1
X_3453_ _3779_/A vssd1 vssd1 vccd1 vccd1 _3453_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3022_ clkbuf_0__3022_/X vssd1 vssd1 vccd1 vccd1 _6154__10/A sky130_fd_sc_hd__clkbuf_4
X_6172_ _6172_/A _6172_/B _6172_/C _6171_/X vssd1 vssd1 vccd1 vccd1 _6172_/X sky130_fd_sc_hd__or4b_1
X_3384_ _3782_/A vssd1 vssd1 vccd1 vccd1 _3384_/X sky130_fd_sc_hd__buf_2
XFILLER_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5054_ _5054_/A vssd1 vssd1 vccd1 vccd1 _6445_/D sky130_fd_sc_hd__clkbuf_1
X_4005_ _3702_/X _6760_/Q _4007_/S vssd1 vssd1 vccd1 vccd1 _4006_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ _5953_/X _5954_/Y _5976_/A vssd1 vssd1 vccd1 vccd1 _6873_/D sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_1_0__2737_ clkbuf_0__2737_/X vssd1 vssd1 vccd1 vccd1 _5508__342/A sky130_fd_sc_hd__clkbuf_4
X_4907_ _6475_/Q _6627_/Q _7060_/Q _6785_/Q _4906_/X _3966_/X vssd1 vssd1 vccd1 vccd1
+ _4908_/B sky130_fd_sc_hd__mux4_2
X_4838_ _6497_/Q _6513_/Q _4898_/A vssd1 vssd1 vccd1 vccd1 _4838_/X sky130_fd_sc_hd__mux2_1
X_4769_ _6899_/Q _6559_/Q _6907_/Q _6487_/Q _4709_/X _4701_/X vssd1 vssd1 vccd1 vccd1
+ _4770_/B sky130_fd_sc_hd__mux4_1
X_6508_ _6508_/CLK _6508_/D vssd1 vssd1 vccd1 vccd1 _6508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6439_ _6439_/CLK _6439_/D vssd1 vssd1 vccd1 vccd1 _6439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6144__178 _6145__179/A vssd1 vssd1 vccd1 vccd1 _6986_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6790_ _6790_/CLK _6790_/D vssd1 vssd1 vccd1 vccd1 _6790_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__2522_ clkbuf_0__2522_/X vssd1 vssd1 vccd1 vccd1 _5186__243/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__2453_ clkbuf_0__2453_/X vssd1 vssd1 vccd1 vccd1 _5597_/A sky130_fd_sc_hd__clkbuf_4
X_5672_ _7014_/Q _7013_/Q _7012_/Q _6271_/B vssd1 vssd1 vccd1 vccd1 _6272_/B sky130_fd_sc_hd__and4_1
XFILLER_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4623_ _4623_/A vssd1 vssd1 vccd1 vccd1 _6487_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4554_ _4499_/X _6518_/Q _4554_/S vssd1 vssd1 vccd1 vccd1 _4555_/A sky130_fd_sc_hd__mux2_1
X_6323__14 _6323__14/A vssd1 vssd1 vccd1 vccd1 _7034_/CLK sky130_fd_sc_hd__inv_2
X_3505_ _4350_/A vssd1 vssd1 vccd1 vccd1 _3827_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4485_ _4484_/X _6547_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6224_ _7001_/Q _6224_/B vssd1 vssd1 vccd1 vccd1 _6225_/B sky130_fd_sc_hd__or2_1
Xclkbuf_1_1_0__3005_ clkbuf_0__3005_/X vssd1 vssd1 vccd1 vccd1 _6069__117/A sky130_fd_sc_hd__clkbuf_4
X_3436_ _3436_/A vssd1 vssd1 vccd1 vccd1 _7031_/D sky130_fd_sc_hd__clkbuf_1
X_6155_ _6155_/A vssd1 vssd1 vccd1 vccd1 _6155_/Y sky130_fd_sc_hd__inv_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _7029_/Q vssd1 vssd1 vccd1 vccd1 _3770_/A sky130_fd_sc_hd__clkbuf_4
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _6013_/A vssd1 vssd1 vccd1 vccd1 _5972_/A sky130_fd_sc_hd__clkbuf_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3298_ _4167_/A vssd1 vssd1 vccd1 vccd1 _3990_/B sky130_fd_sc_hd__clkbuf_4
X_5037_ _5037_/A vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__buf_1
XFILLER_45_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3152_ clkbuf_0__3152_/X vssd1 vssd1 vccd1 vccd1 _6334__23/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6988_ _6988_/CLK _6988_/D vssd1 vssd1 vccd1 vccd1 _6988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5939_ _5945_/C _5936_/X _5938_/X _5406_/X vssd1 vssd1 vccd1 vccd1 _6870_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5798__490 _5799__491/A vssd1 vssd1 vccd1 vccd1 _6796_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput100 wbs_data_i[9] vssd1 vssd1 vccd1 vccd1 _7134_/A sky130_fd_sc_hd__buf_4
XFILLER_103_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5501__336 _5502__337/A vssd1 vssd1 vccd1 vccd1 _6626_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5766__467 _5766__467/A vssd1 vssd1 vccd1 vccd1 _6771_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A vssd1 vssd1 vccd1 vccd1 _6649_/D sky130_fd_sc_hd__clkbuf_1
X_3221_ _3221_/A _3221_/B vssd1 vssd1 vccd1 vccd1 _4068_/B sky130_fd_sc_hd__or2_1
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6911_ _6911_/CLK _6911_/D vssd1 vssd1 vccd1 vccd1 _6911_/Q sky130_fd_sc_hd__dfxtp_1
X_6842_ _6842_/CLK _6842_/D vssd1 vssd1 vccd1 vccd1 _6842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5556__381 _5557__382/A vssd1 vssd1 vccd1 vccd1 _6671_/CLK sky130_fd_sc_hd__inv_2
XFILLER_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3985_ _4851_/S vssd1 vssd1 vccd1 vccd1 _3986_/A sky130_fd_sc_hd__clkinv_2
X_6773_ _6773_/CLK _6773_/D vssd1 vssd1 vccd1 vccd1 _6773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5724_ _5724_/A vssd1 vssd1 vccd1 vccd1 _6743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5655_ _5663_/A _7004_/Q vssd1 vssd1 vccd1 vccd1 _6178_/A sky130_fd_sc_hd__xor2_1
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4606_ _6494_/Q _4032_/A _4606_/S vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__mux2_1
X_5586_ _6695_/Q _7158_/A _5586_/S vssd1 vssd1 vccd1 vccd1 _5587_/A sky130_fd_sc_hd__mux2_1
X_4537_ _4537_/A vssd1 vssd1 vccd1 vccd1 _6526_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4468_ _4023_/X _6553_/Q _4468_/S vssd1 vssd1 vccd1 vccd1 _4469_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6093__136 _6094__137/A vssd1 vssd1 vccd1 vccd1 _6944_/CLK sky130_fd_sc_hd__inv_2
X_6207_ _6217_/B _6216_/B _6207_/C vssd1 vssd1 vccd1 vccd1 _6213_/B sky130_fd_sc_hd__and3_1
XFILLER_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3419_ _3623_/A _4040_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _3435_/S sky130_fd_sc_hd__or3_4
X_4399_ _4399_/A vssd1 vssd1 vccd1 vccd1 _6592_/D sky130_fd_sc_hd__clkbuf_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5692__425 _5694__427/A vssd1 vssd1 vccd1 vccd1 _6719_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3770_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3770_/X sky130_fd_sc_hd__buf_2
X_5848__531 _5849__532/A vssd1 vssd1 vccd1 vccd1 _6837_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5440_ _6961_/Q _6945_/Q _7070_/Q _6937_/Q _5266_/X _5268_/X vssd1 vssd1 vccd1 vccd1
+ _5440_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5371_ _5369_/X _5370_/X _5410_/S vssd1 vssd1 vccd1 vccd1 _5371_/X sky130_fd_sc_hd__mux2_1
X_7110_ _7110_/A vssd1 vssd1 vccd1 vccd1 _7110_/X sky130_fd_sc_hd__clkbuf_1
X_4322_ _6626_/Q _3883_/X _4324_/S vssd1 vssd1 vccd1 vccd1 _4323_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7041_ _7041_/CLK _7041_/D vssd1 vssd1 vccd1 vccd1 _7041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4253_ _3782_/X _6656_/Q _4257_/S vssd1 vssd1 vccd1 vccd1 _4254_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3204_ _6736_/Q vssd1 vssd1 vccd1 vccd1 _3361_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4184_ _4032_/X _6686_/Q _4184_/S vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
X_6825_ _6825_/CLK _6825_/D vssd1 vssd1 vccd1 vccd1 _6825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6756_ _6756_/CLK _6756_/D vssd1 vssd1 vccd1 vccd1 _6756_/Q sky130_fd_sc_hd__dfxtp_1
X_3968_ _3968_/A _3977_/A _3977_/B vssd1 vssd1 vccd1 vccd1 _3978_/B sky130_fd_sc_hd__and3_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6368__50 _6370__52/A vssd1 vssd1 vccd1 vccd1 _7070_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6687_ _6687_/CLK _6687_/D vssd1 vssd1 vccd1 vccd1 _6687_/Q sky130_fd_sc_hd__dfxtp_1
X_3899_ _3914_/S vssd1 vssd1 vccd1 vccd1 _3908_/S sky130_fd_sc_hd__buf_2
X_5233__281 _5236__284/A vssd1 vssd1 vccd1 vccd1 _6563_/CLK sky130_fd_sc_hd__inv_2
X_5638_ _6998_/Q _5906_/B _5906_/C vssd1 vssd1 vccd1 vccd1 _5638_/Y sky130_fd_sc_hd__nand3b_1
X_6101__143 _6102__144/A vssd1 vssd1 vccd1 vccd1 _6951_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240__285 _5242__287/A vssd1 vssd1 vccd1 vccd1 _6567_/CLK sky130_fd_sc_hd__inv_2
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5700__432 _5701__433/A vssd1 vssd1 vccd1 vccd1 _6726_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4940_ _4726_/X _4933_/X _4939_/X _3971_/X vssd1 vssd1 vccd1 vccd1 _4940_/X sky130_fd_sc_hd__a211o_1
XFILLER_91_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4871_ _4909_/A _4866_/X _4870_/X _3953_/A vssd1 vssd1 vccd1 vccd1 _4871_/X sky130_fd_sc_hd__o211a_1
X_6610_ _6610_/CLK _6610_/D vssd1 vssd1 vccd1 vccd1 _6610_/Q sky130_fd_sc_hd__dfxtp_1
X_3822_ _3822_/A vssd1 vssd1 vccd1 vccd1 _6822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6541_ _6541_/CLK _6541_/D vssd1 vssd1 vccd1 vccd1 _6541_/Q sky130_fd_sc_hd__dfxtp_1
X_3753_ _3753_/A vssd1 vssd1 vccd1 vccd1 _6849_/D sky130_fd_sc_hd__clkbuf_1
X_3684_ _3706_/S vssd1 vssd1 vccd1 vccd1 _3697_/S sky130_fd_sc_hd__clkbuf_2
X_6472_ _6472_/CLK _6472_/D vssd1 vssd1 vccd1 vccd1 _6472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput201 _4861_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[3] sky130_fd_sc_hd__buf_2
X_5423_ _5334_/X _5416_/X _5418_/Y _5420_/X _5422_/Y vssd1 vssd1 vccd1 vccd1 _5423_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_114_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5354_ _6925_/Q _6917_/Q _7034_/Q _7050_/Q _5281_/X _5282_/X vssd1 vssd1 vccd1 vccd1
+ _5354_/X sky130_fd_sc_hd__mux4_2
XFILLER_114_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4305_ _4305_/A vssd1 vssd1 vccd1 vccd1 _6634_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_7 _4014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__3152_ _6330_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3152_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5285_ _6922_/Q _6914_/Q _7031_/Q _7047_/Q _4066_/A _4063_/A vssd1 vssd1 vccd1 vccd1
+ _5285_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7024_ _7030_/CLK _7024_/D vssd1 vssd1 vccd1 vccd1 _7024_/Q sky130_fd_sc_hd__dfxtp_1
X_4236_ _4236_/A vssd1 vssd1 vccd1 vccd1 _6664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ _4167_/A _4167_/B _3708_/A vssd1 vssd1 vccd1 vccd1 _4662_/B sky130_fd_sc_hd__or3b_4
XFILLER_67_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4098_ _4098_/A vssd1 vssd1 vccd1 vccd1 _6725_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6808_ _6808_/CLK _6808_/D vssd1 vssd1 vccd1 vccd1 _6808_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2867_ _5821_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2867_/X sky130_fd_sc_hd__clkbuf_16
X_6739_ _6739_/CLK _6739_/D vssd1 vssd1 vccd1 vccd1 _6739_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_109_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5569__391 _5569__391/A vssd1 vssd1 vccd1 vccd1 _6681_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6108__149 _6108__149/A vssd1 vssd1 vccd1 vccd1 _6957_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6362__45 _6363__46/A vssd1 vssd1 vccd1 vccd1 _7065_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5070_ _5070_/A vssd1 vssd1 vccd1 vccd1 _6452_/D sky130_fd_sc_hd__clkbuf_1
X_4021_ _4020_/X _6755_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5972_ _5972_/A _5972_/B vssd1 vssd1 vccd1 vccd1 _5973_/A sky130_fd_sc_hd__and2_1
X_4923_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__buf_6
X_4854_ _4850_/X _4852_/X _4853_/X _4909_/A _3953_/A vssd1 vssd1 vccd1 vccd1 _4854_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3805_ _3702_/X _6829_/Q _3807_/S vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__mux2_1
X_4785_ _4878_/S vssd1 vssd1 vccd1 vccd1 _4900_/S sky130_fd_sc_hd__buf_4
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6524_ _6524_/CLK _6524_/D vssd1 vssd1 vccd1 vccd1 _6524_/Q sky130_fd_sc_hd__dfxtp_1
X_3736_ _3693_/X _6856_/Q _3738_/S vssd1 vssd1 vccd1 vccd1 _3737_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3667_ _3667_/A vssd1 vssd1 vccd1 vccd1 _6904_/D sky130_fd_sc_hd__clkbuf_1
X_6455_ _7096_/CLK _6455_/D vssd1 vssd1 vccd1 vccd1 _6455_/Q sky130_fd_sc_hd__dfxtp_1
X_6386_ _6389_/A _6386_/B vssd1 vssd1 vccd1 vccd1 _6387_/A sky130_fd_sc_hd__and2_1
X_5406_ _6019_/B vssd1 vssd1 vccd1 vccd1 _5406_/X sky130_fd_sc_hd__clkbuf_2
X_3598_ _3623_/A _4040_/A _4368_/A vssd1 vssd1 vccd1 vccd1 _3621_/S sky130_fd_sc_hd__nor3_4
XFILLER_102_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5337_ _5337_/A vssd1 vssd1 vccd1 vccd1 _5337_/X sky130_fd_sc_hd__buf_2
XFILLER_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5268_ _5330_/A vssd1 vssd1 vccd1 vccd1 _5268_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7007_ _7011_/CLK _7007_/D vssd1 vssd1 vccd1 vccd1 _7007_/Q sky130_fd_sc_hd__dfxtp_2
X_4219_ _6671_/Q _4161_/X _4221_/S vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5456__300 _5458__302/A vssd1 vssd1 vccd1 vccd1 _6590_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5792__485 _5796__489/A vssd1 vssd1 vccd1 vccd1 _6791_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5855__55 _5857__57/A vssd1 vssd1 vccd1 vccd1 _6841_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6032__88 _6032__88/A vssd1 vssd1 vccd1 vccd1 _6895_/CLK sky130_fd_sc_hd__inv_2
X_5550__376 _5550__376/A vssd1 vssd1 vccd1 vccd1 _6666_/CLK sky130_fd_sc_hd__inv_2
X_4570_ _6510_/Q _4032_/A _4570_/S vssd1 vssd1 vccd1 vccd1 _4571_/A sky130_fd_sc_hd__mux2_1
X_3521_ _3521_/A vssd1 vssd1 vccd1 vccd1 _6963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3021_ clkbuf_0__3021_/X vssd1 vssd1 vccd1 vccd1 _6150__7/A sky130_fd_sc_hd__clkbuf_4
X_6240_ _7005_/Q vssd1 vssd1 vccd1 vccd1 _6250_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3452_ _3452_/A vssd1 vssd1 vccd1 vccd1 _6990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6171_ _4978_/X _6163_/Y _6162_/Y _4974_/X _6170_/Y vssd1 vssd1 vccd1 vccd1 _6171_/X
+ sky130_fd_sc_hd__o221a_1
X_3383_ _7025_/Q vssd1 vssd1 vccd1 vccd1 _3782_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _6445_/Q _7099_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__mux2_1
X_4004_ _4004_/A vssd1 vssd1 vccd1 vccd1 _6761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__2736_ clkbuf_0__2736_/X vssd1 vssd1 vccd1 vccd1 _5502__337/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5713__442 _5713__442/A vssd1 vssd1 vccd1 vccd1 _6736_/CLK sky130_fd_sc_hd__inv_2
X_5955_ _7126_/A _3242_/X _6433_/A vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__a21o_4
X_4906_ _4906_/A vssd1 vssd1 vccd1 vccd1 _4906_/X sky130_fd_sc_hd__buf_4
XFILLER_80_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4837_ _4878_/S vssd1 vssd1 vccd1 vccd1 _4898_/A sky130_fd_sc_hd__buf_2
X_5451__296 _5454__299/A vssd1 vssd1 vccd1 vccd1 _6586_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4768_ _4909_/A vssd1 vssd1 vccd1 vccd1 _4933_/S sky130_fd_sc_hd__buf_2
X_5189__245 _5190__246/A vssd1 vssd1 vccd1 vccd1 _6527_/CLK sky130_fd_sc_hd__inv_2
X_6507_ _6507_/CLK _6507_/D vssd1 vssd1 vccd1 vccd1 _6507_/Q sky130_fd_sc_hd__dfxtp_1
X_3719_ _3696_/X _6863_/Q _3719_/S vssd1 vssd1 vccd1 vccd1 _3720_/A sky130_fd_sc_hd__mux2_1
X_4699_ _4845_/A vssd1 vssd1 vccd1 vccd1 _4914_/A sky130_fd_sc_hd__buf_4
XFILLER_107_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6438_ _6438_/CLK _6438_/D vssd1 vssd1 vccd1 vccd1 _6438_/Q sky130_fd_sc_hd__dfxtp_1
X_6057__107 _6059__109/A vssd1 vssd1 vccd1 vccd1 _6915_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5800__492 _5802__494/A vssd1 vssd1 vccd1 vccd1 _6798_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5133__200 _5137__204/A vssd1 vssd1 vccd1 vccd1 _6482_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5842__526 _5845__529/A vssd1 vssd1 vccd1 vccd1 _6832_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6148__5 _6150__7/A vssd1 vssd1 vccd1 vccd1 _6988_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2521_ clkbuf_0__2521_/X vssd1 vssd1 vccd1 vccd1 _5181__239/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5740_ _5740_/A vssd1 vssd1 vccd1 vccd1 _6750_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ _6180_/A _6994_/Q vssd1 vssd1 vccd1 vccd1 _6271_/B sky130_fd_sc_hd__nor2_1
X_4622_ _3865_/X _6487_/Q _4624_/S vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4553_ _4553_/A vssd1 vssd1 vccd1 vccd1 _6519_/D sky130_fd_sc_hd__clkbuf_1
X_4484_ _6746_/Q vssd1 vssd1 vccd1 vccd1 _4484_/X sky130_fd_sc_hd__buf_2
X_3504_ _3504_/A vssd1 vssd1 vccd1 vccd1 _6970_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6223_ _7001_/Q _6249_/C _6250_/C vssd1 vssd1 vccd1 vccd1 _6228_/B sky130_fd_sc_hd__and3_1
Xclkbuf_1_1_0__3004_ clkbuf_0__3004_/X vssd1 vssd1 vccd1 vccd1 _6065__114/A sky130_fd_sc_hd__clkbuf_4
X_3435_ _3392_/X _7031_/Q _3435_/S vssd1 vssd1 vccd1 vccd1 _3436_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3366_ _3366_/A vssd1 vssd1 vccd1 vccd1 _7054_/D sky130_fd_sc_hd__clkbuf_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _6775_/Q vssd1 vssd1 vccd1 vccd1 _4167_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _7126_/A _3242_/X _6433_/A vssd1 vssd1 vccd1 vccd1 _6013_/A sky130_fd_sc_hd__a21oi_4
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6085_/X sky130_fd_sc_hd__buf_1
X_5036_ _5206_/A vssd1 vssd1 vccd1 vccd1 _5036_/X sky130_fd_sc_hd__buf_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3151_ clkbuf_0__3151_/X vssd1 vssd1 vccd1 vccd1 _6328__18/A sky130_fd_sc_hd__clkbuf_4
X_6987_ _6987_/CLK _6987_/D vssd1 vssd1 vccd1 vccd1 _6987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5938_ _5937_/Y _5936_/X _5954_/B vssd1 vssd1 vccd1 vccd1 _5938_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput101 wbs_sel_i[0] vssd1 vssd1 vccd1 vccd1 _7157_/A sky130_fd_sc_hd__buf_4
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5469__310 _5470__311/A vssd1 vssd1 vccd1 vccd1 _6600_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5807__498 _5808__499/A vssd1 vssd1 vccd1 vccd1 _6804_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7095_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_3220_ _6737_/Q vssd1 vssd1 vccd1 vccd1 _4277_/C sky130_fd_sc_hd__clkinv_2
XFILLER_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6910_ _6910_/CLK _6910_/D vssd1 vssd1 vccd1 vccd1 _6910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6841_ _6841_/CLK _6841_/D vssd1 vssd1 vccd1 vccd1 _6841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ _4868_/S vssd1 vssd1 vccd1 vccd1 _4851_/S sky130_fd_sc_hd__clkbuf_2
X_6772_ _6772_/CLK _6772_/D vssd1 vssd1 vccd1 vccd1 _6772_/Q sky130_fd_sc_hd__dfxtp_1
X_5723_ _7017_/Q _5723_/B vssd1 vssd1 vccd1 vccd1 _5724_/A sky130_fd_sc_hd__and2_1
X_5654_ _7002_/Q _5917_/B _5917_/C vssd1 vssd1 vccd1 vccd1 _5657_/C sky130_fd_sc_hd__and3_1
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4605_ _4605_/A vssd1 vssd1 vccd1 vccd1 _6495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5585_ _5585_/A vssd1 vssd1 vccd1 vccd1 _6694_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4536_ _4499_/X _6526_/Q _4536_/S vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__mux2_1
X_4467_ _4467_/A vssd1 vssd1 vccd1 vccd1 _6554_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5563__386 _5564__387/A vssd1 vssd1 vccd1 vccd1 _6676_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6206_ _6206_/A vssd1 vssd1 vccd1 vccd1 _6997_/D sky130_fd_sc_hd__clkbuf_1
X_4398_ _3263_/X _6592_/Q _4402_/S vssd1 vssd1 vccd1 vccd1 _4399_/A sky130_fd_sc_hd__mux2_1
X_3418_ _4048_/A _4051_/A _3418_/C vssd1 vssd1 vccd1 vccd1 _4422_/B sky130_fd_sc_hd__or3_4
XFILLER_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3349_ _4029_/A vssd1 vssd1 vccd1 vccd1 _3349_/X sky130_fd_sc_hd__clkbuf_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5019_ _5019_/A vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5772__472 _5773__473/A vssd1 vssd1 vccd1 vccd1 _6776_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5370_ _6674_/Q _6666_/Q _6658_/Q _6650_/Q _5257_/X _5259_/X vssd1 vssd1 vccd1 vccd1
+ _5370_/X sky130_fd_sc_hd__mux4_2
X_4321_ _4321_/A vssd1 vssd1 vccd1 vccd1 _6627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7040_ _7040_/CLK _7040_/D vssd1 vssd1 vccd1 vccd1 _7040_/Q sky130_fd_sc_hd__dfxtp_1
X_4252_ _4252_/A vssd1 vssd1 vccd1 vccd1 _6657_/D sky130_fd_sc_hd__clkbuf_1
X_5146__210 _5147__211/A vssd1 vssd1 vccd1 vccd1 _6492_/CLK sky130_fd_sc_hd__inv_2
X_3203_ _4204_/A _4044_/A _6739_/Q vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__or3b_2
X_4183_ _4183_/A vssd1 vssd1 vccd1 vccd1 _6687_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6824_ _6824_/CLK _6824_/D vssd1 vssd1 vccd1 vccd1 _6824_/Q sky130_fd_sc_hd__dfxtp_1
X_6755_ _6755_/CLK _6755_/D vssd1 vssd1 vccd1 vccd1 _6755_/Q sky130_fd_sc_hd__dfxtp_1
X_3967_ _3983_/A _3983_/B _3966_/X _6779_/Q vssd1 vssd1 vccd1 vccd1 _3977_/B sky130_fd_sc_hd__o211a_1
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6686_ _6686_/CLK _6686_/D vssd1 vssd1 vccd1 vccd1 _6686_/Q sky130_fd_sc_hd__dfxtp_1
X_3898_ _4205_/A _3898_/B vssd1 vssd1 vccd1 vccd1 _3914_/S sky130_fd_sc_hd__nor2_2
X_5637_ _5906_/B _5906_/C _6217_/B vssd1 vssd1 vccd1 vccd1 _5637_/X sky130_fd_sc_hd__a21bo_1
X_4519_ _4519_/A vssd1 vssd1 vccd1 vccd1 _6534_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5499_ _5499_/A vssd1 vssd1 vccd1 vccd1 _5499_/X sky130_fd_sc_hd__buf_1
XFILLER_77_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4870_ _4719_/X _4867_/X _4869_/X vssd1 vssd1 vccd1 vccd1 _4870_/X sky130_fd_sc_hd__a21o_1
XFILLER_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5514__347 _5514__347/A vssd1 vssd1 vccd1 vccd1 _6637_/CLK sky130_fd_sc_hd__inv_2
X_3821_ _6822_/Q _3614_/X _3825_/S vssd1 vssd1 vccd1 vccd1 _3822_/A sky130_fd_sc_hd__mux2_1
X_6540_ _6540_/CLK _6540_/D vssd1 vssd1 vccd1 vccd1 _6540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3752_ _6849_/Q _3605_/X _3756_/S vssd1 vssd1 vccd1 vccd1 _3753_/A sky130_fd_sc_hd__mux2_1
X_3683_ _4572_/A _4590_/B vssd1 vssd1 vccd1 vccd1 _3706_/S sky130_fd_sc_hd__or2_2
X_6471_ _6471_/CLK _6471_/D vssd1 vssd1 vccd1 vccd1 _6471_/Q sky130_fd_sc_hd__dfxtp_1
X_5422_ _5289_/X _5421_/X _5292_/X vssd1 vssd1 vccd1 vccd1 _5422_/Y sky130_fd_sc_hd__o21ai_1
Xoutput202 _4887_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[4] sky130_fd_sc_hd__buf_2
X_5353_ _5355_/B _5353_/B vssd1 vssd1 vccd1 vccd1 _5353_/Y sky130_fd_sc_hd__nor2_1
X_4304_ _3776_/X _6634_/Q _4306_/S vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3151_ _6324_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3151_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5284_ _5351_/B _5284_/B vssd1 vssd1 vccd1 vccd1 _5284_/Y sky130_fd_sc_hd__nor2_1
XINSDIODE2_8 _4026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4235_ _3782_/X _6664_/Q _4239_/S vssd1 vssd1 vccd1 vccd1 _4236_/A sky130_fd_sc_hd__mux2_1
X_7023_ _7079_/CLK _7023_/D vssd1 vssd1 vccd1 vccd1 _7023_/Q sky130_fd_sc_hd__dfxtp_1
X_5595__408 _5596__409/A vssd1 vssd1 vccd1 vccd1 _6701_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4166_ _4166_/A vssd1 vssd1 vccd1 vccd1 _6697_/D sky130_fd_sc_hd__clkbuf_1
X_4097_ _4023_/X _6725_/Q _4097_/S vssd1 vssd1 vccd1 vccd1 _4098_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6807_ _6807_/CLK _6807_/D vssd1 vssd1 vccd1 vccd1 _6807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4999_ _5003_/A _4999_/B vssd1 vssd1 vccd1 vccd1 _5000_/A sky130_fd_sc_hd__and2_1
XFILLER_23_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2866_ _5815_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2866_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6738_ _6738_/CLK _6738_/D vssd1 vssd1 vccd1 vccd1 _6738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6669_ _6669_/CLK _6669_/D vssd1 vssd1 vccd1 vccd1 _6669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5882__78 _5882__78/A vssd1 vssd1 vccd1 vccd1 _6864_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044__97 _6046__99/A vssd1 vssd1 vccd1 vccd1 _6905_/CLK sky130_fd_sc_hd__inv_2
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6050__102 _6052__104/A vssd1 vssd1 vccd1 vccd1 _6910_/CLK sky130_fd_sc_hd__inv_2
X_4020_ _4020_/A vssd1 vssd1 vccd1 vccd1 _4020_/X sky130_fd_sc_hd__buf_4
XFILLER_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5971_ _6876_/Q _5966_/X _5969_/Y _5970_/X vssd1 vssd1 vccd1 vccd1 _5972_/B sky130_fd_sc_hd__a22o_1
XFILLER_18_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4922_ _4944_/A _4922_/B vssd1 vssd1 vccd1 vccd1 _4922_/X sky130_fd_sc_hd__or2_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4853_ _6762_/Q _6754_/Q _6717_/Q _6709_/Q _4957_/S _4845_/X vssd1 vssd1 vccd1 vccd1
+ _4853_/X sky130_fd_sc_hd__mux4_2
X_4784_ _4726_/X _4770_/X _4777_/X _4783_/X _3971_/X vssd1 vssd1 vccd1 vccd1 _4784_/X
+ sky130_fd_sc_hd__a311o_1
X_3804_ _3804_/A vssd1 vssd1 vccd1 vccd1 _6830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6523_ _6523_/CLK _6523_/D vssd1 vssd1 vccd1 vccd1 _6523_/Q sky130_fd_sc_hd__dfxtp_1
X_3735_ _3735_/A vssd1 vssd1 vccd1 vccd1 _6857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6454_ _7096_/CLK _6454_/D vssd1 vssd1 vccd1 vccd1 _6454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3666_ _3329_/X _6904_/Q _3672_/S vssd1 vssd1 vccd1 vccd1 _3667_/A sky130_fd_sc_hd__mux2_1
X_5405_ _5324_/X _5394_/X _5404_/Y vssd1 vssd1 vccd1 vccd1 _5405_/X sky130_fd_sc_hd__a21o_1
X_6385_ _7140_/A _6161_/A _6401_/S vssd1 vssd1 vccd1 vccd1 _6386_/B sky130_fd_sc_hd__mux2_1
X_3597_ _7030_/Q vssd1 vssd1 vccd1 vccd1 _3597_/X sky130_fd_sc_hd__buf_4
XFILLER_114_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5336_ _5335_/X _5364_/S vssd1 vssd1 vccd1 vccd1 _5336_/X sky130_fd_sc_hd__and2b_1
XFILLER_102_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5267_ _5337_/A vssd1 vssd1 vccd1 vccd1 _5330_/A sky130_fd_sc_hd__clkbuf_4
X_7006_ _7019_/CLK _7006_/D vssd1 vssd1 vccd1 vccd1 _7006_/Q sky130_fd_sc_hd__dfxtp_1
X_4218_ _4218_/A vssd1 vssd1 vccd1 vccd1 _6672_/D sky130_fd_sc_hd__clkbuf_1
X_4149_ _7028_/Q vssd1 vssd1 vccd1 vccd1 _4149_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_28_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6374__2 _6376__4/A vssd1 vssd1 vccd1 vccd1 _7076_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7008_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6114__154 _6114__154/A vssd1 vssd1 vccd1 vccd1 _6962_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6335__24 _6335__24/A vssd1 vssd1 vccd1 vccd1 _7044_/CLK sky130_fd_sc_hd__inv_2
X_3520_ _6963_/Q _3459_/X _3522_/S vssd1 vssd1 vccd1 vccd1 _3521_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3020_ clkbuf_0__3020_/X vssd1 vssd1 vccd1 vccd1 _6330_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3451_ _6990_/Q _3450_/X _3454_/S vssd1 vssd1 vccd1 vccd1 _3452_/A sky130_fd_sc_hd__mux2_1
X_6170_ _6170_/A _7008_/Q vssd1 vssd1 vccd1 vccd1 _6170_/Y sky130_fd_sc_hd__xnor2_1
X_3382_ _3382_/A vssd1 vssd1 vccd1 vccd1 _7050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5052_ _5061_/A vssd1 vssd1 vccd1 vccd1 _5116_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4003_ _3699_/X _6761_/Q _4007_/S vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5954_ _6873_/Q _5954_/B vssd1 vssd1 vccd1 vccd1 _5954_/Y sky130_fd_sc_hd__nand2_1
X_5885_ _6028_/A vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__buf_1
X_4905_ _4905_/A vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4836_ _4834_/X _4835_/X _4875_/S vssd1 vssd1 vccd1 vccd1 _4836_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6506_ _6506_/CLK _6506_/D vssd1 vssd1 vccd1 vccd1 _6506_/Q sky130_fd_sc_hd__dfxtp_1
X_4767_ _6769_/Q vssd1 vssd1 vccd1 vccd1 _4909_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3718_ _3718_/A vssd1 vssd1 vccd1 vccd1 _6864_/D sky130_fd_sc_hd__clkbuf_1
X_4698_ _4865_/A vssd1 vssd1 vccd1 vccd1 _4954_/S sky130_fd_sc_hd__clkbuf_4
X_6437_ _6437_/CLK _6437_/D vssd1 vssd1 vccd1 vccd1 _6437_/Q sky130_fd_sc_hd__dfxtp_1
X_3649_ _3333_/X _6911_/Q _3653_/S vssd1 vssd1 vccd1 vccd1 _3650_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5319_ _5315_/X _5318_/X _5433_/S vssd1 vssd1 vccd1 vccd1 _5320_/B sky130_fd_sc_hd__mux2_1
X_6299_ _7022_/Q _6284_/A _6298_/X _6290_/X vssd1 vssd1 vccd1 vccd1 _7021_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2520_ clkbuf_0__2520_/X vssd1 vssd1 vccd1 vccd1 _5200_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5670_ _6995_/Q vssd1 vssd1 vccd1 vccd1 _6180_/A sky130_fd_sc_hd__inv_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4621_ _4621_/A vssd1 vssd1 vccd1 vccd1 _6488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4552_ _4496_/X _6519_/Q _4554_/S vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__mux2_1
X_4483_ _4483_/A vssd1 vssd1 vccd1 vccd1 _6548_/D sky130_fd_sc_hd__clkbuf_1
X_3503_ _3353_/X _6970_/Q _3503_/S vssd1 vssd1 vccd1 vccd1 _3504_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6222_ _6222_/A vssd1 vssd1 vccd1 vccd1 _7000_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3003_ clkbuf_0__3003_/X vssd1 vssd1 vccd1 vccd1 _6055__105/A sky130_fd_sc_hd__clkbuf_4
X_3434_ _3434_/A vssd1 vssd1 vccd1 vccd1 _7032_/D sky130_fd_sc_hd__clkbuf_1
X_6153_ _6336_/A vssd1 vssd1 vccd1 vccd1 _6153_/X sky130_fd_sc_hd__buf_1
X_3365_ _3357_/X _7054_/Q _3381_/S vssd1 vssd1 vccd1 vccd1 _3366_/A sky130_fd_sc_hd__mux2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3296_ _3708_/A vssd1 vssd1 vccd1 vccd1 _3990_/C sky130_fd_sc_hd__clkbuf_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6084_/A vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__buf_1
X_5104_ _5248_/B vssd1 vssd1 vccd1 vccd1 _5929_/B sky130_fd_sc_hd__clkbuf_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6986_ _6986_/CLK _6986_/D vssd1 vssd1 vccd1 vccd1 _6986_/Q sky130_fd_sc_hd__dfxtp_1
X_5195__250 _5196__251/A vssd1 vssd1 vccd1 vccd1 _6532_/CLK sky130_fd_sc_hd__inv_2
X_5937_ _5945_/C vssd1 vssd1 vccd1 vccd1 _5937_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6063__112 _6064__113/A vssd1 vssd1 vccd1 vccd1 _6920_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4819_ _4815_/X _4817_/X _4818_/X _4716_/A _4711_/X vssd1 vssd1 vccd1 vccd1 _4819_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2865_ clkbuf_0__2865_/X vssd1 vssd1 vccd1 vccd1 _5813__503/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput102 wbs_sel_i[1] vssd1 vssd1 vccd1 vccd1 _7158_/A sky130_fd_sc_hd__buf_4
XFILLER_102_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6150__7 _6150__7/A vssd1 vssd1 vccd1 vccd1 _6990_/CLK sky130_fd_sc_hd__inv_2
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6840_ _6840_/CLK _6840_/D vssd1 vssd1 vccd1 vccd1 _6840_/Q sky130_fd_sc_hd__dfxtp_1
X_6771_ _6771_/CLK _6771_/D vssd1 vssd1 vccd1 vccd1 _6771_/Q sky130_fd_sc_hd__dfxtp_1
X_5722_ _5722_/A vssd1 vssd1 vccd1 vccd1 _6742_/D sky130_fd_sc_hd__clkbuf_1
X_3983_ _3983_/A _3983_/B vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__nor2_2
X_6127__164 _6127__164/A vssd1 vssd1 vccd1 vccd1 _6972_/CLK sky130_fd_sc_hd__inv_2
X_5653_ _5653_/A _5653_/B _5653_/C vssd1 vssd1 vccd1 vccd1 _5657_/B sky130_fd_sc_hd__or3_1
XFILLER_31_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4604_ _6495_/Q _4029_/A _4606_/S vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__mux2_1
X_5584_ _6427_/A _7157_/A _5586_/S vssd1 vssd1 vccd1 vccd1 _5585_/A sky130_fd_sc_hd__mux2_1
X_4535_ _4535_/A vssd1 vssd1 vccd1 vccd1 _6527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4466_ _4020_/X _6554_/Q _4468_/S vssd1 vssd1 vccd1 vccd1 _4467_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6205_ _6238_/A _6205_/B _6205_/C vssd1 vssd1 vccd1 vccd1 _6206_/A sky130_fd_sc_hd__and3_1
X_3417_ _3417_/A vssd1 vssd1 vccd1 vccd1 _7039_/D sky130_fd_sc_hd__clkbuf_1
X_4397_ _4397_/A vssd1 vssd1 vccd1 vccd1 _6593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3348_ _6742_/Q vssd1 vssd1 vccd1 vccd1 _4029_/A sky130_fd_sc_hd__buf_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3279_ _7069_/Q _3251_/X _3285_/S vssd1 vssd1 vccd1 vccd1 _3280_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5018_ _5018_/A _5018_/B vssd1 vssd1 vccd1 vccd1 _5019_/A sky130_fd_sc_hd__and2_2
XFILLER_26_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6969_ _6969_/CLK _6969_/D vssd1 vssd1 vccd1 vccd1 _6969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4320_ _6627_/Q _3880_/X _4324_/S vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4251_ _3779_/X _6657_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3202_ _6737_/Q vssd1 vssd1 vccd1 vccd1 _4044_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4182_ _4029_/X _6687_/Q _4184_/S vssd1 vssd1 vccd1 vccd1 _4183_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6823_ _6823_/CLK _6823_/D vssd1 vssd1 vccd1 vccd1 _6823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6754_ _6754_/CLK _6754_/D vssd1 vssd1 vccd1 vccd1 _6754_/Q sky130_fd_sc_hd__dfxtp_1
X_3966_ _4807_/S vssd1 vssd1 vccd1 vccd1 _3966_/X sky130_fd_sc_hd__buf_4
X_6685_ _6685_/CLK _6685_/D vssd1 vssd1 vccd1 vccd1 _6685_/Q sky130_fd_sc_hd__dfxtp_1
X_3897_ _3897_/A vssd1 vssd1 vccd1 vccd1 _6796_/D sky130_fd_sc_hd__clkbuf_1
X_5636_ _6998_/Q vssd1 vssd1 vccd1 vccd1 _6217_/B sky130_fd_sc_hd__clkbuf_2
X_5567_ _5573_/A vssd1 vssd1 vccd1 vccd1 _5567_/X sky130_fd_sc_hd__buf_1
X_4518_ _4499_/X _6534_/Q _4518_/S vssd1 vssd1 vccd1 vccd1 _4519_/A sky130_fd_sc_hd__mux2_1
X_5498_ _5560_/A vssd1 vssd1 vccd1 vccd1 _5498_/X sky130_fd_sc_hd__buf_1
X_4449_ _4449_/A vssd1 vssd1 vccd1 vccd1 _6562_/D sky130_fd_sc_hd__clkbuf_1
X_7099_ _7099_/A vssd1 vssd1 vccd1 vccd1 _7099_/X sky130_fd_sc_hd__clkbuf_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3820_ _3820_/A vssd1 vssd1 vccd1 vccd1 _6823_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3751_ _3751_/A vssd1 vssd1 vccd1 vccd1 _6850_/D sky130_fd_sc_hd__clkbuf_1
X_3682_ _3990_/C _3990_/B _3727_/B vssd1 vssd1 vccd1 vccd1 _4590_/B sky130_fd_sc_hd__nand3b_4
X_6470_ _6470_/CLK _6470_/D vssd1 vssd1 vccd1 vccd1 _6470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5421_ _6960_/Q _6944_/Q _7069_/Q _6936_/Q _5266_/X _5268_/X vssd1 vssd1 vccd1 vccd1
+ _5421_/X sky130_fd_sc_hd__mux4_2
Xoutput203 _4920_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[5] sky130_fd_sc_hd__buf_2
X_5352_ _6949_/Q _6681_/Q _6593_/Q _6815_/Q _4083_/X _4070_/A vssd1 vssd1 vccd1 vccd1
+ _5353_/B sky130_fd_sc_hd__mux4_1
X_4303_ _4303_/A vssd1 vssd1 vccd1 vccd1 _6635_/D sky130_fd_sc_hd__clkbuf_1
X_7022_ _7022_/CLK _7022_/D vssd1 vssd1 vccd1 vccd1 _7022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5283_ _6946_/Q _6678_/Q _6590_/Q _6812_/Q _5281_/X _5282_/X vssd1 vssd1 vccd1 vccd1
+ _5284_/B sky130_fd_sc_hd__mux4_1
X_4234_ _4234_/A vssd1 vssd1 vccd1 vccd1 _6665_/D sky130_fd_sc_hd__clkbuf_1
XINSDIODE2_9 _4152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4165_ _6697_/Q _4164_/X _4165_/S vssd1 vssd1 vccd1 vccd1 _4166_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4096_ _4096_/A vssd1 vssd1 vccd1 vccd1 _6726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2865_ _5809_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2865_/X sky130_fd_sc_hd__clkbuf_16
X_6806_ _6806_/CLK _6806_/D vssd1 vssd1 vccd1 vccd1 _6806_/Q sky130_fd_sc_hd__dfxtp_1
X_4998_ _4998_/A vssd1 vssd1 vccd1 vccd1 _4998_/X sky130_fd_sc_hd__clkbuf_1
X_3949_ _3949_/A _5774_/C _3949_/C vssd1 vssd1 vccd1 vccd1 _3950_/A sky130_fd_sc_hd__and3_1
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6737_ _6737_/CLK _6737_/D vssd1 vssd1 vccd1 vccd1 _6737_/Q sky130_fd_sc_hd__dfxtp_2
X_6668_ _6668_/CLK _6668_/D vssd1 vssd1 vccd1 vccd1 _6668_/Q sky130_fd_sc_hd__dfxtp_1
X_5619_ _5619_/A vssd1 vssd1 vccd1 vccd1 _5913_/A sky130_fd_sc_hd__buf_2
X_6599_ _6599_/CLK _6599_/D vssd1 vssd1 vccd1 vccd1 _6599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5867__65 _5870__68/A vssd1 vssd1 vccd1 vccd1 _6851_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5576__397 _5578__399/A vssd1 vssd1 vccd1 vccd1 _6687_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6347__33 _6347__33/A vssd1 vssd1 vccd1 vccd1 _7053_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5520__352 _5522__354/A vssd1 vssd1 vccd1 vccd1 _6642_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__2751_ clkbuf_0__2751_/X vssd1 vssd1 vccd1 vccd1 _5583__403/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5970_ _5970_/A vssd1 vssd1 vccd1 vccd1 _5970_/X sky130_fd_sc_hd__clkbuf_2
X_4921_ _6508_/Q _6442_/Q _6540_/Q _6692_/Q _4778_/X _4914_/X vssd1 vssd1 vccd1 vccd1
+ _4922_/B sky130_fd_sc_hd__mux4_2
X_4852_ _4808_/X _4851_/X _4718_/A vssd1 vssd1 vccd1 vccd1 _4852_/X sky130_fd_sc_hd__a21o_1
X_3803_ _3699_/X _6830_/Q _3807_/S vssd1 vssd1 vccd1 vccd1 _3804_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4783_ _4954_/S _4779_/X _4781_/X _4782_/X vssd1 vssd1 vccd1 vccd1 _4783_/X sky130_fd_sc_hd__o211a_1
X_6522_ _6522_/CLK _6522_/D vssd1 vssd1 vccd1 vccd1 _6522_/Q sky130_fd_sc_hd__dfxtp_1
X_3734_ _3690_/X _6857_/Q _3738_/S vssd1 vssd1 vccd1 vccd1 _3735_/A sky130_fd_sc_hd__mux2_1
X_3665_ _3665_/A vssd1 vssd1 vccd1 vccd1 _6905_/D sky130_fd_sc_hd__clkbuf_1
X_6453_ _6750_/CLK _6453_/D vssd1 vssd1 vccd1 vccd1 _6453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5404_ _5324_/A _5403_/X _5321_/A vssd1 vssd1 vccd1 vccd1 _5404_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6384_ _6407_/S vssd1 vssd1 vccd1 vccd1 _6401_/S sky130_fd_sc_hd__clkbuf_2
X_3596_ _3596_/A vssd1 vssd1 vccd1 vccd1 _6930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5335_ _6790_/Q _6980_/Q _6988_/Q _6964_/Q _5264_/A _5276_/X vssd1 vssd1 vccd1 vccd1
+ _5335_/X sky130_fd_sc_hd__mux4_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5266_ _5329_/A vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__buf_4
X_7005_ _7019_/CLK _7005_/D vssd1 vssd1 vccd1 vccd1 _7005_/Q sky130_fd_sc_hd__dfxtp_2
X_4217_ _6672_/Q _4158_/X _4221_/S vssd1 vssd1 vccd1 vccd1 _4218_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ _4148_/A vssd1 vssd1 vccd1 vccd1 _6703_/D sky130_fd_sc_hd__clkbuf_1
X_4079_ _4071_/B _4081_/A _4078_/Y vssd1 vssd1 vccd1 vccd1 _6732_/D sky130_fd_sc_hd__o21a_1
X_5159__221 _5160__222/A vssd1 vssd1 vccd1 vccd1 _6503_/CLK sky130_fd_sc_hd__inv_2
XFILLER_71_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5463__306 _5464__307/A vssd1 vssd1 vccd1 vccd1 _6596_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5812__502 _5814__504/A vssd1 vssd1 vccd1 vccd1 _6808_/CLK sky130_fd_sc_hd__inv_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6121__159 _6121__159/A vssd1 vssd1 vccd1 vccd1 _6967_/CLK sky130_fd_sc_hd__inv_2
X_3450_ _3776_/A vssd1 vssd1 vccd1 vccd1 _3450_/X sky130_fd_sc_hd__clkbuf_4
X_3381_ _3380_/X _7050_/Q _3381_/S vssd1 vssd1 vccd1 vccd1 _3382_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5120_ _5138_/A vssd1 vssd1 vccd1 vccd1 _5120_/X sky130_fd_sc_hd__buf_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5051_ _6391_/A _5113_/B _5113_/C vssd1 vssd1 vccd1 vccd1 _5061_/A sky130_fd_sc_hd__and3_1
XFILLER_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4002_ _4002_/A vssd1 vssd1 vccd1 vccd1 _6762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2734_ clkbuf_0__2734_/X vssd1 vssd1 vccd1 vccd1 _5497__334/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5953_ _5961_/C _5953_/B _5952_/X vssd1 vssd1 vccd1 vccd1 _5953_/X sky130_fd_sc_hd__or3b_1
X_4904_ _4904_/A _4904_/B _4904_/C vssd1 vssd1 vccd1 vccd1 _4904_/X sky130_fd_sc_hd__or3_1
X_5884_ _6115_/A vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__buf_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4835_ _6481_/Q _6553_/Q _7042_/Q _6973_/Q _4923_/A _3958_/A vssd1 vssd1 vccd1 vccd1
+ _4835_/X sky130_fd_sc_hd__mux4_1
XFILLER_61_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4766_ _4795_/B _4766_/B _4766_/C vssd1 vssd1 vccd1 vccd1 _4766_/Y sky130_fd_sc_hd__nor3_1
XFILLER_119_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6505_ _6505_/CLK _6505_/D vssd1 vssd1 vccd1 vccd1 _6505_/Q sky130_fd_sc_hd__dfxtp_1
X_3717_ _3693_/X _6864_/Q _3719_/S vssd1 vssd1 vccd1 vccd1 _3718_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4697_ _4732_/A vssd1 vssd1 vccd1 vccd1 _4865_/A sky130_fd_sc_hd__buf_2
X_3648_ _3648_/A vssd1 vssd1 vccd1 vccd1 _6912_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2881_ clkbuf_0__2881_/X vssd1 vssd1 vccd1 vccd1 _6027__84/A sky130_fd_sc_hd__clkbuf_4
X_6436_ _6436_/CLK _6436_/D vssd1 vssd1 vccd1 vccd1 _6436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6367_ _6367_/A vssd1 vssd1 vccd1 vccd1 _6367_/X sky130_fd_sc_hd__buf_1
X_3579_ _3579_/A _3827_/A vssd1 vssd1 vccd1 vccd1 _3595_/S sky130_fd_sc_hd__nor2_2
X_5527__358 _5527__358/A vssd1 vssd1 vccd1 vccd1 _6648_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5318_ _5316_/X _5317_/X _5364_/S vssd1 vssd1 vccd1 vccd1 _5318_/X sky130_fd_sc_hd__mux2_1
X_6298_ _7021_/Q _6300_/B vssd1 vssd1 vccd1 vccd1 _6298_/X sky130_fd_sc_hd__or2_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5249_ _5321_/A vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5140__206 _5140__206/A vssd1 vssd1 vccd1 vccd1 _6488_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _3862_/X _6488_/Q _4624_/S vssd1 vssd1 vccd1 vccd1 _4621_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4551_ _4551_/A vssd1 vssd1 vccd1 vccd1 _6520_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4482_ _4481_/X _6548_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__mux2_1
X_3502_ _3502_/A vssd1 vssd1 vccd1 vccd1 _6971_/D sky130_fd_sc_hd__clkbuf_1
X_6221_ _6224_/B _6267_/A _6221_/C vssd1 vssd1 vccd1 vccd1 _6222_/A sky130_fd_sc_hd__and3b_1
Xclkbuf_1_1_0__3002_ clkbuf_0__3002_/X vssd1 vssd1 vccd1 vccd1 _6072_/A sky130_fd_sc_hd__clkbuf_4
X_3433_ _3388_/X _7032_/Q _3435_/S vssd1 vssd1 vccd1 vccd1 _3434_/A sky130_fd_sc_hd__mux2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3364_ _3393_/S vssd1 vssd1 vccd1 vccd1 _3381_/S sky130_fd_sc_hd__clkbuf_2
X_5819__508 _5820__509/A vssd1 vssd1 vccd1 vccd1 _6814_/CLK sky130_fd_sc_hd__inv_2
X_5103_ _6868_/Q vssd1 vssd1 vccd1 vccd1 _5248_/B sky130_fd_sc_hd__inv_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3295_ _6776_/Q vssd1 vssd1 vccd1 vccd1 _3708_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6985_ _6985_/CLK _6985_/D vssd1 vssd1 vccd1 vccd1 _6985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5936_ _5970_/A vssd1 vssd1 vccd1 vccd1 _5936_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5533__362 _5535__364/A vssd1 vssd1 vccd1 vccd1 _6652_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4818_ _6544_/Q _6724_/Q _6862_/Q _6528_/Q _3958_/A _4807_/S vssd1 vssd1 vccd1 vccd1
+ _4818_/X sky130_fd_sc_hd__mux4_1
X_4749_ _5736_/B _4766_/B vssd1 vssd1 vccd1 vccd1 _4762_/C sky130_fd_sc_hd__and2_1
XFILLER_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6419_ _6425_/A _6419_/B vssd1 vssd1 vccd1 vccd1 _6420_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_0_0__2864_ clkbuf_0__2864_/X vssd1 vssd1 vccd1 vccd1 _5808__499/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput103 wbs_sel_i[2] vssd1 vssd1 vccd1 vccd1 _7159_/A sky130_fd_sc_hd__buf_4
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5204__258 _5205__259/A vssd1 vssd1 vccd1 vccd1 _6540_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5476__316 _5479__319/A vssd1 vssd1 vccd1 vccd1 _6606_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6770_ _6770_/CLK _6770_/D vssd1 vssd1 vccd1 vccd1 _6770_/Q sky130_fd_sc_hd__dfxtp_2
X_3982_ _6779_/Q vssd1 vssd1 vccd1 vccd1 _3982_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5721_ _7016_/Q _5723_/B vssd1 vssd1 vccd1 vccd1 _5722_/A sky130_fd_sc_hd__and2_1
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5652_ _5918_/A _5918_/B _5652_/C vssd1 vssd1 vccd1 vccd1 _5653_/C sky130_fd_sc_hd__and3b_1
XFILLER_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4603_ _4603_/A vssd1 vssd1 vccd1 vccd1 _6496_/D sky130_fd_sc_hd__clkbuf_1
X_5825__512 _5825__512/A vssd1 vssd1 vccd1 vccd1 _6818_/CLK sky130_fd_sc_hd__inv_2
X_4534_ _4496_/X _6527_/Q _4536_/S vssd1 vssd1 vccd1 vccd1 _4535_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4465_ _4465_/A vssd1 vssd1 vccd1 vccd1 _6555_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6204_ _6216_/B _6207_/C vssd1 vssd1 vccd1 vccd1 _6205_/C sky130_fd_sc_hd__or2_1
X_3416_ _3353_/X _7039_/Q _3416_/S vssd1 vssd1 vccd1 vccd1 _3417_/A sky130_fd_sc_hd__mux2_1
X_4396_ _3260_/X _6593_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4397_/A sky130_fd_sc_hd__mux2_1
X_3347_ _3347_/A vssd1 vssd1 vccd1 vccd1 _7057_/D sky130_fd_sc_hd__clkbuf_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6066_ _6078_/A vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__buf_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _3278_/A vssd1 vssd1 vccd1 vccd1 _7070_/D sky130_fd_sc_hd__clkbuf_1
X_5017_ _5017_/A vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6968_ _6968_/CLK _6968_/D vssd1 vssd1 vccd1 vccd1 _6968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6899_ _6899_/CLK _6899_/D vssd1 vssd1 vccd1 vccd1 _6899_/Q sky130_fd_sc_hd__dfxtp_1
X_5919_ _6874_/Q _5919_/B vssd1 vssd1 vccd1 vccd1 _5919_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5210__262 _5210__262/A vssd1 vssd1 vccd1 vccd1 _6544_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4250_ _4250_/A vssd1 vssd1 vccd1 vccd1 _6658_/D sky130_fd_sc_hd__clkbuf_1
X_4181_ _4181_/A vssd1 vssd1 vccd1 vccd1 _6688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3201_ _6738_/Q vssd1 vssd1 vccd1 vccd1 _4204_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6822_ _6822_/CLK _6822_/D vssd1 vssd1 vccd1 vccd1 _6822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2881_ _5885_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2881_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6753_ _6753_/CLK _6753_/D vssd1 vssd1 vccd1 vccd1 _6753_/Q sky130_fd_sc_hd__dfxtp_1
X_3965_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4807_/S sky130_fd_sc_hd__buf_4
X_5749__454 _5749__454/A vssd1 vssd1 vccd1 vccd1 _6758_/CLK sky130_fd_sc_hd__inv_2
X_5153__216 _5156__219/A vssd1 vssd1 vccd1 vccd1 _6498_/CLK sky130_fd_sc_hd__inv_2
X_3896_ _6796_/Q _3895_/X _3896_/S vssd1 vssd1 vccd1 vccd1 _3897_/A sky130_fd_sc_hd__mux2_1
X_5704_ _5716_/A vssd1 vssd1 vccd1 vccd1 _5704_/X sky130_fd_sc_hd__buf_1
X_6684_ _6684_/CLK _6684_/D vssd1 vssd1 vccd1 vccd1 _6684_/Q sky130_fd_sc_hd__dfxtp_1
X_5635_ _4760_/X _5910_/A _6173_/A vssd1 vssd1 vccd1 vccd1 _5906_/C sky130_fd_sc_hd__o21ai_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4517_ _4517_/A vssd1 vssd1 vccd1 vccd1 _6535_/D sky130_fd_sc_hd__clkbuf_1
X_4448_ _4020_/X _6562_/Q _4450_/S vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4379_ _4379_/A vssd1 vssd1 vccd1 vccd1 _6601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7098_ _7098_/A vssd1 vssd1 vccd1 vccd1 _7098_/X sky130_fd_sc_hd__buf_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6076__123 _6077__124/A vssd1 vssd1 vccd1 vccd1 _6931_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3750_ _6850_/Q _3602_/X _3756_/S vssd1 vssd1 vccd1 vccd1 _3751_/A sky130_fd_sc_hd__mux2_1
X_5217__268 _5218__269/A vssd1 vssd1 vccd1 vccd1 _6550_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3681_ _4644_/B vssd1 vssd1 vccd1 vccd1 _4572_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5420_ _5419_/X _5439_/B vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__and2b_1
XFILLER_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput204 _4942_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[6] sky130_fd_sc_hd__buf_2
X_5351_ _5350_/X _5351_/B vssd1 vssd1 vccd1 vccd1 _5351_/X sky130_fd_sc_hd__and2b_1
X_4302_ _3773_/X _6635_/Q _4306_/S vssd1 vssd1 vccd1 vccd1 _4303_/A sky130_fd_sc_hd__mux2_1
X_5282_ _5338_/A vssd1 vssd1 vccd1 vccd1 _5282_/X sky130_fd_sc_hd__clkbuf_4
X_7021_ _7022_/CLK _7021_/D vssd1 vssd1 vccd1 vccd1 _7021_/Q sky130_fd_sc_hd__dfxtp_1
X_4233_ _3779_/X _6665_/Q _4233_/S vssd1 vssd1 vccd1 vccd1 _4234_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4164_ _7023_/Q vssd1 vssd1 vccd1 vccd1 _4164_/X sky130_fd_sc_hd__buf_4
X_4095_ _4020_/X _6726_/Q _4097_/S vssd1 vssd1 vccd1 vccd1 _4096_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6805_ _6805_/CLK _6805_/D vssd1 vssd1 vccd1 vccd1 _6805_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2864_ _5803_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2864_/X sky130_fd_sc_hd__clkbuf_16
X_4997_ _5003_/A _4997_/B vssd1 vssd1 vccd1 vccd1 _4998_/A sky130_fd_sc_hd__and2_1
XFILLER_23_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6736_ _6736_/CLK _6736_/D vssd1 vssd1 vccd1 vccd1 _6736_/Q sky130_fd_sc_hd__dfxtp_1
X_3948_ _3948_/A _3948_/B vssd1 vssd1 vccd1 vccd1 _3949_/C sky130_fd_sc_hd__or2_1
X_5118__188 _5119__189/A vssd1 vssd1 vccd1 vccd1 _6470_/CLK sky130_fd_sc_hd__inv_2
X_3879_ _3879_/A vssd1 vssd1 vccd1 vccd1 _6802_/D sky130_fd_sc_hd__clkbuf_1
X_6667_ _6667_/CLK _6667_/D vssd1 vssd1 vccd1 vccd1 _6667_/Q sky130_fd_sc_hd__dfxtp_1
X_5618_ _5663_/A vssd1 vssd1 vccd1 vccd1 _5890_/A sky130_fd_sc_hd__inv_2
X_6598_ _6598_/CLK _6598_/D vssd1 vssd1 vccd1 vccd1 _6598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6029__85 _6032__88/A vssd1 vssd1 vccd1 vccd1 _6892_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2750_ clkbuf_0__2750_/X vssd1 vssd1 vccd1 vccd1 _5578__399/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4920_ _4888_/X input30/X _4890_/X _4919_/X vssd1 vssd1 vccd1 vccd1 _4920_/X sky130_fd_sc_hd__a22o_2
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4851_ _6473_/Q _7058_/Q _4851_/S vssd1 vssd1 vccd1 vccd1 _4851_/X sky130_fd_sc_hd__mux2_1
X_3802_ _3802_/A vssd1 vssd1 vccd1 vccd1 _6831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4782_ _6770_/Q vssd1 vssd1 vccd1 vccd1 _4782_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6521_ _6521_/CLK _6521_/D vssd1 vssd1 vccd1 vccd1 _6521_/Q sky130_fd_sc_hd__dfxtp_1
X_3733_ _3733_/A vssd1 vssd1 vccd1 vccd1 _6858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3664_ _3294_/X _6905_/Q _3672_/S vssd1 vssd1 vccd1 vccd1 _3665_/A sky130_fd_sc_hd__mux2_1
X_6452_ _6750_/CLK _6452_/D vssd1 vssd1 vccd1 vccd1 _6452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5403_ _5334_/X _5396_/X _5398_/Y _5400_/X _5402_/Y vssd1 vssd1 vccd1 vccd1 _5403_/X
+ sky130_fd_sc_hd__o32a_2
X_6383_ _6695_/Q _6427_/C vssd1 vssd1 vccd1 vccd1 _6407_/S sky130_fd_sc_hd__nand2_2
X_3595_ _6930_/Q _3462_/X _3595_/S vssd1 vssd1 vccd1 vccd1 _3596_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5334_ _5334_/A vssd1 vssd1 vccd1 vccd1 _5334_/X sky130_fd_sc_hd__clkbuf_2
X_5265_ _6638_/Q _6630_/Q _6614_/Q _6606_/Q _5263_/X _5264_/X vssd1 vssd1 vccd1 vccd1
+ _5265_/X sky130_fd_sc_hd__mux4_1
X_7004_ _7011_/CLK _7004_/D vssd1 vssd1 vccd1 vccd1 _7004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4216_ _4216_/A vssd1 vssd1 vccd1 vccd1 _6673_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4147_ _6703_/Q _4146_/X _4156_/S vssd1 vssd1 vccd1 vccd1 _4148_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4078_ _4071_/B _4081_/A _6303_/B vssd1 vssd1 vccd1 vccd1 _4078_/Y sky130_fd_sc_hd__a21boi_1
Xclkbuf_1_1_0__2879_ clkbuf_0__2879_/X vssd1 vssd1 vccd1 vccd1 _5882__78/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6719_ _6719_/CLK _6719_/D vssd1 vssd1 vccd1 vccd1 _6719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2529_ clkbuf_0__2529_/X vssd1 vssd1 vccd1 vccd1 _5224__274/A sky130_fd_sc_hd__clkbuf_4
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3380_ _3779_/A vssd1 vssd1 vccd1 vccd1 _3380_/X sky130_fd_sc_hd__buf_2
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5050_ _6435_/Q _5050_/B _5050_/C vssd1 vssd1 vccd1 vccd1 _5113_/C sky130_fd_sc_hd__and3_1
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4001_ _3696_/X _6762_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _4002_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6089__133 _6090__134/A vssd1 vssd1 vccd1 vccd1 _6941_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5952_ _6873_/Q _5952_/B vssd1 vssd1 vccd1 vccd1 _5952_/X sky130_fd_sc_hd__or2_1
Xclkbuf_1_1_0__2733_ clkbuf_0__2733_/X vssd1 vssd1 vccd1 vccd1 _5488__326/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4903_ _4899_/X _4901_/X _4902_/X _4933_/S _4782_/X vssd1 vssd1 vccd1 vccd1 _4904_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4834_ _6901_/Q _6561_/Q _6909_/Q _6489_/Q _4845_/A _4900_/S vssd1 vssd1 vccd1 vccd1
+ _4834_/X sky130_fd_sc_hd__mux4_1
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4765_ _4765_/A vssd1 vssd1 vccd1 vccd1 _4765_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6504_ _6504_/CLK _6504_/D vssd1 vssd1 vccd1 vccd1 _6504_/Q sky130_fd_sc_hd__dfxtp_1
X_3716_ _3716_/A vssd1 vssd1 vccd1 vccd1 _6865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4696_ _6769_/Q vssd1 vssd1 vccd1 vccd1 _4732_/A sky130_fd_sc_hd__inv_2
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _3329_/X _6912_/Q _3653_/S vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__2880_ clkbuf_0__2880_/X vssd1 vssd1 vccd1 vccd1 _6047_/A sky130_fd_sc_hd__clkbuf_4
X_6435_ _7096_/CLK _6435_/D vssd1 vssd1 vccd1 vccd1 _6435_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3578_ _3578_/A vssd1 vssd1 vccd1 vccd1 _6938_/D sky130_fd_sc_hd__clkbuf_1
X_6341__29 _6341__29/A vssd1 vssd1 vccd1 vccd1 _7049_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5317_ _6599_/Q _6583_/Q _6837_/Q _6821_/Q _5338_/A _5281_/X vssd1 vssd1 vccd1 vccd1
+ _5317_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6297_ _7021_/Q _6284_/A _6296_/X _6290_/X vssd1 vssd1 vccd1 vccd1 _7020_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5248_ _5929_/A _5248_/B _5739_/C vssd1 vssd1 vccd1 vccd1 _5321_/A sky130_fd_sc_hd__and3_1
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5688__422 _5688__422/A vssd1 vssd1 vccd1 vccd1 _6716_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4550_ _4493_/X _6520_/Q _4554_/S vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__mux2_1
X_4481_ _6747_/Q vssd1 vssd1 vccd1 vccd1 _4481_/X sky130_fd_sc_hd__buf_2
X_5743__449 _5743__449/A vssd1 vssd1 vccd1 vccd1 _6753_/CLK sky130_fd_sc_hd__inv_2
X_3501_ _3349_/X _6971_/Q _3503_/S vssd1 vssd1 vccd1 vccd1 _3502_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3001_ clkbuf_0__3001_/X vssd1 vssd1 vccd1 vccd1 _6052__104/A sky130_fd_sc_hd__clkbuf_4
X_6220_ _6216_/A _6213_/B _7000_/Q vssd1 vssd1 vccd1 vccd1 _6221_/C sky130_fd_sc_hd__a21o_1
X_3432_ _3432_/A vssd1 vssd1 vccd1 vccd1 _7033_/D sky130_fd_sc_hd__clkbuf_1
X_3363_ _3623_/A _4040_/A _4350_/A vssd1 vssd1 vccd1 vccd1 _3393_/S sky130_fd_sc_hd__or3_4
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _6869_/Q vssd1 vssd1 vccd1 vccd1 _5924_/D sky130_fd_sc_hd__clkbuf_2
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _4009_/A vssd1 vssd1 vccd1 vccd1 _3294_/X sky130_fd_sc_hd__buf_2
XFILLER_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6984_ _6984_/CLK _6984_/D vssd1 vssd1 vccd1 vccd1 _6984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5935_ _6013_/B _6017_/A vssd1 vssd1 vccd1 vccd1 _5970_/A sky130_fd_sc_hd__and2_1
X_5866_ _5866_/A vssd1 vssd1 vccd1 vccd1 _5866_/X sky130_fd_sc_hd__buf_1
XFILLER_34_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4817_ _4808_/X _4816_/X _4718_/A vssd1 vssd1 vccd1 vccd1 _4817_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5797_ _5809_/A vssd1 vssd1 vccd1 vccd1 _5797_/X sky130_fd_sc_hd__buf_1
XFILLER_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4748_ _4798_/A _4748_/B _4754_/B vssd1 vssd1 vccd1 vccd1 _4856_/B sky130_fd_sc_hd__or3_1
X_4679_ _4679_/A vssd1 vssd1 vccd1 vccd1 _6436_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2863_ clkbuf_0__2863_/X vssd1 vssd1 vccd1 vccd1 _5799__491/A sky130_fd_sc_hd__clkbuf_4
X_6418_ _7130_/A _5918_/A _6424_/S vssd1 vssd1 vccd1 vccd1 _6419_/B sky130_fd_sc_hd__mux2_1
X_6349_ _6355_/A vssd1 vssd1 vccd1 vccd1 _6349_/X sky130_fd_sc_hd__buf_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput104 wbs_sel_i[3] vssd1 vssd1 vccd1 vccd1 _7160_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6070__118 _6071__119/A vssd1 vssd1 vccd1 vccd1 _6926_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3981_ _3981_/A _3981_/B vssd1 vssd1 vccd1 vccd1 _6768_/D sky130_fd_sc_hd__nor2_1
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5720_ _5720_/A vssd1 vssd1 vccd1 vccd1 _6741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _5648_/X _5649_/X _6174_/A vssd1 vssd1 vccd1 vccd1 _5653_/B sky130_fd_sc_hd__mux2_1
X_4602_ _6496_/Q _4026_/A _4606_/S vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4533_ _4533_/A vssd1 vssd1 vccd1 vccd1 _6528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4464_ _4017_/X _6555_/Q _4468_/S vssd1 vssd1 vccd1 vccd1 _4465_/A sky130_fd_sc_hd__mux2_1
X_6203_ _6216_/B _6207_/C vssd1 vssd1 vccd1 vccd1 _6205_/B sky130_fd_sc_hd__nand2_1
X_3415_ _3415_/A vssd1 vssd1 vccd1 vccd1 _7040_/D sky130_fd_sc_hd__clkbuf_1
X_4395_ _4395_/A vssd1 vssd1 vccd1 vccd1 _6594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3346_ _3345_/X _7057_/Q _3354_/S vssd1 vssd1 vccd1 vccd1 _3347_/A sky130_fd_sc_hd__mux2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _6140_/A vssd1 vssd1 vccd1 vccd1 _6134_/X sky130_fd_sc_hd__buf_1
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5016_ _5018_/A _5016_/B vssd1 vssd1 vccd1 vccd1 _5017_/A sky130_fd_sc_hd__and2_2
X_3277_ _7070_/Q _3200_/X _3285_/S vssd1 vssd1 vccd1 vccd1 _3278_/A sky130_fd_sc_hd__mux2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _6967_/CLK _6967_/D vssd1 vssd1 vccd1 vccd1 _6967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5918_ _5918_/A _5918_/B vssd1 vssd1 vccd1 vccd1 _5919_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6898_ _6898_/CLK _6898_/D vssd1 vssd1 vccd1 vccd1 _6898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5581__401 _5590__404/A vssd1 vssd1 vccd1 vccd1 _6691_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2529_ _5219_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2529_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5482__321 _5483__322/A vssd1 vssd1 vccd1 vccd1 _6611_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4180_ _4026_/X _6688_/Q _4184_/S vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3200_ _7030_/Q vssd1 vssd1 vccd1 vccd1 _3200_/X sky130_fd_sc_hd__buf_2
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6821_ _6821_/CLK _6821_/D vssd1 vssd1 vccd1 vccd1 _6821_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2880_ _5884_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2880_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6752_ _6752_/CLK _6752_/D vssd1 vssd1 vccd1 vccd1 _6752_/Q sky130_fd_sc_hd__dfxtp_1
X_3964_ _4868_/S vssd1 vssd1 vccd1 vccd1 _4923_/A sky130_fd_sc_hd__clkbuf_2
X_3895_ _6741_/Q vssd1 vssd1 vccd1 vccd1 _3895_/X sky130_fd_sc_hd__clkbuf_4
X_5703_ _5756_/A vssd1 vssd1 vccd1 vccd1 _5703_/X sky130_fd_sc_hd__buf_1
XFILLER_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6683_ _6683_/CLK _6683_/D vssd1 vssd1 vccd1 vccd1 _6683_/Q sky130_fd_sc_hd__dfxtp_1
X_5634_ _6216_/A _5908_/B vssd1 vssd1 vccd1 vccd1 _5642_/C sky130_fd_sc_hd__nor2_1
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4516_ _4496_/X _6535_/Q _4518_/S vssd1 vssd1 vccd1 vccd1 _4517_/A sky130_fd_sc_hd__mux2_1
X_4447_ _4447_/A vssd1 vssd1 vccd1 vccd1 _6563_/D sky130_fd_sc_hd__clkbuf_1
X_5879__75 _5882__78/A vssd1 vssd1 vccd1 vccd1 _6861_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4378_ _6601_/Q _3779_/A _4378_/S vssd1 vssd1 vccd1 vccd1 _4379_/A sky130_fd_sc_hd__mux2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _4014_/A vssd1 vssd1 vccd1 vccd1 _3329_/X sky130_fd_sc_hd__buf_2
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7097_ _7097_/A vssd1 vssd1 vccd1 vccd1 _7097_/X sky130_fd_sc_hd__buf_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6888_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6359__43 _6360__44/A vssd1 vssd1 vccd1 vccd1 _7063_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5546__373 _5547__374/A vssd1 vssd1 vccd1 vccd1 _6663_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3680_ _4009_/A vssd1 vssd1 vccd1 vccd1 _3680_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput205 _4964_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[7] sky130_fd_sc_hd__buf_2
X_5350_ _6791_/Q _6981_/Q _6989_/Q _6965_/Q _5290_/X _4069_/A vssd1 vssd1 vccd1 vccd1
+ _5350_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4301_ _4301_/A vssd1 vssd1 vccd1 vccd1 _6636_/D sky130_fd_sc_hd__clkbuf_1
X_5281_ _5281_/A vssd1 vssd1 vccd1 vccd1 _5281_/X sky130_fd_sc_hd__buf_4
X_7020_ _7022_/CLK _7020_/D vssd1 vssd1 vccd1 vccd1 _7020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4232_ _4232_/A vssd1 vssd1 vccd1 vccd1 _6666_/D sky130_fd_sc_hd__clkbuf_1
X_5447__293 _5447__293/A vssd1 vssd1 vccd1 vccd1 _6583_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4163_ _4163_/A vssd1 vssd1 vccd1 vccd1 _6698_/D sky130_fd_sc_hd__clkbuf_1
X_4094_ _4094_/A vssd1 vssd1 vccd1 vccd1 _6727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2863_ _5797_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2863_/X sky130_fd_sc_hd__clkbuf_16
X_6804_ _6804_/CLK _6804_/D vssd1 vssd1 vccd1 vccd1 _6804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4996_ _4996_/A vssd1 vssd1 vccd1 vccd1 _4996_/X sky130_fd_sc_hd__clkbuf_1
X_3947_ _3947_/A vssd1 vssd1 vccd1 vccd1 _5774_/C sky130_fd_sc_hd__buf_4
XFILLER_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6735_ _6735_/CLK _6735_/D vssd1 vssd1 vccd1 vccd1 _6735_/Q sky130_fd_sc_hd__dfxtp_1
X_5489__327 _5491__329/A vssd1 vssd1 vccd1 vccd1 _6617_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5682__417 _5682__417/A vssd1 vssd1 vccd1 vccd1 _6711_/CLK sky130_fd_sc_hd__inv_2
X_3878_ _6802_/Q _3877_/X _3887_/S vssd1 vssd1 vccd1 vccd1 _3879_/A sky130_fd_sc_hd__mux2_1
X_6666_ _6666_/CLK _6666_/D vssd1 vssd1 vccd1 vccd1 _6666_/Q sky130_fd_sc_hd__dfxtp_1
X_5617_ _5664_/A _5620_/A _5664_/C _5617_/D vssd1 vssd1 vccd1 vccd1 _5892_/B sky130_fd_sc_hd__or4_4
X_6597_ _6597_/CLK _6597_/D vssd1 vssd1 vccd1 vccd1 _6597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5548_ _5548_/A vssd1 vssd1 vccd1 vccd1 _5548_/X sky130_fd_sc_hd__buf_1
XFILLER_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5838__523 _5839__524/A vssd1 vssd1 vccd1 vccd1 _6829_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7149_ _7149_/A vssd1 vssd1 vccd1 vccd1 _7149_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5223__273 _5223__273/A vssd1 vssd1 vccd1 vccd1 _6555_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4850_ _6783_/Q _3986_/A _4849_/X _4806_/A vssd1 vssd1 vccd1 vccd1 _4850_/X sky130_fd_sc_hd__o211a_1
X_3801_ _3696_/X _6831_/Q _3801_/S vssd1 vssd1 vccd1 vccd1 _3802_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6520_ _6520_/CLK _6520_/D vssd1 vssd1 vccd1 vccd1 _6520_/Q sky130_fd_sc_hd__dfxtp_1
X_4781_ _4804_/A _4781_/B vssd1 vssd1 vccd1 vccd1 _4781_/X sky130_fd_sc_hd__or2_1
X_3732_ _3687_/X _6858_/Q _3738_/S vssd1 vssd1 vccd1 vccd1 _3733_/A sky130_fd_sc_hd__mux2_1
X_3663_ _3678_/S vssd1 vssd1 vccd1 vccd1 _3672_/S sky130_fd_sc_hd__buf_2
X_6451_ _6750_/CLK _6451_/D vssd1 vssd1 vccd1 vccd1 _6451_/Q sky130_fd_sc_hd__dfxtp_1
X_6353__38 _6354__39/A vssd1 vssd1 vccd1 vccd1 _7058_/CLK sky130_fd_sc_hd__inv_2
X_6382_ _7141_/A _6381_/B _6381_/Y _6389_/A vssd1 vssd1 vccd1 vccd1 _7080_/D sky130_fd_sc_hd__o211a_1
X_5402_ _5289_/X _5401_/X _5292_/X vssd1 vssd1 vccd1 vccd1 _5402_/Y sky130_fd_sc_hd__o21ai_1
X_3594_ _3594_/A vssd1 vssd1 vccd1 vccd1 _6931_/D sky130_fd_sc_hd__clkbuf_1
X_5333_ _5327_/X _5332_/X _5394_/S vssd1 vssd1 vccd1 vccd1 _5333_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5264_ _5264_/A vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7003_ _7011_/CLK _7003_/D vssd1 vssd1 vccd1 vccd1 _7003_/Q sky130_fd_sc_hd__dfxtp_1
X_4215_ _6673_/Q _4155_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__mux2_1
X_4146_ _7029_/Q vssd1 vssd1 vccd1 vccd1 _4146_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4077_ _4077_/A vssd1 vssd1 vccd1 vccd1 _6733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__2878_ clkbuf_0__2878_/X vssd1 vssd1 vccd1 vccd1 _5876__73/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124__193 _5125__194/A vssd1 vssd1 vccd1 vccd1 _6475_/CLK sky130_fd_sc_hd__inv_2
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4979_ _4973_/X input6/X _4970_/X _4978_/X vssd1 vssd1 vccd1 vccd1 _4979_/X sky130_fd_sc_hd__a22o_2
X_6718_ _6718_/CLK _6718_/D vssd1 vssd1 vccd1 vccd1 _6718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6649_ _6649_/CLK _6649_/D vssd1 vssd1 vccd1 vccd1 _6649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5166__227 _5166__227/A vssd1 vssd1 vccd1 vccd1 _6509_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2528_ clkbuf_0__2528_/X vssd1 vssd1 vccd1 vccd1 _5218__269/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4000_ _4000_/A vssd1 vssd1 vccd1 vccd1 _6763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5951_ _6873_/Q _5951_/B _5951_/C _6870_/Q vssd1 vssd1 vccd1 vccd1 _5961_/C sky130_fd_sc_hd__and4_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__2732_ clkbuf_0__2732_/X vssd1 vssd1 vccd1 vccd1 _5485__324/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4902_ _6547_/Q _6727_/Q _6865_/Q _6531_/Q _4728_/X _4701_/X vssd1 vssd1 vccd1 vccd1
+ _4902_/X sky130_fd_sc_hd__mux4_2
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4833_ _4691_/X input25/X _4832_/X vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__a21o_2
XFILLER_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4764_ _4760_/X _4763_/X _4695_/A vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__o21a_1
X_6503_ _6503_/CLK _6503_/D vssd1 vssd1 vccd1 vccd1 _6503_/Q sky130_fd_sc_hd__dfxtp_1
X_3715_ _3690_/X _6865_/Q _3719_/S vssd1 vssd1 vccd1 vccd1 _3716_/A sky130_fd_sc_hd__mux2_1
X_6326__16 _6328__18/A vssd1 vssd1 vccd1 vccd1 _7036_/CLK sky130_fd_sc_hd__inv_2
X_6434_ _6434_/A vssd1 vssd1 vccd1 vccd1 _7096_/D sky130_fd_sc_hd__clkbuf_1
X_4695_ _4695_/A vssd1 vssd1 vccd1 vccd1 _4695_/X sky130_fd_sc_hd__clkbuf_2
X_3646_ _3646_/A vssd1 vssd1 vccd1 vccd1 _6913_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3577_ _3392_/X _6938_/Q _3577_/S vssd1 vssd1 vccd1 vccd1 _3578_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6296_ _7020_/Q _6300_/B vssd1 vssd1 vccd1 vccd1 _6296_/X sky130_fd_sc_hd__or2_1
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5316_ _6639_/Q _6631_/Q _6615_/Q _6607_/Q _5330_/A _5312_/X vssd1 vssd1 vccd1 vccd1
+ _5316_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4129_ _6711_/Q _3880_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3500_ _3500_/A vssd1 vssd1 vccd1 vccd1 _6972_/D sky130_fd_sc_hd__clkbuf_1
X_4480_ _4480_/A vssd1 vssd1 vccd1 vccd1 _6549_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3000_ clkbuf_0__3000_/X vssd1 vssd1 vccd1 vccd1 _6043__96/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__3154_ clkbuf_0__3154_/X vssd1 vssd1 vccd1 vccd1 _6367_/A sky130_fd_sc_hd__clkbuf_16
X_3431_ _3384_/X _7033_/Q _3435_/S vssd1 vssd1 vccd1 vccd1 _3432_/A sky130_fd_sc_hd__mux2_1
X_3362_ _4036_/A _4044_/B vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__nand2_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5101_/A vssd1 vssd1 vccd1 vccd1 _6466_/D sky130_fd_sc_hd__clkbuf_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3293_ _6748_/Q vssd1 vssd1 vccd1 vccd1 _4009_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_97_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6883_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6983_ _6983_/CLK _6983_/D vssd1 vssd1 vccd1 vccd1 _6983_/Q sky130_fd_sc_hd__dfxtp_1
X_5934_ _6870_/Q vssd1 vssd1 vccd1 vccd1 _5945_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4816_ _6891_/Q _6520_/Q _4876_/A vssd1 vssd1 vccd1 vccd1 _4816_/X sky130_fd_sc_hd__mux2_1
X_4747_ _4752_/B _4747_/B vssd1 vssd1 vccd1 vccd1 _4754_/B sky130_fd_sc_hd__or2_1
X_6104__145 _6104__145/A vssd1 vssd1 vccd1 vccd1 _6953_/CLK sky130_fd_sc_hd__inv_2
X_4678_ _3868_/X _6436_/Q _4678_/S vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6417_ _6417_/A vssd1 vssd1 vccd1 vccd1 _7090_/D sky130_fd_sc_hd__clkbuf_1
X_3629_ _3372_/X _6919_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _3630_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__2862_ clkbuf_0__2862_/X vssd1 vssd1 vccd1 vccd1 _5796__489/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6279_ _7013_/Q _6276_/A _6278_/X _6192_/X vssd1 vssd1 vccd1 vccd1 _7013_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput105 wbs_stb_i vssd1 vssd1 vccd1 vccd1 _5050_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5540__368 _5541__369/A vssd1 vssd1 vccd1 vccd1 _6658_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5179__237 _5179__237/A vssd1 vssd1 vccd1 vccd1 _6519_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3980_ _3977_/A _3977_/B _5723_/B vssd1 vssd1 vccd1 vccd1 _3981_/B sky130_fd_sc_hd__o21ai_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5650_ _7094_/Q _6997_/Q vssd1 vssd1 vccd1 vccd1 _6174_/A sky130_fd_sc_hd__xnor2_1
XFILLER_31_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4601_ _4601_/A vssd1 vssd1 vccd1 vccd1 _6497_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4532_ _4493_/X _6528_/Q _4536_/S vssd1 vssd1 vccd1 vccd1 _4533_/A sky130_fd_sc_hd__mux2_1
X_4463_ _4463_/A vssd1 vssd1 vccd1 vccd1 _6556_/D sky130_fd_sc_hd__clkbuf_1
X_6202_ _6997_/Q vssd1 vssd1 vccd1 vccd1 _6216_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3414_ _3349_/X _7040_/Q _3416_/S vssd1 vssd1 vccd1 vccd1 _3415_/A sky130_fd_sc_hd__mux2_1
X_4394_ _3257_/X _6594_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3345_ _4026_/A vssd1 vssd1 vccd1 vccd1 _3345_/X sky130_fd_sc_hd__buf_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3276_ _3291_/S vssd1 vssd1 vccd1 vccd1 _3285_/S sky130_fd_sc_hd__clkbuf_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5015_/A vssd1 vssd1 vccd1 vccd1 _5015_/X sky130_fd_sc_hd__clkbuf_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5832__518 _5833__519/A vssd1 vssd1 vccd1 vccd1 _6824_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6966_ _6966_/CLK _6966_/D vssd1 vssd1 vccd1 vccd1 _6966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5917_ _6876_/Q _5917_/B _5917_/C vssd1 vssd1 vccd1 vccd1 _5917_/X sky130_fd_sc_hd__and3_1
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6897_ _6897_/CLK _6897_/D vssd1 vssd1 vccd1 vccd1 _6897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2528_ _5213_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2528_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6820_ _6820_/CLK _6820_/D vssd1 vssd1 vccd1 vccd1 _6820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6751_ _6751_/CLK _6751_/D vssd1 vssd1 vccd1 vccd1 _6751_/Q sky130_fd_sc_hd__dfxtp_1
X_3963_ _6767_/Q vssd1 vssd1 vccd1 vccd1 _4868_/S sky130_fd_sc_hd__buf_2
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3894_ _3894_/A vssd1 vssd1 vccd1 vccd1 _6797_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_6682_ _6682_/CLK _6682_/D vssd1 vssd1 vccd1 vccd1 _6682_/Q sky130_fd_sc_hd__dfxtp_1
X_5788__483 _5789__484/A vssd1 vssd1 vccd1 vccd1 _6789_/CLK sky130_fd_sc_hd__inv_2
X_5633_ _4885_/X _5906_/B _5918_/B vssd1 vssd1 vccd1 vccd1 _5908_/B sky130_fd_sc_hd__a21oi_2
XFILLER_117_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4515_ _4515_/A vssd1 vssd1 vccd1 vccd1 _6536_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4446_ _4017_/X _6563_/Q _4450_/S vssd1 vssd1 vccd1 vccd1 _4447_/A sky130_fd_sc_hd__mux2_1
X_4377_ _4377_/A vssd1 vssd1 vccd1 vccd1 _6602_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3328_ _6747_/Q vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6116_ _6140_/A vssd1 vssd1 vccd1 vccd1 _6116_/X sky130_fd_sc_hd__buf_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7096_ _7096_/CLK _7096_/D vssd1 vssd1 vccd1 vccd1 _7096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6047_ _6047_/A vssd1 vssd1 vccd1 vccd1 _6047_/X sky130_fd_sc_hd__buf_1
XFILLER_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3259_ _3259_/A vssd1 vssd1 vccd1 vccd1 _7075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6949_ _6949_/CLK _6949_/D vssd1 vssd1 vccd1 vccd1 _6949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6117__155 _6119__157/A vssd1 vssd1 vccd1 vccd1 _6963_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6083__129 _6083__129/A vssd1 vssd1 vccd1 vccd1 _6937_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput206 _4968_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4300_ _3770_/X _6636_/Q _4306_/S vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5280_ _5286_/A vssd1 vssd1 vccd1 vccd1 _5351_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ _3776_/X _6666_/Q _4233_/S vssd1 vssd1 vccd1 vccd1 _4232_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4162_ _6698_/Q _4161_/X _4165_/S vssd1 vssd1 vccd1 vccd1 _4163_/A sky130_fd_sc_hd__mux2_1
X_4093_ _4017_/X _6727_/Q _4097_/S vssd1 vssd1 vccd1 vccd1 _4094_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6803_ _6803_/CLK _6803_/D vssd1 vssd1 vccd1 vccd1 _6803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4995_ _5003_/A _4995_/B vssd1 vssd1 vccd1 vccd1 _4996_/A sky130_fd_sc_hd__and2_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2862_ _5791_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2862_/X sky130_fd_sc_hd__clkbuf_16
X_3946_ _5776_/A _3946_/B _3946_/C vssd1 vssd1 vccd1 vccd1 _6773_/D sky130_fd_sc_hd__nor3_1
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6734_ _6734_/CLK _6734_/D vssd1 vssd1 vccd1 vccd1 _6734_/Q sky130_fd_sc_hd__dfxtp_2
X_3877_ _6747_/Q vssd1 vssd1 vccd1 vccd1 _3877_/X sky130_fd_sc_hd__clkbuf_4
X_6665_ _6665_/CLK _6665_/D vssd1 vssd1 vccd1 vccd1 _6665_/Q sky130_fd_sc_hd__dfxtp_1
X_5616_ _7087_/Q _7086_/Q vssd1 vssd1 vccd1 vccd1 _5617_/D sky130_fd_sc_hd__or2_1
X_6596_ _6596_/CLK _6596_/D vssd1 vssd1 vccd1 vccd1 _6596_/Q sky130_fd_sc_hd__dfxtp_1
X_5762__464 _5762__464/A vssd1 vssd1 vccd1 vccd1 _6768_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4429_ _4429_/A vssd1 vssd1 vccd1 vccd1 _6571_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7148_ _7148_/A vssd1 vssd1 vccd1 vccd1 _7148_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7079_ _7079_/CLK _7079_/D vssd1 vssd1 vccd1 vccd1 _7079_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2757_ clkbuf_0__2757_/X vssd1 vssd1 vccd1 vccd1 _5697_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_77_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4780_ _6543_/Q _6723_/Q _6861_/Q _6527_/Q _4719_/A _4936_/S vssd1 vssd1 vccd1 vccd1
+ _4781_/B sky130_fd_sc_hd__mux4_2
X_3800_ _3800_/A vssd1 vssd1 vccd1 vccd1 _6832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3731_ _3731_/A vssd1 vssd1 vccd1 vccd1 _6859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3662_ _4608_/B _4644_/B vssd1 vssd1 vccd1 vccd1 _3678_/S sky130_fd_sc_hd__or2_2
X_6450_ _6750_/CLK _6450_/D vssd1 vssd1 vccd1 vccd1 _6450_/Q sky130_fd_sc_hd__dfxtp_1
X_6381_ _6381_/A _6381_/B vssd1 vssd1 vccd1 vccd1 _6381_/Y sky130_fd_sc_hd__nand2_1
X_5401_ _6959_/Q _6943_/Q _7068_/Q _6935_/Q _5266_/X _5268_/X vssd1 vssd1 vccd1 vccd1
+ _5401_/X sky130_fd_sc_hd__mux4_2
X_3593_ _6931_/Q _3459_/X _3595_/S vssd1 vssd1 vccd1 vccd1 _3594_/A sky130_fd_sc_hd__mux2_1
X_5332_ _5328_/X _5331_/X _5429_/S vssd1 vssd1 vccd1 vccd1 _5332_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5263_ _5337_/A vssd1 vssd1 vccd1 vccd1 _5263_/X sky130_fd_sc_hd__clkbuf_4
X_5194_ _5200_/A vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__buf_1
X_7002_ _7011_/CLK _7002_/D vssd1 vssd1 vccd1 vccd1 _7002_/Q sky130_fd_sc_hd__dfxtp_1
X_4214_ _4214_/A vssd1 vssd1 vccd1 vccd1 _6674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4145_ _4145_/A vssd1 vssd1 vccd1 vccd1 _6704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5495__332 _5497__334/A vssd1 vssd1 vccd1 vccd1 _6622_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4076_ _4071_/X _4076_/B _6318_/B vssd1 vssd1 vccd1 vccd1 _4077_/A sky130_fd_sc_hd__and3b_1
Xclkbuf_1_1_0__2877_ clkbuf_0__2877_/X vssd1 vssd1 vccd1 vccd1 _5871__69/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4978_ _7084_/Q vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6717_ _6717_/CLK _6717_/D vssd1 vssd1 vccd1 vccd1 _6717_/Q sky130_fd_sc_hd__dfxtp_1
X_3929_ _3929_/A vssd1 vssd1 vccd1 vccd1 _6782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6648_ _6648_/CLK _6648_/D vssd1 vssd1 vccd1 vccd1 _6648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6579_ _6888_/CLK _6579_/D vssd1 vssd1 vccd1 vccd1 _6579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5504__339 _5504__339/A vssd1 vssd1 vccd1 vccd1 _6629_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2527_ clkbuf_0__2527_/X vssd1 vssd1 vccd1 vccd1 _5212__264/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2458_ clkbuf_0__2458_/X vssd1 vssd1 vccd1 vccd1 _5119__189/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5559__384 _5559__384/A vssd1 vssd1 vccd1 vccd1 _6674_/CLK sky130_fd_sc_hd__inv_2
X_5950_ _5950_/A vssd1 vssd1 vccd1 vccd1 _6872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2731_ clkbuf_0__2731_/X vssd1 vssd1 vccd1 vccd1 _5478__318/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4901_ _4774_/X _4900_/X _4905_/A vssd1 vssd1 vccd1 vccd1 _4901_/X sky130_fd_sc_hd__a21o_1
XFILLER_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4832_ _5910_/A _4763_/X _4695_/A _4831_/X vssd1 vssd1 vccd1 vccd1 _4832_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4763_ _4798_/A _4798_/B vssd1 vssd1 vccd1 vccd1 _4763_/X sky130_fd_sc_hd__or2_1
XFILLER_119_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6502_ _6502_/CLK _6502_/D vssd1 vssd1 vccd1 vccd1 _6502_/Q sky130_fd_sc_hd__dfxtp_1
X_3714_ _3714_/A vssd1 vssd1 vccd1 vccd1 _6866_/D sky130_fd_sc_hd__clkbuf_1
X_4694_ _4987_/A _6427_/A _5736_/B vssd1 vssd1 vccd1 vccd1 _4695_/A sky130_fd_sc_hd__and3_1
XFILLER_119_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6433_ _6433_/A _6433_/B vssd1 vssd1 vccd1 vccd1 _6434_/A sky130_fd_sc_hd__or2_1
X_3645_ _3294_/X _6913_/Q _3653_/S vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6096__139 _6096__139/A vssd1 vssd1 vccd1 vccd1 _6947_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3576_ _3576_/A vssd1 vssd1 vccd1 vccd1 _6939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6295_ _7020_/Q _6284_/X _6294_/X _6290_/X vssd1 vssd1 vccd1 vccd1 _7019_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5315_ _5313_/X _5314_/X _5439_/B vssd1 vssd1 vccd1 vccd1 _5315_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4128_ _4128_/A vssd1 vssd1 vccd1 vccd1 _6712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4059_ _5286_/A vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5172__232 _5172__232/A vssd1 vssd1 vccd1 vccd1 _6514_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5695__428 _5696__429/A vssd1 vssd1 vccd1 vccd1 _6722_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5782__478 _5783__479/A vssd1 vssd1 vccd1 vccd1 _6784_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3430_ _3430_/A vssd1 vssd1 vccd1 vccd1 _7034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6331__20 _6334__23/A vssd1 vssd1 vccd1 vccd1 _7040_/CLK sky130_fd_sc_hd__inv_2
X_3361_ _3361_/A _4051_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _4044_/B sky130_fd_sc_hd__and3_2
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5100_ _6466_/Q _7120_/A _5586_/S vssd1 vssd1 vccd1 vccd1 _5101_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3292_ _3292_/A vssd1 vssd1 vccd1 vccd1 _7063_/D sky130_fd_sc_hd__clkbuf_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6982_ _6982_/CLK _6982_/D vssd1 vssd1 vccd1 vccd1 _6982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5933_ _5933_/A vssd1 vssd1 vccd1 vccd1 _6869_/D sky130_fd_sc_hd__clkbuf_1
X_4815_ _3986_/X _6512_/Q _4814_/X _4719_/X vssd1 vssd1 vccd1 vccd1 _4815_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5236__284 _5236__284/A vssd1 vssd1 vccd1 vccd1 _6566_/CLK sky130_fd_sc_hd__inv_2
XFILLER_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4746_ _4795_/A _4762_/D _4693_/A vssd1 vssd1 vccd1 vccd1 _4747_/B sky130_fd_sc_hd__o21a_1
X_4677_ _4677_/A vssd1 vssd1 vccd1 vccd1 _6437_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2861_ clkbuf_0__2861_/X vssd1 vssd1 vccd1 vccd1 _5815_/A sky130_fd_sc_hd__clkbuf_4
X_6416_ _6430_/A _6416_/B vssd1 vssd1 vccd1 vccd1 _6417_/A sky130_fd_sc_hd__or2_1
X_3628_ _3628_/A vssd1 vssd1 vccd1 vccd1 _6920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3559_ _6946_/Q _3462_/X _3559_/S vssd1 vssd1 vccd1 vccd1 _3560_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6278_ _6995_/Q _6277_/Y _6272_/B _6271_/X _6272_/A vssd1 vssd1 vccd1 vccd1 _6278_/X
+ sky130_fd_sc_hd__a2111o_1
Xinput106 wbs_we_i vssd1 vssd1 vccd1 vccd1 _7161_/A sky130_fd_sc_hd__buf_6
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5243__288 _5244__289/A vssd1 vssd1 vccd1 vccd1 _6570_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_79_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4600_ _6497_/Q _4023_/A _4600_/S vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4531_ _4531_/A vssd1 vssd1 vccd1 vccd1 _6529_/D sky130_fd_sc_hd__clkbuf_1
X_4462_ _4014_/X _6556_/Q _4468_/S vssd1 vssd1 vccd1 vccd1 _4463_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6201_ _6229_/C vssd1 vssd1 vccd1 vccd1 _6238_/A sky130_fd_sc_hd__clkbuf_2
X_3413_ _3413_/A vssd1 vssd1 vccd1 vccd1 _7041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4393_ _4393_/A vssd1 vssd1 vccd1 vccd1 _6595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3344_ _6743_/Q vssd1 vssd1 vccd1 vccd1 _4026_/A sky130_fd_sc_hd__buf_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3275_ _3579_/A _4186_/A vssd1 vssd1 vccd1 vccd1 _3291_/S sky130_fd_sc_hd__nor2_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5014_ _5014_/A _5014_/B vssd1 vssd1 vccd1 vccd1 _5015_/A sky130_fd_sc_hd__and2_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6110__150 _6113__153/A vssd1 vssd1 vccd1 vccd1 _6958_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6965_ _6965_/CLK _6965_/D vssd1 vssd1 vccd1 vccd1 _6965_/Q sky130_fd_sc_hd__dfxtp_1
X_5916_ _5915_/B _5915_/C _6875_/Q vssd1 vssd1 vccd1 vccd1 _5916_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6896_ _6896_/CLK _6896_/D vssd1 vssd1 vccd1 vccd1 _6896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5778_ _5778_/A vssd1 vssd1 vccd1 vccd1 _5778_/X sky130_fd_sc_hd__buf_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4729_ _6478_/Q _6550_/Q _7039_/Q _6970_/Q _4701_/A _4728_/X vssd1 vssd1 vccd1 vccd1
+ _4729_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_0__2527_ _5207_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2527_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__2458_ _5037_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2458_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5185__242 _5186__243/A vssd1 vssd1 vccd1 vccd1 _6524_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6750_ _6750_/CLK _6750_/D vssd1 vssd1 vccd1 vccd1 _6750_/Q sky130_fd_sc_hd__dfxtp_1
X_3962_ _3962_/A _3962_/B _3309_/X vssd1 vssd1 vccd1 vccd1 _3983_/B sky130_fd_sc_hd__or3b_1
XFILLER_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3893_ _6797_/Q _3892_/X _3896_/S vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__mux2_1
X_6681_ _6681_/CLK _6681_/D vssd1 vssd1 vccd1 vccd1 _6681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5632_ _5648_/A _5910_/A _6173_/A _7092_/Q vssd1 vssd1 vccd1 vccd1 _5918_/B sky130_fd_sc_hd__nor4_2
X_4514_ _4493_/X _6536_/Q _4518_/S vssd1 vssd1 vccd1 vccd1 _4515_/A sky130_fd_sc_hd__mux2_1
X_4445_ _4445_/A vssd1 vssd1 vccd1 vccd1 _6564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4376_ _6602_/Q _3776_/A _4378_/S vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3327_ _3327_/A vssd1 vssd1 vccd1 vccd1 _7062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6115_ _6115_/A vssd1 vssd1 vccd1 vccd1 _6115_/X sky130_fd_sc_hd__buf_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7095_ _7095_/CLK _7095_/D vssd1 vssd1 vccd1 vccd1 _7095_/Q sky130_fd_sc_hd__dfxtp_1
X_5795__488 _5795__488/A vssd1 vssd1 vccd1 vccd1 _6794_/CLK sky130_fd_sc_hd__inv_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5459__303 _5460__304/A vssd1 vssd1 vccd1 vccd1 _6593_/CLK sky130_fd_sc_hd__inv_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _7075_/Q _3257_/X _3261_/S vssd1 vssd1 vccd1 vccd1 _3259_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6948_ _6948_/CLK _6948_/D vssd1 vssd1 vccd1 vccd1 _6948_/Q sky130_fd_sc_hd__dfxtp_1
X_6879_ _6883_/CLK _6879_/D vssd1 vssd1 vccd1 vccd1 _6879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2758_ clkbuf_0__2758_/X vssd1 vssd1 vccd1 vccd1 _5601__411/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5553__379 _5553__379/A vssd1 vssd1 vccd1 vccd1 _6669_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6365__48 _6366__49/A vssd1 vssd1 vccd1 vccd1 _7068_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput207 _4972_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_4_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4230_ _4230_/A vssd1 vssd1 vccd1 vccd1 _6667_/D sky130_fd_sc_hd__clkbuf_1
X_4161_ _7024_/Q vssd1 vssd1 vccd1 vccd1 _4161_/X sky130_fd_sc_hd__buf_2
XFILLER_68_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4092_ _4092_/A vssd1 vssd1 vccd1 vccd1 _6728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6802_ _6802_/CLK _6802_/D vssd1 vssd1 vccd1 vccd1 _6802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2861_ _5790_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2861_/X sky130_fd_sc_hd__clkbuf_16
X_4994_ _5005_/A vssd1 vssd1 vccd1 vccd1 _5003_/A sky130_fd_sc_hd__clkbuf_1
X_3945_ _3948_/A _3948_/B _3661_/A vssd1 vssd1 vccd1 vccd1 _3946_/C sky130_fd_sc_hd__a21oi_1
X_5454__299 _5454__299/A vssd1 vssd1 vccd1 vccd1 _6589_/CLK sky130_fd_sc_hd__inv_2
X_6733_ _6733_/CLK _6733_/D vssd1 vssd1 vccd1 vccd1 _6733_/Q sky130_fd_sc_hd__dfxtp_1
X_6664_ _6664_/CLK _6664_/D vssd1 vssd1 vccd1 vccd1 _6664_/Q sky130_fd_sc_hd__dfxtp_1
X_3876_ _3876_/A vssd1 vssd1 vccd1 vccd1 _6803_/D sky130_fd_sc_hd__clkbuf_1
X_5615_ _7009_/Q _5609_/Y _5610_/X _7011_/Q _5614_/X vssd1 vssd1 vccd1 vccd1 _5669_/A
+ sky130_fd_sc_hd__a221o_1
X_6595_ _6595_/CLK _6595_/D vssd1 vssd1 vccd1 vccd1 _6595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4428_ _3254_/X _6571_/Q _4432_/S vssd1 vssd1 vccd1 vccd1 _4429_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7147_ _7147_/A vssd1 vssd1 vccd1 vccd1 _7147_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4359_ _4359_/A vssd1 vssd1 vccd1 vccd1 _6610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7078_ _7078_/CLK _7078_/D vssd1 vssd1 vccd1 vccd1 _7078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5136__203 _5136__203/A vssd1 vssd1 vccd1 vccd1 _6485_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5845__529 _5845__529/A vssd1 vssd1 vccd1 vccd1 _6835_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6123__160 _6124__161/A vssd1 vssd1 vccd1 vccd1 _6968_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5858__58 _5859__59/A vssd1 vssd1 vccd1 vccd1 _6844_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _3680_/X _6859_/Q _3738_/S vssd1 vssd1 vccd1 vccd1 _3731_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6338__26 _6338__26/A vssd1 vssd1 vccd1 vccd1 _7046_/CLK sky130_fd_sc_hd__inv_2
X_3661_ _3661_/A _3948_/A _3661_/C vssd1 vssd1 vccd1 vccd1 _4644_/B sky130_fd_sc_hd__or3_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6380_ _7142_/A _6381_/B _6379_/X _6389_/A vssd1 vssd1 vccd1 vccd1 _7079_/D sky130_fd_sc_hd__o211a_1
X_3592_ _3592_/A vssd1 vssd1 vccd1 vccd1 _6932_/D sky130_fd_sc_hd__clkbuf_1
X_5400_ _5399_/X _5439_/B vssd1 vssd1 vccd1 vccd1 _5400_/X sky130_fd_sc_hd__and2b_1
XFILLER_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5230__279 _5230__279/A vssd1 vssd1 vccd1 vccd1 _6561_/CLK sky130_fd_sc_hd__inv_2
X_5331_ _6600_/Q _6584_/Q _6838_/Q _6822_/Q _5329_/X _5330_/X vssd1 vssd1 vccd1 vccd1
+ _5331_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7001_ _7019_/CLK _7001_/D vssd1 vssd1 vccd1 vccd1 _7001_/Q sky130_fd_sc_hd__dfxtp_1
X_5262_ _5255_/X _5260_/X _5410_/S vssd1 vssd1 vccd1 vccd1 _5262_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4213_ _6674_/Q _4152_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4214_/A sky130_fd_sc_hd__mux2_1
X_4144_ _6704_/Q _4141_/X _4156_/S vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4075_ _6305_/A vssd1 vssd1 vccd1 vccd1 _6318_/B sky130_fd_sc_hd__buf_2
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2876_ clkbuf_0__2876_/X vssd1 vssd1 vccd1 vccd1 _5865__64/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6716_ _6716_/CLK _6716_/D vssd1 vssd1 vccd1 vccd1 _6716_/Q sky130_fd_sc_hd__dfxtp_1
X_4977_ _4973_/X input5/X _4970_/X _5892_/A vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__a22o_2
X_3928_ _6782_/Q _3889_/X _3932_/S vssd1 vssd1 vccd1 vccd1 _3929_/A sky130_fd_sc_hd__mux2_1
X_3859_ _6744_/Q vssd1 vssd1 vccd1 vccd1 _3859_/X sky130_fd_sc_hd__buf_4
X_6647_ _6647_/CLK _6647_/D vssd1 vssd1 vccd1 vccd1 _6647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6578_ _6888_/CLK _6578_/D vssd1 vssd1 vccd1 vccd1 _6578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5529_ _5529_/A vssd1 vssd1 vccd1 vccd1 _5529_/X sky130_fd_sc_hd__buf_1
X_5131__199 _5131__199/A vssd1 vssd1 vccd1 vccd1 _6481_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2526_ clkbuf_0__2526_/X vssd1 vssd1 vccd1 vccd1 _5231_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2457_ clkbuf_0__2457_/X vssd1 vssd1 vccd1 vccd1 _5138_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6040__94 _6040__94/A vssd1 vssd1 vccd1 vccd1 _6902_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3009_ clkbuf_0__3009_/X vssd1 vssd1 vccd1 vccd1 _6090__134/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2730_ clkbuf_0__2730_/X vssd1 vssd1 vccd1 vccd1 _5470__311/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _6894_/Q _6523_/Q _4900_/S vssd1 vssd1 vccd1 vccd1 _4900_/X sky130_fd_sc_hd__mux2_2
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4831_ _6777_/Q _4766_/Y _4820_/X _4830_/Y _4798_/Y vssd1 vssd1 vccd1 vccd1 _4831_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4762_ _4795_/A _4795_/B _4762_/C _4762_/D vssd1 vssd1 vccd1 vccd1 _4798_/B sky130_fd_sc_hd__or4_1
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3713_ _3687_/X _6866_/Q _3719_/S vssd1 vssd1 vccd1 vccd1 _3714_/A sky130_fd_sc_hd__mux2_1
X_6501_ _6501_/CLK _6501_/D vssd1 vssd1 vccd1 vccd1 _6501_/Q sky130_fd_sc_hd__dfxtp_1
X_4693_ _4693_/A vssd1 vssd1 vccd1 vccd1 _5736_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3644_ _3659_/S vssd1 vssd1 vccd1 vccd1 _3653_/S sky130_fd_sc_hd__clkbuf_2
X_6432_ _7125_/A _7096_/Q _6432_/S vssd1 vssd1 vccd1 vccd1 _6433_/B sky130_fd_sc_hd__mux2_1
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5566__389 _5566__389/A vssd1 vssd1 vccd1 vccd1 _6679_/CLK sky130_fd_sc_hd__inv_2
X_3575_ _3388_/X _6939_/Q _3577_/S vssd1 vssd1 vccd1 vccd1 _3576_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6294_ _7019_/Q _6300_/B vssd1 vssd1 vccd1 vccd1 _6294_/X sky130_fd_sc_hd__or2_1
X_5314_ _6671_/Q _6663_/Q _6655_/Q _6647_/Q _5311_/X _5312_/X vssd1 vssd1 vccd1 vccd1
+ _5314_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5245_ _5449_/A vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__buf_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5176_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5176_/X sky130_fd_sc_hd__buf_1
XFILLER_110_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4127_ _6712_/Q _3877_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4128_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4058_ _5302_/A vssd1 vssd1 vccd1 vccd1 _5286_/A sky130_fd_sc_hd__buf_2
XFILLER_44_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__2859_ clkbuf_0__2859_/X vssd1 vssd1 vccd1 vccd1 _5783__479/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_24_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__2758_ _5599_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2758_/X sky130_fd_sc_hd__clkbuf_16
X_5510__344 _5510__344/A vssd1 vssd1 vccd1 vccd1 _6634_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5149__213 _5150__214/A vssd1 vssd1 vccd1 vccd1 _6495_/CLK sky130_fd_sc_hd__inv_2
X_3360_ _3623_/B vssd1 vssd1 vccd1 vccd1 _4040_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5030_ _5030_/A vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__buf_1
X_3291_ _7063_/Q _3269_/X _3291_/S vssd1 vssd1 vccd1 vccd1 _3292_/A sky130_fd_sc_hd__mux2_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6981_ _6981_/CLK _6981_/D vssd1 vssd1 vccd1 vccd1 _6981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2867_ clkbuf_0__2867_/X vssd1 vssd1 vccd1 vccd1 _5846_/A sky130_fd_sc_hd__clkbuf_16
X_5932_ _5954_/B _6019_/B _5932_/C vssd1 vssd1 vccd1 vccd1 _5933_/A sky130_fd_sc_hd__and3b_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4814_ _4814_/A _6496_/Q vssd1 vssd1 vccd1 vccd1 _4814_/X sky130_fd_sc_hd__or2_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4745_ _6445_/Q _6453_/Q _6454_/Q vssd1 vssd1 vccd1 vccd1 _4762_/D sky130_fd_sc_hd__or3_1
XFILLER_119_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4676_ _3865_/X _6437_/Q _4678_/S vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__mux2_1
X_6415_ _7131_/A _7090_/Q _6432_/S vssd1 vssd1 vccd1 vccd1 _6416_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__2860_ clkbuf_0__2860_/X vssd1 vssd1 vccd1 vccd1 _5789__484/A sky130_fd_sc_hd__clkbuf_4
X_3627_ _3368_/X _6920_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _3628_/A sky130_fd_sc_hd__mux2_1
X_3558_ _3558_/A vssd1 vssd1 vccd1 vccd1 _6947_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6277_ _7013_/Q _7012_/Q vssd1 vssd1 vccd1 vccd1 _6277_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3489_ _3294_/X _6977_/Q _3497_/S vssd1 vssd1 vccd1 vccd1 _3490_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4530_ _4490_/X _6529_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4461_ _4461_/A vssd1 vssd1 vccd1 vccd1 _6557_/D sky130_fd_sc_hd__clkbuf_1
X_6200_ _6270_/A _6282_/A vssd1 vssd1 vccd1 vccd1 _6229_/C sky130_fd_sc_hd__nor2_2
X_3412_ _3345_/X _7041_/Q _3416_/S vssd1 vssd1 vccd1 vccd1 _3413_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4392_ _3254_/X _6595_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4393_/A sky130_fd_sc_hd__mux2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3343_ _3343_/A vssd1 vssd1 vccd1 vccd1 _7058_/D sky130_fd_sc_hd__clkbuf_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3274_ _4296_/A vssd1 vssd1 vccd1 vccd1 _4186_/A sky130_fd_sc_hd__clkbuf_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5013_ _5013_/A vssd1 vssd1 vccd1 vccd1 _5013_/X sky130_fd_sc_hd__clkbuf_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6964_ _6964_/CLK _6964_/D vssd1 vssd1 vccd1 vccd1 _6964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6895_ _6895_/CLK _6895_/D vssd1 vssd1 vccd1 vccd1 _6895_/Q sky130_fd_sc_hd__dfxtp_1
X_5915_ _6875_/Q _5915_/B _5915_/C vssd1 vssd1 vccd1 vccd1 _5915_/X sky130_fd_sc_hd__or3_1
XFILLER_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5846_ _5846_/A vssd1 vssd1 vccd1 vccd1 _5846_/X sky130_fd_sc_hd__buf_1
XFILLER_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4728_ _4906_/A vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__buf_6
Xclkbuf_0__2526_ _5206_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2526_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4659_ _4659_/A vssd1 vssd1 vccd1 vccd1 _6471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2457_ _5036_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2457_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_115_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3009_ _6085_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3009_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3961_ _3961_/A _3961_/B vssd1 vssd1 vccd1 vccd1 _3962_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3892_ _6742_/Q vssd1 vssd1 vccd1 vccd1 _3892_/X sky130_fd_sc_hd__buf_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6680_ _6680_/CLK _6680_/D vssd1 vssd1 vccd1 vccd1 _6680_/Q sky130_fd_sc_hd__dfxtp_1
X_5631_ _5648_/A _7094_/Q _7093_/Q vssd1 vssd1 vccd1 vccd1 _5906_/B sky130_fd_sc_hd__or3_2
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4513_ _4513_/A vssd1 vssd1 vccd1 vccd1 _6537_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4444_ _4014_/X _6564_/Q _4450_/S vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__mux2_1
X_4375_ _4375_/A vssd1 vssd1 vccd1 vccd1 _6603_/D sky130_fd_sc_hd__clkbuf_1
X_3326_ _3294_/X _7062_/Q _3342_/S vssd1 vssd1 vccd1 vccd1 _3327_/A sky130_fd_sc_hd__mux2_1
X_7094_ _7095_/CLK _7094_/D vssd1 vssd1 vccd1 vccd1 _7094_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _7027_/Q vssd1 vssd1 vccd1 vccd1 _3257_/X sky130_fd_sc_hd__clkbuf_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6947_ _6947_/CLK _6947_/D vssd1 vssd1 vccd1 vccd1 _6947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6878_ _6883_/CLK _6878_/D vssd1 vssd1 vccd1 vccd1 _6878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4160_ _4160_/A vssd1 vssd1 vccd1 vccd1 _6699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4091_ _4014_/X _6728_/Q _4097_/S vssd1 vssd1 vccd1 vccd1 _4092_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6801_ _6801_/CLK _6801_/D vssd1 vssd1 vccd1 vccd1 _6801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__2860_ _5784_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2860_/X sky130_fd_sc_hd__clkbuf_16
X_4993_ _4993_/A vssd1 vssd1 vccd1 vccd1 _4993_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3944_ _3727_/B _3946_/B _3943_/Y vssd1 vssd1 vccd1 vccd1 _6774_/D sky130_fd_sc_hd__o21a_1
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6732_ _6732_/CLK _6732_/D vssd1 vssd1 vccd1 vccd1 _6732_/Q sky130_fd_sc_hd__dfxtp_1
X_3875_ _6803_/Q _3871_/X _3887_/S vssd1 vssd1 vccd1 vccd1 _3876_/A sky130_fd_sc_hd__mux2_1
X_6663_ _6663_/CLK _6663_/D vssd1 vssd1 vccd1 vccd1 _6663_/Q sky130_fd_sc_hd__dfxtp_1
X_5614_ _6269_/A _6266_/A _5888_/C vssd1 vssd1 vccd1 vccd1 _5614_/X sky130_fd_sc_hd__and3_1
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6594_ _6594_/CLK _6594_/D vssd1 vssd1 vccd1 vccd1 _6594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4427_ _4427_/A vssd1 vssd1 vccd1 vccd1 _6572_/D sky130_fd_sc_hd__clkbuf_1
X_7146_ _7146_/A vssd1 vssd1 vccd1 vccd1 _7146_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4358_ _6610_/Q _3776_/A _4360_/S vssd1 vssd1 vccd1 vccd1 _4359_/A sky130_fd_sc_hd__mux2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3309_ _6767_/Q _3315_/D vssd1 vssd1 vccd1 vccd1 _3309_/X sky130_fd_sc_hd__or2b_1
XFILLER_59_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4289_/A vssd1 vssd1 vccd1 vccd1 _6641_/D sky130_fd_sc_hd__clkbuf_1
X_7077_ _7077_/CLK _7077_/D vssd1 vssd1 vccd1 vccd1 _7077_/Q sky130_fd_sc_hd__dfxtp_1
X_6028_ _6028_/A vssd1 vssd1 vccd1 vccd1 _6028_/X sky130_fd_sc_hd__buf_1
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6370__52 _6370__52/A vssd1 vssd1 vccd1 vccd1 _7072_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3660_ _3660_/A vssd1 vssd1 vccd1 vccd1 _6906_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3591_ _6932_/Q _3456_/X _3595_/S vssd1 vssd1 vccd1 vccd1 _3592_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _5330_/A vssd1 vssd1 vccd1 vccd1 _5330_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7096_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_5261_ _5286_/A vssd1 vssd1 vccd1 vccd1 _5410_/S sky130_fd_sc_hd__clkbuf_2
X_7000_ _7093_/CLK _7000_/D vssd1 vssd1 vccd1 vccd1 _7000_/Q sky130_fd_sc_hd__dfxtp_1
X_4212_ _4212_/A vssd1 vssd1 vccd1 vccd1 _6675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4143_ _4165_/S vssd1 vssd1 vccd1 vccd1 _4156_/S sky130_fd_sc_hd__buf_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4074_ _4071_/B _4070_/A _4070_/B _4071_/A vssd1 vssd1 vccd1 vccd1 _4076_/B sky130_fd_sc_hd__a31o_1
XFILLER_95_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5198__253 _5199__254/A vssd1 vssd1 vccd1 vccd1 _6535_/CLK sky130_fd_sc_hd__inv_2
XFILLER_24_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6715_ _6715_/CLK _6715_/D vssd1 vssd1 vccd1 vccd1 _6715_/Q sky130_fd_sc_hd__dfxtp_1
X_4976_ _7085_/Q vssd1 vssd1 vccd1 vccd1 _5892_/A sky130_fd_sc_hd__buf_4
X_3927_ _3927_/A vssd1 vssd1 vccd1 vccd1 _6783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3858_ _3858_/A vssd1 vssd1 vccd1 vccd1 _6808_/D sky130_fd_sc_hd__clkbuf_1
X_6646_ _6646_/CLK _6646_/D vssd1 vssd1 vccd1 vccd1 _6646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3789_ _3788_/X _6836_/Q _3789_/S vssd1 vssd1 vccd1 vccd1 _3790_/A sky130_fd_sc_hd__mux2_1
X_6577_ _6897_/CLK _6577_/D vssd1 vssd1 vccd1 vccd1 _6577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7129_ _7129_/A vssd1 vssd1 vccd1 vccd1 _7129_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2525_ clkbuf_0__2525_/X vssd1 vssd1 vccd1 vccd1 _5205__259/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5863__62 _5865__64/A vssd1 vssd1 vccd1 vccd1 _6848_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5851__534 _5851__534/A vssd1 vssd1 vccd1 vccd1 _6840_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2456_ clkbuf_0__2456_/X vssd1 vssd1 vccd1 vccd1 _5033__182/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3008_ clkbuf_0__3008_/X vssd1 vssd1 vccd1 vccd1 _6109_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5745__450 _5747__452/A vssd1 vssd1 vccd1 vccd1 _6754_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4830_ _4918_/A _4830_/B vssd1 vssd1 vccd1 vccd1 _4830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _5113_/B _4761_/B _4761_/C _4761_/D vssd1 vssd1 vccd1 vccd1 _4795_/B sky130_fd_sc_hd__or4_1
XFILLER_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3712_ _3712_/A vssd1 vssd1 vccd1 vccd1 _6867_/D sky130_fd_sc_hd__clkbuf_1
X_6500_ _6500_/CLK _6500_/D vssd1 vssd1 vccd1 vccd1 _6500_/Q sky130_fd_sc_hd__dfxtp_1
X_4692_ _6694_/Q vssd1 vssd1 vccd1 vccd1 _6427_/A sky130_fd_sc_hd__buf_2
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3643_ _4458_/A _4608_/B vssd1 vssd1 vccd1 vccd1 _3659_/S sky130_fd_sc_hd__or2_2
X_6431_ _6431_/A vssd1 vssd1 vccd1 vccd1 _7095_/D sky130_fd_sc_hd__clkbuf_1
X_3574_ _3574_/A vssd1 vssd1 vccd1 vccd1 _6940_/D sky130_fd_sc_hd__clkbuf_1
X_5313_ _7072_/Q _6698_/Q _6567_/Q _6845_/Q _5311_/X _5312_/X vssd1 vssd1 vccd1 vccd1
+ _5313_/X sky130_fd_sc_hd__mux4_1
X_6293_ _7019_/Q _6284_/X _6292_/X _6290_/X vssd1 vssd1 vccd1 vccd1 _7018_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5175_ _5175_/A vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__buf_1
XFILLER_96_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4126_ _4126_/A vssd1 vssd1 vccd1 vccd1 _6713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4057_ _5334_/A vssd1 vssd1 vccd1 vccd1 _4071_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4959_ _3977_/A _4956_/X _4958_/X vssd1 vssd1 vccd1 vccd1 _4959_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_0__2757_ _5598_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2757_/X sky130_fd_sc_hd__clkbuf_16
X_6629_ _6629_/CLK _6629_/D vssd1 vssd1 vccd1 vccd1 _6629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1__f__2454_ clkbuf_0__2454_/X vssd1 vssd1 vccd1 vccd1 _5175_/A sky130_fd_sc_hd__clkbuf_16
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3290_ _3290_/A vssd1 vssd1 vccd1 vccd1 _7064_/D sky130_fd_sc_hd__clkbuf_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6136__171 _6137__172/A vssd1 vssd1 vccd1 vccd1 _6979_/CLK sky130_fd_sc_hd__inv_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6980_ _6980_/CLK _6980_/D vssd1 vssd1 vccd1 vccd1 _6980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2866_ clkbuf_0__2866_/X vssd1 vssd1 vccd1 vccd1 _5820__509/A sky130_fd_sc_hd__clkbuf_16
X_5931_ _5929_/B _5926_/B _5929_/A vssd1 vssd1 vccd1 vccd1 _5932_/C sky130_fd_sc_hd__o21ai_1
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5572__394 _5572__394/A vssd1 vssd1 vccd1 vccd1 _6684_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4813_ _4851_/S vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__buf_4
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4744_ _6446_/Q vssd1 vssd1 vccd1 vccd1 _4795_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4675_ _4675_/A vssd1 vssd1 vccd1 vccd1 _6438_/D sky130_fd_sc_hd__clkbuf_1
X_6414_ _6414_/A vssd1 vssd1 vccd1 vccd1 _7089_/D sky130_fd_sc_hd__clkbuf_1
X_3626_ _3626_/A vssd1 vssd1 vccd1 vccd1 _6921_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3557_ _6947_/Q _3459_/X _3559_/S vssd1 vssd1 vccd1 vccd1 _3558_/A sky130_fd_sc_hd__mux2_1
X_6276_ _6276_/A _6276_/B vssd1 vssd1 vccd1 vccd1 _7012_/D sky130_fd_sc_hd__nor2_1
XFILLER_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3488_ _3503_/S vssd1 vssd1 vccd1 vccd1 _3497_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _6720_/Q _3877_/X _4115_/S vssd1 vssd1 vccd1 vccd1 _4110_/A sky130_fd_sc_hd__mux2_1
X_5089_ _6461_/Q _7115_/A _5093_/S vssd1 vssd1 vccd1 vccd1 _5090_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6079__125 _6083__129/A vssd1 vssd1 vccd1 vccd1 _6933_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5033__182 _5033__182/A vssd1 vssd1 vccd1 vccd1 _6438_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4460_ _4009_/X _6557_/Q _4468_/S vssd1 vssd1 vccd1 vccd1 _4461_/A sky130_fd_sc_hd__mux2_1
X_3411_ _3411_/A vssd1 vssd1 vccd1 vccd1 _7042_/D sky130_fd_sc_hd__clkbuf_1
X_4391_ _4391_/A vssd1 vssd1 vccd1 vccd1 _6596_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3342_ _3341_/X _7058_/Q _3342_/S vssd1 vssd1 vccd1 vccd1 _3343_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5678__414 _5678__414/A vssd1 vssd1 vccd1 vccd1 _6708_/CLK sky130_fd_sc_hd__inv_2
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3361_/A _3273_/B _3418_/C vssd1 vssd1 vccd1 vccd1 _4296_/A sky130_fd_sc_hd__or3_4
X_5758__460 _5760__462/A vssd1 vssd1 vccd1 vccd1 _6764_/CLK sky130_fd_sc_hd__inv_2
X_5012_ _5014_/A _5012_/B vssd1 vssd1 vccd1 vccd1 _5013_/A sky130_fd_sc_hd__and2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6963_ _6963_/CLK _6963_/D vssd1 vssd1 vccd1 vccd1 _6963_/Q sky130_fd_sc_hd__dfxtp_1
X_6894_ _6894_/CLK _6894_/D vssd1 vssd1 vccd1 vccd1 _6894_/Q sky130_fd_sc_hd__dfxtp_1
X_5914_ _5918_/A _5913_/A _7090_/Q vssd1 vssd1 vccd1 vccd1 _5915_/C sky130_fd_sc_hd__o21a_1
XFILLER_21_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5776_ _5776_/A _5776_/B vssd1 vssd1 vccd1 vccd1 _6779_/D sky130_fd_sc_hd__nor2_1
XFILLER_22_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4727_ _6768_/Q vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__2525_ _5200_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2525_/X sky130_fd_sc_hd__clkbuf_16
X_4658_ _3865_/X _6471_/Q _4660_/S vssd1 vssd1 vccd1 vccd1 _4659_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2456_ _5030_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2456_/X sky130_fd_sc_hd__clkbuf_16
Xinput90 wbs_data_i[29] vssd1 vssd1 vccd1 vccd1 _7154_/A sky130_fd_sc_hd__buf_4
X_3609_ _6926_/Q _3608_/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3610_/A sky130_fd_sc_hd__mux2_1
X_4589_ _4589_/A vssd1 vssd1 vccd1 vccd1 _6502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6259_ _6267_/A _6259_/B _6262_/B vssd1 vssd1 vccd1 vccd1 _6260_/A sky130_fd_sc_hd__and3_1
XFILLER_76_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3008_ _6084_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3008_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3960_ _3960_/A _3308_/X vssd1 vssd1 vccd1 vccd1 _3983_/A sky130_fd_sc_hd__or2b_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5192__248 _5193__249/A vssd1 vssd1 vccd1 vccd1 _6530_/CLK sky130_fd_sc_hd__inv_2
X_3891_ _3891_/A vssd1 vssd1 vccd1 vccd1 _6798_/D sky130_fd_sc_hd__clkbuf_1
X_5630_ _6999_/Q vssd1 vssd1 vccd1 vccd1 _6216_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5561_ _5573_/A vssd1 vssd1 vccd1 vccd1 _5561_/X sky130_fd_sc_hd__buf_1
X_4512_ _4490_/X _6537_/Q _4512_/S vssd1 vssd1 vccd1 vccd1 _4513_/A sky130_fd_sc_hd__mux2_1
X_5492_ _5492_/A vssd1 vssd1 vccd1 vccd1 _5492_/X sky130_fd_sc_hd__buf_1
XFILLER_117_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4443_ _4443_/A vssd1 vssd1 vccd1 vccd1 _6565_/D sky130_fd_sc_hd__clkbuf_1
X_4374_ _6603_/Q _3773_/A _4378_/S vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__mux2_1
X_7093_ _7093_/CLK _7093_/D vssd1 vssd1 vccd1 vccd1 _7093_/Q sky130_fd_sc_hd__dfxtp_1
X_3325_ _3354_/S vssd1 vssd1 vccd1 vccd1 _3342_/S sky130_fd_sc_hd__clkbuf_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3256_/A vssd1 vssd1 vccd1 vccd1 _7076_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6946_ _6946_/CLK _6946_/D vssd1 vssd1 vccd1 vccd1 _6946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6877_ _6883_/CLK _6877_/D vssd1 vssd1 vccd1 vccd1 _6877_/Q sky130_fd_sc_hd__dfxtp_2
X_5828_ _5846_/A vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__buf_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5466__309 _5466__309/A vssd1 vssd1 vccd1 vccd1 _6599_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2756_ clkbuf_0__2756_/X vssd1 vssd1 vccd1 vccd1 _5821_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4090_ _4090_/A vssd1 vssd1 vccd1 vccd1 _6729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6800_ _6800_/CLK _6800_/D vssd1 vssd1 vccd1 vccd1 _6800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4992_ _4992_/A _4992_/B vssd1 vssd1 vccd1 vccd1 _4993_/A sky130_fd_sc_hd__and2_2
XFILLER_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3943_ _5776_/A _3943_/B vssd1 vssd1 vccd1 vccd1 _3943_/Y sky130_fd_sc_hd__nor2_1
X_6731_ _6731_/CLK _6731_/D vssd1 vssd1 vccd1 vccd1 _6731_/Q sky130_fd_sc_hd__dfxtp_1
X_3874_ _3896_/S vssd1 vssd1 vccd1 vccd1 _3887_/S sky130_fd_sc_hd__clkbuf_2
X_6662_ _6662_/CLK _6662_/D vssd1 vssd1 vccd1 vccd1 _6662_/Q sky130_fd_sc_hd__dfxtp_1
X_5613_ _6170_/A _7082_/Q _5659_/B _6161_/A vssd1 vssd1 vccd1 vccd1 _5888_/C sky130_fd_sc_hd__o31ai_4
X_6593_ _6593_/CLK _6593_/D vssd1 vssd1 vccd1 vccd1 _6593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4426_ _3251_/X _6572_/Q _4432_/S vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__mux2_1
X_7145_ _7145_/A vssd1 vssd1 vccd1 vccd1 _7145_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _4357_/A vssd1 vssd1 vccd1 vccd1 _6611_/D sky130_fd_sc_hd__clkbuf_1
X_3308_ _6772_/Q _6767_/Q vssd1 vssd1 vccd1 vccd1 _3308_/X sky130_fd_sc_hd__or2b_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _6641_/Q _4155_/X _4288_/S vssd1 vssd1 vccd1 vccd1 _4289_/A sky130_fd_sc_hd__mux2_1
X_7076_ _7076_/CLK _7076_/D vssd1 vssd1 vccd1 vccd1 _7076_/Q sky130_fd_sc_hd__dfxtp_1
X_3239_ _5113_/B _4761_/B _4761_/C _4761_/D vssd1 vssd1 vccd1 vccd1 _4752_/B sky130_fd_sc_hd__or4_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5472__313 _5473__314/A vssd1 vssd1 vccd1 vccd1 _6603_/CLK sky130_fd_sc_hd__inv_2
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _6929_/CLK _6929_/D vssd1 vssd1 vccd1 vccd1 _6929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5143__209 _5143__209/A vssd1 vssd1 vccd1 vccd1 _6491_/CLK sky130_fd_sc_hd__inv_2
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2739_ clkbuf_0__2739_/X vssd1 vssd1 vccd1 vccd1 _5522__354/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6130__166 _6133__169/A vssd1 vssd1 vccd1 vccd1 _6974_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3590_ _3590_/A vssd1 vssd1 vccd1 vccd1 _6933_/D sky130_fd_sc_hd__clkbuf_1
X_5260_ _6670_/Q _6662_/Q _6654_/Q _6646_/Q _5257_/X _5259_/X vssd1 vssd1 vccd1 vccd1
+ _5260_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4211_ _6675_/Q _4149_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4142_ _4422_/A _4186_/A vssd1 vssd1 vccd1 vccd1 _4165_/S sky130_fd_sc_hd__nor2_2
XFILLER_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4073_ _4055_/X _4071_/X _4072_/Y vssd1 vssd1 vccd1 vccd1 _6734_/D sky130_fd_sc_hd__o21a_1
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2874_ clkbuf_0__2874_/X vssd1 vssd1 vccd1 vccd1 _5878_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4975_ _4973_/X input4/X _4970_/X _4974_/X vssd1 vssd1 vccd1 vccd1 _4975_/X sky130_fd_sc_hd__a22o_2
X_6714_ _6714_/CLK _6714_/D vssd1 vssd1 vccd1 vccd1 _6714_/Q sky130_fd_sc_hd__dfxtp_1
X_3926_ _6783_/Q _3886_/X _3926_/S vssd1 vssd1 vccd1 vccd1 _3927_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3857_ _6808_/Q _3856_/X _3860_/S vssd1 vssd1 vccd1 vccd1 _3858_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6645_ _6645_/CLK _6645_/D vssd1 vssd1 vccd1 vccd1 _6645_/Q sky130_fd_sc_hd__dfxtp_1
X_3788_ _3788_/A vssd1 vssd1 vccd1 vccd1 _3788_/X sky130_fd_sc_hd__buf_2
X_6576_ _6897_/CLK _6576_/D vssd1 vssd1 vccd1 vccd1 _6576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4409_ _4409_/A vssd1 vssd1 vccd1 vccd1 _6588_/D sky130_fd_sc_hd__clkbuf_1
X_5389_ _6675_/Q _6667_/Q _6659_/Q _6651_/Q _5263_/X _5259_/X vssd1 vssd1 vccd1 vccd1
+ _5389_/X sky130_fd_sc_hd__mux4_2
X_7128_ _7128_/A vssd1 vssd1 vccd1 vccd1 _7128_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2524_ clkbuf_0__2524_/X vssd1 vssd1 vccd1 vccd1 _5196__251/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7059_ _7059_/CLK _7059_/D vssd1 vssd1 vccd1 vccd1 _7059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2455_ clkbuf_0__2455_/X vssd1 vssd1 vccd1 vccd1 _6376__4/A sky130_fd_sc_hd__clkbuf_4
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6025__82 _6027__84/A vssd1 vssd1 vccd1 vccd1 _6889_/CLK sky130_fd_sc_hd__inv_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__3007_ clkbuf_0__3007_/X vssd1 vssd1 vccd1 vccd1 _6082__128/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5479__319 _5479__319/A vssd1 vssd1 vccd1 vccd1 _6609_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4760_ _5648_/A vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_119_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3711_ _3680_/X _6867_/Q _3719_/S vssd1 vssd1 vccd1 vccd1 _3712_/A sky130_fd_sc_hd__mux2_1
X_4691_ _5018_/A vssd1 vssd1 vccd1 vccd1 _4691_/X sky130_fd_sc_hd__clkbuf_2
X_3642_ _3708_/A _4167_/A _4167_/B vssd1 vssd1 vccd1 vccd1 _4608_/B sky130_fd_sc_hd__or3_1
X_6430_ _6430_/A _6430_/B vssd1 vssd1 vccd1 vccd1 _6431_/A sky130_fd_sc_hd__or2_2
X_6361_ _6367_/A vssd1 vssd1 vccd1 vccd1 _6361_/X sky130_fd_sc_hd__buf_1
X_3573_ _3384_/X _6940_/Q _3577_/S vssd1 vssd1 vccd1 vccd1 _3574_/A sky130_fd_sc_hd__mux2_1
X_5312_ _5329_/A vssd1 vssd1 vccd1 vccd1 _5312_/X sky130_fd_sc_hd__clkbuf_4
X_6292_ _7018_/Q _6292_/B vssd1 vssd1 vccd1 vccd1 _6292_/X sky130_fd_sc_hd__or2_1
XFILLER_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4125_ _6713_/Q _3871_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4126_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4056_ _6733_/Q vssd1 vssd1 vccd1 vccd1 _5334_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_45_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2857_ clkbuf_0__2857_/X vssd1 vssd1 vccd1 vccd1 _5777__474/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _4774_/X _4957_/X _4865_/A vssd1 vssd1 vccd1 vccd1 _4958_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4889_ _7091_/Q vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__2756_ _5597_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2756_/X sky130_fd_sc_hd__clkbuf_16
X_3909_ _3909_/A vssd1 vssd1 vccd1 vccd1 _6791_/D sky130_fd_sc_hd__clkbuf_1
X_6628_ _6628_/CLK _6628_/D vssd1 vssd1 vccd1 vccd1 _6628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6559_ _6559_/CLK _6559_/D vssd1 vssd1 vccd1 vccd1 _6559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5930_ _5966_/A vssd1 vssd1 vccd1 vccd1 _5954_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5156__219 _5156__219/A vssd1 vssd1 vccd1 vccd1 _6501_/CLK sky130_fd_sc_hd__inv_2
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4812_ _4806_/X _4807_/X _4811_/X vssd1 vssd1 vccd1 vccd1 _4812_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4743_ _5044_/C vssd1 vssd1 vccd1 vccd1 _4748_/B sky130_fd_sc_hd__inv_2
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4674_ _3862_/X _6438_/Q _4678_/S vssd1 vssd1 vccd1 vccd1 _4675_/A sky130_fd_sc_hd__mux2_1
X_6413_ _6425_/A _6413_/B vssd1 vssd1 vccd1 vccd1 _6414_/A sky130_fd_sc_hd__and2_1
X_3625_ _3357_/X _6921_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _3626_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3556_ _3556_/A vssd1 vssd1 vccd1 vccd1 _6948_/D sky130_fd_sc_hd__clkbuf_1
X_6275_ _7012_/Q _6292_/B _6247_/A vssd1 vssd1 vccd1 vccd1 _6276_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3487_ _4626_/A _4608_/A vssd1 vssd1 vccd1 vccd1 _3503_/S sky130_fd_sc_hd__or2_2
X_5157_ _5163_/A vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__buf_1
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4108_ _4108_/A vssd1 vssd1 vccd1 vccd1 _6721_/D sky130_fd_sc_hd__clkbuf_1
X_5088_ _5088_/A vssd1 vssd1 vccd1 vccd1 _6460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4039_ _4044_/B vssd1 vssd1 vccd1 vccd1 _4049_/B sky130_fd_sc_hd__inv_2
XFILLER_71_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2739_ _5517_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2739_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5549__375 _5550__376/A vssd1 vssd1 vccd1 vccd1 _6665_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5040__187 _5040__187/A vssd1 vssd1 vccd1 vccd1 _6443_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3410_ _3341_/X _7042_/Q _3410_/S vssd1 vssd1 vccd1 vccd1 _3411_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4390_ _3251_/X _6596_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4391_/A sky130_fd_sc_hd__mux2_1
X_3341_ _4023_/A vssd1 vssd1 vccd1 vccd1 _3341_/X sky130_fd_sc_hd__buf_2
XFILLER_112_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6060_ _6078_/A vssd1 vssd1 vccd1 vccd1 _6060_/X sky130_fd_sc_hd__buf_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _6739_/Q _6737_/Q _4204_/A vssd1 vssd1 vccd1 vccd1 _3579_/A sky130_fd_sc_hd__or3b_4
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5011_ _5011_/A vssd1 vssd1 vccd1 vccd1 _5011_/X sky130_fd_sc_hd__clkbuf_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6962_ _6962_/CLK _6962_/D vssd1 vssd1 vccd1 vccd1 _6962_/Q sky130_fd_sc_hd__dfxtp_1
X_6893_ _6893_/CLK _6893_/D vssd1 vssd1 vccd1 vccd1 _6893_/Q sky130_fd_sc_hd__dfxtp_1
X_5913_ _5913_/A _5913_/B vssd1 vssd1 vccd1 vccd1 _5915_/B sky130_fd_sc_hd__nor2_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5775_ _5775_/A vssd1 vssd1 vccd1 vccd1 _6778_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4726_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4726_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__2524_ _5194_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2524_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4657_ _4657_/A vssd1 vssd1 vccd1 vccd1 _6472_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__2455_ _5029_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2455_/X sky130_fd_sc_hd__clkbuf_16
X_3608_ _7027_/Q vssd1 vssd1 vccd1 vccd1 _3608_/X sky130_fd_sc_hd__clkbuf_8
Xinput91 wbs_data_i[2] vssd1 vssd1 vccd1 vccd1 _7127_/A sky130_fd_sc_hd__buf_8
Xinput80 wbs_data_i[1] vssd1 vssd1 vccd1 vccd1 _7126_/A sky130_fd_sc_hd__buf_8
X_4588_ _4499_/X _6502_/Q _4588_/S vssd1 vssd1 vccd1 vccd1 _4589_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3539_ _3539_/A vssd1 vssd1 vccd1 vccd1 _6955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6258_ _7008_/Q _6258_/B vssd1 vssd1 vccd1 vccd1 _6262_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6189_ _6189_/A vssd1 vssd1 vccd1 vccd1 _6994_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__3007_ _6078_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3007_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5226__275 _5230__279/A vssd1 vssd1 vccd1 vccd1 _6557_/CLK sky130_fd_sc_hd__inv_2
X_3890_ _6798_/Q _3889_/X _3896_/S vssd1 vssd1 vccd1 vccd1 _3891_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5560_ _5560_/A vssd1 vssd1 vccd1 vccd1 _5560_/X sky130_fd_sc_hd__buf_1
XFILLER_31_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4511_ _4511_/A vssd1 vssd1 vccd1 vccd1 _6538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4442_ _4009_/X _6565_/Q _4450_/S vssd1 vssd1 vccd1 vccd1 _4443_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7161_ _7161_/A vssd1 vssd1 vccd1 vccd1 _7161_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4373_ _4373_/A vssd1 vssd1 vccd1 vccd1 _6604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3324_ _4644_/A _4662_/A vssd1 vssd1 vccd1 vccd1 _3354_/S sky130_fd_sc_hd__or2_2
X_7092_ _7095_/CLK _7092_/D vssd1 vssd1 vccd1 vccd1 _7092_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _7076_/Q _3254_/X _3261_/S vssd1 vssd1 vccd1 vccd1 _3256_/A sky130_fd_sc_hd__mux2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5127__195 _5131__199/A vssd1 vssd1 vccd1 vccd1 _6477_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _6945_/CLK _6945_/D vssd1 vssd1 vccd1 vccd1 _6945_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_6876_ _7008_/CLK _6876_/D vssd1 vssd1 vccd1 vccd1 _6876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4709_ _4719_/A vssd1 vssd1 vccd1 vccd1 _4709_/X sky130_fd_sc_hd__buf_4
XFILLER_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2755_ clkbuf_0__2755_/X vssd1 vssd1 vccd1 vccd1 _5594__407/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _4991_/A vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__clkbuf_1
X_6730_ _6730_/CLK _6730_/D vssd1 vssd1 vccd1 vccd1 _6730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _3990_/B _3943_/B _3937_/Y vssd1 vssd1 vccd1 vccd1 _6775_/D sky130_fd_sc_hd__o21a_1
X_3873_ _4168_/A _3873_/B vssd1 vssd1 vccd1 vccd1 _3896_/S sky130_fd_sc_hd__nor2_2
X_6661_ _6661_/CLK _6661_/D vssd1 vssd1 vccd1 vccd1 _6661_/Q sky130_fd_sc_hd__dfxtp_1
X_5612_ _7010_/Q vssd1 vssd1 vccd1 vccd1 _6266_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6592_ _6592_/CLK _6592_/D vssd1 vssd1 vccd1 vccd1 _6592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5474_ _5492_/A vssd1 vssd1 vccd1 vccd1 _5474_/X sky130_fd_sc_hd__buf_1
X_4425_ _4425_/A vssd1 vssd1 vccd1 vccd1 _6573_/D sky130_fd_sc_hd__clkbuf_1
X_7144_ _7144_/A vssd1 vssd1 vccd1 vccd1 _7144_/X sky130_fd_sc_hd__clkbuf_1
X_4356_ _6611_/Q _3773_/A _4360_/S vssd1 vssd1 vccd1 vccd1 _4357_/A sky130_fd_sc_hd__mux2_1
X_5506__340 _5510__344/A vssd1 vssd1 vccd1 vccd1 _6630_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3307_ _3941_/B _3961_/A vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__xnor2_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5875__72 _5876__73/A vssd1 vssd1 vccd1 vccd1 _6858_/CLK sky130_fd_sc_hd__inv_2
X_4287_ _4287_/A vssd1 vssd1 vccd1 vccd1 _6642_/D sky130_fd_sc_hd__clkbuf_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7075_ _7075_/CLK _7075_/D vssd1 vssd1 vccd1 vccd1 _7075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3238_ _6456_/Q _6457_/Q _6458_/Q _6455_/Q vssd1 vssd1 vccd1 vccd1 _4761_/D sky130_fd_sc_hd__or4b_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6037__91 _6038__92/A vssd1 vssd1 vccd1 vccd1 _6899_/CLK sky130_fd_sc_hd__inv_2
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6928_ _6928_/CLK _6928_/D vssd1 vssd1 vccd1 vccd1 _6928_/Q sky130_fd_sc_hd__dfxtp_1
X_6859_ _6859_/CLK _6859_/D vssd1 vssd1 vccd1 vccd1 _6859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2738_ clkbuf_0__2738_/X vssd1 vssd1 vccd1 vccd1 _5514__347/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6098__140 _6099__141/A vssd1 vssd1 vccd1 vccd1 _6948_/CLK sky130_fd_sc_hd__inv_2
X_4210_ _4210_/A vssd1 vssd1 vccd1 vccd1 _6676_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4141_ _7030_/Q vssd1 vssd1 vccd1 vccd1 _4141_/X sky130_fd_sc_hd__buf_4
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4072_ _4055_/X _4071_/X _6303_/B vssd1 vssd1 vccd1 vccd1 _4072_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2873_ clkbuf_0__2873_/X vssd1 vssd1 vccd1 vccd1 _6115_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4974_ _7086_/Q vssd1 vssd1 vccd1 vccd1 _4974_/X sky130_fd_sc_hd__clkbuf_4
X_6713_ _6713_/CLK _6713_/D vssd1 vssd1 vccd1 vccd1 _6713_/Q sky130_fd_sc_hd__dfxtp_1
X_3925_ _3925_/A vssd1 vssd1 vccd1 vccd1 _6784_/D sky130_fd_sc_hd__clkbuf_1
X_6644_ _6644_/CLK _6644_/D vssd1 vssd1 vccd1 vccd1 _6644_/Q sky130_fd_sc_hd__dfxtp_1
X_3856_ _6745_/Q vssd1 vssd1 vccd1 vccd1 _3856_/X sky130_fd_sc_hd__buf_6
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3787_ _3787_/A vssd1 vssd1 vccd1 vccd1 _6837_/D sky130_fd_sc_hd__clkbuf_1
X_6575_ _6897_/CLK _6575_/D vssd1 vssd1 vccd1 vccd1 _6575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4408_ _3251_/X _6588_/Q _4414_/S vssd1 vssd1 vccd1 vccd1 _4409_/A sky130_fd_sc_hd__mux2_1
X_5388_ _7076_/Q _6702_/Q _6571_/Q _6849_/Q _5251_/X _5254_/X vssd1 vssd1 vccd1 vccd1
+ _5388_/X sky130_fd_sc_hd__mux4_1
X_7127_ _7127_/A vssd1 vssd1 vccd1 vccd1 _7127_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4339_ _4339_/A vssd1 vssd1 vccd1 vccd1 _6619_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2523_ clkbuf_0__2523_/X vssd1 vssd1 vccd1 vccd1 _5193__249/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7058_ _7058_/CLK _7058_/D vssd1 vssd1 vccd1 vccd1 _7058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6009_ _5936_/X _6012_/B _6012_/D vssd1 vssd1 vccd1 vccd1 _6009_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3006_ clkbuf_0__3006_/X vssd1 vssd1 vccd1 vccd1 _6075__122/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5706__436 _5709__439/A vssd1 vssd1 vccd1 vccd1 _6730_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5752__456 _5752__456/A vssd1 vssd1 vccd1 vccd1 _6760_/CLK sky130_fd_sc_hd__inv_2
XFILLER_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3725_/S vssd1 vssd1 vccd1 vccd1 _3719_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4690_ _5005_/A vssd1 vssd1 vccd1 vccd1 _5018_/A sky130_fd_sc_hd__buf_4
X_3641_ _4662_/A vssd1 vssd1 vccd1 vccd1 _4458_/A sky130_fd_sc_hd__buf_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3572_ _3572_/A vssd1 vssd1 vccd1 vccd1 _6941_/D sky130_fd_sc_hd__clkbuf_1
X_5311_ _5337_/A vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__clkbuf_8
X_6291_ _7018_/Q _6284_/X _6289_/X _6290_/X vssd1 vssd1 vccd1 vccd1 _7017_/D sky130_fd_sc_hd__o211a_1
XFILLER_102_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4124_ _4139_/S vssd1 vssd1 vccd1 vccd1 _4133_/S sky130_fd_sc_hd__buf_2
XFILLER_56_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput1 caravel_uart_rx vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4055_ _5324_/A vssd1 vssd1 vccd1 vccd1 _4055_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0__2856_ clkbuf_0__2856_/X vssd1 vssd1 vccd1 vccd1 _5766__467/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4957_ _6896_/Q _6525_/Q _4957_/S vssd1 vssd1 vccd1 vccd1 _4957_/X sky130_fd_sc_hd__mux2_1
X_4888_ _5018_/A vssd1 vssd1 vccd1 vccd1 _4888_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__2755_ _5591_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2755_/X sky130_fd_sc_hd__clkbuf_16
X_3908_ _6791_/Q _3611_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3909_/A sky130_fd_sc_hd__mux2_1
X_6627_ _6627_/CLK _6627_/D vssd1 vssd1 vccd1 vccd1 _6627_/Q sky130_fd_sc_hd__dfxtp_1
X_3839_ _6814_/Q _3614_/X _3843_/S vssd1 vssd1 vccd1 vccd1 _3840_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6558_ _6558_/CLK _6558_/D vssd1 vssd1 vccd1 vccd1 _6558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6489_ _6489_/CLK _6489_/D vssd1 vssd1 vccd1 vccd1 _6489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6049__101 _6049__101/A vssd1 vssd1 vccd1 vccd1 _6909_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5485__324 _5485__324/A vssd1 vssd1 vccd1 vccd1 _6614_/CLK sky130_fd_sc_hd__inv_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5860_ _5866_/A vssd1 vssd1 vccd1 vccd1 _5860_/X sky130_fd_sc_hd__buf_1
XFILLER_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4808_/X _4810_/X _4865_/A vssd1 vssd1 vccd1 vccd1 _4811_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5791_ _5815_/A vssd1 vssd1 vccd1 vccd1 _5791_/X sky130_fd_sc_hd__buf_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4742_ _6447_/Q _5736_/B _4794_/B vssd1 vssd1 vccd1 vccd1 _5044_/C sky130_fd_sc_hd__and3_1
XFILLER_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _4673_/A vssd1 vssd1 vccd1 vccd1 _6439_/D sky130_fd_sc_hd__clkbuf_1
X_6143__177 _6143__177/A vssd1 vssd1 vccd1 vccd1 _6985_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6412_ _7132_/A _6167_/A _6424_/S vssd1 vssd1 vccd1 vccd1 _6413_/B sky130_fd_sc_hd__mux2_1
X_3624_ _3639_/S vssd1 vssd1 vccd1 vccd1 _3633_/S sky130_fd_sc_hd__clkbuf_2
X_6343_ _6367_/A vssd1 vssd1 vccd1 vccd1 _6343_/X sky130_fd_sc_hd__buf_1
X_3555_ _6948_/Q _3456_/X _3559_/S vssd1 vssd1 vccd1 vccd1 _3556_/A sky130_fd_sc_hd__mux2_1
X_6322__13 _6323__14/A vssd1 vssd1 vccd1 vccd1 _7033_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6274_ _6282_/A vssd1 vssd1 vccd1 vccd1 _6292_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3486_ _3947_/A _3946_/B vssd1 vssd1 vccd1 vccd1 _4608_/A sky130_fd_sc_hd__nand2_4
X_5225_ _5231_/A vssd1 vssd1 vccd1 vccd1 _5225_/X sky130_fd_sc_hd__buf_1
XFILLER_103_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4107_ _6721_/Q _3871_/X _4115_/S vssd1 vssd1 vccd1 vccd1 _4108_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5087_ _6460_/Q _7114_/A _5093_/S vssd1 vssd1 vccd1 vccd1 _5088_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4038_ _6740_/Q _6749_/Q _4035_/Y _4037_/X vssd1 vssd1 vccd1 vccd1 _6740_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1_0__2839_ clkbuf_0__2839_/X vssd1 vssd1 vccd1 vccd1 _5743__449/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5989_ _5989_/A vssd1 vssd1 vccd1 vccd1 _6879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2738_ _5511_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2738_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput190 _5000_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[22] sky130_fd_sc_hd__buf_2
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3340_ _6744_/Q vssd1 vssd1 vccd1 vccd1 _4023_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5014_/A _5010_/B vssd1 vssd1 vccd1 vccd1 _5011_/A sky130_fd_sc_hd__and2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3271_/A vssd1 vssd1 vccd1 vccd1 _7071_/D sky130_fd_sc_hd__clkbuf_1
X_5162__224 _5162__224/A vssd1 vssd1 vccd1 vccd1 _6506_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5500__335 _5502__337/A vssd1 vssd1 vccd1 vccd1 _6625_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6961_ _6961_/CLK _6961_/D vssd1 vssd1 vccd1 vccd1 _6961_/Q sky130_fd_sc_hd__dfxtp_1
X_6892_ _6892_/CLK _6892_/D vssd1 vssd1 vccd1 vccd1 _6892_/Q sky130_fd_sc_hd__dfxtp_1
X_5912_ _5912_/A _5912_/B _5912_/C _5911_/X vssd1 vssd1 vccd1 vccd1 _5921_/C sky130_fd_sc_hd__or4b_1
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5774_ _7079_/Q _6705_/Q _5774_/C vssd1 vssd1 vccd1 vccd1 _5775_/A sky130_fd_sc_hd__and3_1
X_4725_ _4703_/Y _4712_/Y _4716_/Y _4723_/Y _4904_/A vssd1 vssd1 vccd1 vccd1 _4725_/X
+ sky130_fd_sc_hd__o221a_1
X_5765__466 _5766__467/A vssd1 vssd1 vccd1 vccd1 _6770_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__2523_ _5188_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2523_/X sky130_fd_sc_hd__clkbuf_16
X_4656_ _3862_/X _6472_/Q _4660_/S vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__mux2_1
X_4587_ _4587_/A vssd1 vssd1 vccd1 vccd1 _6503_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__2454_ _5028_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2454_/X sky130_fd_sc_hd__clkbuf_16
Xinput70 wbs_data_i[10] vssd1 vssd1 vccd1 vccd1 _7135_/A sky130_fd_sc_hd__buf_4
Xinput81 wbs_data_i[20] vssd1 vssd1 vccd1 vccd1 _7145_/A sky130_fd_sc_hd__buf_4
X_3607_ _3607_/A vssd1 vssd1 vccd1 vccd1 _6927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput92 wbs_data_i[30] vssd1 vssd1 vccd1 vccd1 _7155_/A sky130_fd_sc_hd__buf_4
X_3538_ _6955_/Q _3459_/X _3540_/S vssd1 vssd1 vccd1 vccd1 _3539_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6257_ _7008_/Q _6258_/B vssd1 vssd1 vccd1 vccd1 _6259_/B sky130_fd_sc_hd__or2_1
X_3469_ _3469_/A vssd1 vssd1 vccd1 vccd1 _6985_/D sky130_fd_sc_hd__clkbuf_1
X_6188_ _6290_/A _6188_/B _6188_/C vssd1 vssd1 vccd1 vccd1 _6189_/A sky130_fd_sc_hd__and3_1
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__3006_ _6072_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3006_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5555__380 _5559__384/A vssd1 vssd1 vccd1 vccd1 _6670_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6092__135 _6094__137/A vssd1 vssd1 vccd1 vccd1 _6943_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4510_ _4487_/X _6538_/Q _4512_/S vssd1 vssd1 vccd1 vccd1 _4511_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4441_ _4456_/S vssd1 vssd1 vccd1 vccd1 _4450_/S sky130_fd_sc_hd__buf_2
XFILLER_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7160_ _7160_/A vssd1 vssd1 vccd1 vccd1 _7160_/X sky130_fd_sc_hd__buf_4
X_4372_ _6604_/Q _3770_/A _4378_/S vssd1 vssd1 vccd1 vccd1 _4373_/A sky130_fd_sc_hd__mux2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5887__81 _5887__81/A vssd1 vssd1 vccd1 vccd1 _6867_/CLK sky130_fd_sc_hd__inv_2
X_7091_ _7093_/CLK _7091_/D vssd1 vssd1 vccd1 vccd1 _7091_/Q sky130_fd_sc_hd__dfxtp_1
X_3323_ _3661_/A _3949_/A _3936_/A vssd1 vssd1 vccd1 vccd1 _4662_/A sky130_fd_sc_hd__or3_4
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3254_ _7028_/Q vssd1 vssd1 vccd1 vccd1 _3254_/X sky130_fd_sc_hd__clkbuf_4
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6944_ _6944_/CLK _6944_/D vssd1 vssd1 vccd1 vccd1 _6944_/Q sky130_fd_sc_hd__dfxtp_1
X_6875_ _7008_/CLK _6875_/D vssd1 vssd1 vccd1 vccd1 _6875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5847__530 _5849__532/A vssd1 vssd1 vccd1 vccd1 _6836_/CLK sky130_fd_sc_hd__inv_2
X_5757_ _5778_/A vssd1 vssd1 vccd1 vccd1 _5757_/X sky130_fd_sc_hd__buf_1
X_4708_ _6768_/Q vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4639_ _4639_/A vssd1 vssd1 vccd1 vccd1 _6480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6309_ _6309_/A vssd1 vssd1 vccd1 vccd1 _7025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5232__280 _5235__283/A vssd1 vssd1 vccd1 vccd1 _6562_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6100__142 _6102__144/A vssd1 vssd1 vccd1 vccd1 _6950_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _4992_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4991_/A sky130_fd_sc_hd__and2_2
X_3941_ _6778_/Q _3941_/B _4765_/A vssd1 vssd1 vccd1 vccd1 _3943_/B sky130_fd_sc_hd__and3_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3872_ _4608_/A vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__clkbuf_4
X_6660_ _6660_/CLK _6660_/D vssd1 vssd1 vccd1 vccd1 _6660_/Q sky130_fd_sc_hd__dfxtp_1
X_5611_ _7011_/Q vssd1 vssd1 vccd1 vccd1 _6269_/A sky130_fd_sc_hd__inv_2
X_6591_ _6591_/CLK _6591_/D vssd1 vssd1 vccd1 vccd1 _6591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5542_ _5548_/A vssd1 vssd1 vccd1 vccd1 _5542_/X sky130_fd_sc_hd__buf_1
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4424_ _3200_/X _6573_/Q _4432_/S vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__mux2_1
X_7143_ _7143_/A vssd1 vssd1 vccd1 vccd1 _7143_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4355_ _4355_/A vssd1 vssd1 vccd1 vccd1 _6612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3306_ _6775_/Q _6770_/Q vssd1 vssd1 vccd1 vccd1 _3961_/A sky130_fd_sc_hd__xnor2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7074_ _7074_/CLK _7074_/D vssd1 vssd1 vccd1 vccd1 _7074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4286_ _6642_/Q _4152_/X _4288_/S vssd1 vssd1 vccd1 vccd1 _4287_/A sky130_fd_sc_hd__mux2_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3237_ _6463_/Q _6464_/Q _6465_/Q _6466_/Q vssd1 vssd1 vccd1 vccd1 _4761_/C sky130_fd_sc_hd__or4_4
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6927_ _6927_/CLK _6927_/D vssd1 vssd1 vccd1 vccd1 _6927_/Q sky130_fd_sc_hd__dfxtp_1
X_6858_ _6858_/CLK _6858_/D vssd1 vssd1 vccd1 vccd1 _6858_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3022_ clkbuf_0__3022_/X vssd1 vssd1 vccd1 vccd1 _6323__14/A sky130_fd_sc_hd__clkbuf_4
X_5809_ _5809_/A vssd1 vssd1 vccd1 vccd1 _5809_/X sky130_fd_sc_hd__buf_1
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6789_ _6789_/CLK _6789_/D vssd1 vssd1 vccd1 vccd1 _6789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2737_ clkbuf_0__2737_/X vssd1 vssd1 vccd1 vccd1 _5510__344/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_50 _7055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5568__390 _5569__391/A vssd1 vssd1 vccd1 vccd1 _6680_/CLK sky130_fd_sc_hd__inv_2
X_4140_ _4140_/A vssd1 vssd1 vccd1 vccd1 _6706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4071_ _4071_/A _4071_/B _4081_/A vssd1 vssd1 vccd1 vccd1 _4071_/X sky130_fd_sc_hd__and3_1
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2872_ clkbuf_0__2872_/X vssd1 vssd1 vccd1 vccd1 _5849__532/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4973_ _5018_/A vssd1 vssd1 vccd1 vccd1 _4973_/X sky130_fd_sc_hd__clkbuf_2
X_6712_ _6712_/CLK _6712_/D vssd1 vssd1 vccd1 vccd1 _6712_/Q sky130_fd_sc_hd__dfxtp_1
X_3924_ _6784_/Q _3883_/X _3926_/S vssd1 vssd1 vccd1 vccd1 _3925_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6329__19 _6329__19/A vssd1 vssd1 vccd1 vccd1 _7039_/CLK sky130_fd_sc_hd__inv_2
X_6643_ _6643_/CLK _6643_/D vssd1 vssd1 vccd1 vccd1 _6643_/Q sky130_fd_sc_hd__dfxtp_1
X_6107__148 _6108__149/A vssd1 vssd1 vccd1 vccd1 _6956_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3855_ _3855_/A vssd1 vssd1 vccd1 vccd1 _6809_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6574_ _6897_/CLK _6574_/D vssd1 vssd1 vccd1 vccd1 _6574_/Q sky130_fd_sc_hd__dfxtp_1
X_3786_ _3785_/X _6837_/Q _3789_/S vssd1 vssd1 vccd1 vccd1 _3787_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4407_ _4407_/A vssd1 vssd1 vccd1 vccd1 _6589_/D sky130_fd_sc_hd__clkbuf_1
X_5387_ _6578_/Q _5250_/X _5386_/X _5298_/X vssd1 vssd1 vccd1 vccd1 _6578_/D sky130_fd_sc_hd__o211a_1
X_7126_ _7126_/A vssd1 vssd1 vccd1 vccd1 _7126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4338_ _3773_/X _6619_/Q _4342_/S vssd1 vssd1 vccd1 vccd1 _4339_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__2522_ clkbuf_0__2522_/X vssd1 vssd1 vccd1 vccd1 _5187__244/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7057_ _7057_/CLK _7057_/D vssd1 vssd1 vccd1 vccd1 _7057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4269_ _6649_/Q _4155_/X _4269_/S vssd1 vssd1 vccd1 vccd1 _4270_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__2453_ clkbuf_0__2453_/X vssd1 vssd1 vccd1 vccd1 _6342_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6008_ _6008_/A vssd1 vssd1 vccd1 vccd1 _6883_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3005_ clkbuf_0__3005_/X vssd1 vssd1 vccd1 vccd1 _6071__119/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2735_ clkbuf_0__2735_/X vssd1 vssd1 vccd1 vccd1 _5499_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6031__87 _6033__89/A vssd1 vssd1 vccd1 vccd1 _6894_/CLK sky130_fd_sc_hd__inv_2
X_3640_ _3640_/A vssd1 vssd1 vccd1 vccd1 _6914_/D sky130_fd_sc_hd__clkbuf_1
X_3571_ _3380_/X _6941_/Q _3571_/S vssd1 vssd1 vccd1 vccd1 _3572_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6290_ _6290_/A vssd1 vssd1 vccd1 vccd1 _6290_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5310_ _4071_/A _5301_/X _5305_/Y _5307_/X _5309_/Y vssd1 vssd1 vccd1 vccd1 _5310_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4123_ _4168_/A _4123_/B vssd1 vssd1 vccd1 vccd1 _4139_/S sky130_fd_sc_hd__nor2_2
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput2 caravel_wb_ack_i vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
XFILLER_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4054_ _6734_/Q vssd1 vssd1 vccd1 vccd1 _5324_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__2855_ clkbuf_0__2855_/X vssd1 vssd1 vccd1 vccd1 _5760__462/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4956_ _6501_/Q _6517_/Q _4956_/S vssd1 vssd1 vccd1 vccd1 _4956_/X sky130_fd_sc_hd__mux2_1
X_4887_ _4691_/X input29/X _4695_/X _4886_/X vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__a22o_2
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3907_ _3907_/A vssd1 vssd1 vccd1 vccd1 _6792_/D sky130_fd_sc_hd__clkbuf_1
X_6626_ _6626_/CLK _6626_/D vssd1 vssd1 vccd1 vccd1 _6626_/Q sky130_fd_sc_hd__dfxtp_1
X_3838_ _3838_/A vssd1 vssd1 vccd1 vccd1 _6815_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6557_ _6557_/CLK _6557_/D vssd1 vssd1 vccd1 vccd1 _6557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3769_ _3769_/A vssd1 vssd1 vccd1 vccd1 _6843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6488_ _6488_/CLK _6488_/D vssd1 vssd1 vccd1 vccd1 _6488_/Q sky130_fd_sc_hd__dfxtp_1
X_5439_ _5438_/X _5439_/B vssd1 vssd1 vccd1 vccd1 _5439_/X sky130_fd_sc_hd__and2b_1
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7109_ _7109_/A vssd1 vssd1 vccd1 vccd1 _7109_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6750_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_5519__351 _5519__351/A vssd1 vssd1 vccd1 vccd1 _6641_/CLK sky130_fd_sc_hd__inv_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5712__441 _5713__442/A vssd1 vssd1 vccd1 vccd1 _6735_/CLK sky130_fd_sc_hd__inv_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5450__295 _5454__299/A vssd1 vssd1 vccd1 vccd1 _6585_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6056__106 _6059__109/A vssd1 vssd1 vccd1 vccd1 _6914_/CLK sky130_fd_sc_hd__inv_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _6480_/Q _6552_/Q _4957_/S vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5790_ _5821_/A vssd1 vssd1 vccd1 vccd1 _5790_/X sky130_fd_sc_hd__buf_1
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _6448_/Q _4741_/B vssd1 vssd1 vccd1 vccd1 _4794_/B sky130_fd_sc_hd__nor2_1
X_4672_ _3859_/X _6439_/Q _4672_/S vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__mux2_1
X_6411_ _6432_/S vssd1 vssd1 vccd1 vccd1 _6424_/S sky130_fd_sc_hd__clkbuf_2
X_3623_ _3623_/A _3623_/B _4296_/A vssd1 vssd1 vccd1 vccd1 _3639_/S sky130_fd_sc_hd__or3_4
X_5841__525 _5843__527/A vssd1 vssd1 vccd1 vccd1 _6831_/CLK sky130_fd_sc_hd__inv_2
X_6342_ _6342_/A vssd1 vssd1 vccd1 vccd1 _6342_/X sky130_fd_sc_hd__buf_1
X_3554_ _3554_/A vssd1 vssd1 vccd1 vccd1 _6949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6273_ _6271_/X _6280_/B _7012_/Q vssd1 vssd1 vccd1 vccd1 _6276_/A sky130_fd_sc_hd__and3b_1
X_3485_ _3485_/A _3485_/B vssd1 vssd1 vccd1 vccd1 _3946_/B sky130_fd_sc_hd__nor2_2
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3022_ _6153_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3022_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4106_ _4121_/S vssd1 vssd1 vccd1 vccd1 _4115_/S sky130_fd_sc_hd__buf_2
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5086_ _5086_/A vssd1 vssd1 vccd1 vccd1 _6459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4037_ _6305_/A vssd1 vssd1 vccd1 vccd1 _4037_/X sky130_fd_sc_hd__buf_2
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__2838_ clkbuf_0__2838_/X vssd1 vssd1 vccd1 vccd1 _5713__442/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5988_ _6002_/A _5988_/B vssd1 vssd1 vccd1 vccd1 _5989_/A sky130_fd_sc_hd__and2_1
X_4939_ _4935_/X _4937_/X _4938_/X _3968_/A _3974_/A vssd1 vssd1 vccd1 vccd1 _4939_/X
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__2737_ _5505_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2737_/X sky130_fd_sc_hd__clkbuf_16
X_6609_ _6609_/CLK _6609_/D vssd1 vssd1 vccd1 vccd1 _6609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput191 _5002_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput180 _4981_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[13] sky130_fd_sc_hd__buf_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _7071_/Q _3269_/X _3270_/S vssd1 vssd1 vccd1 vccd1 _3271_/A sky130_fd_sc_hd__mux2_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6960_ _6960_/CLK _6960_/D vssd1 vssd1 vccd1 vccd1 _6960_/Q sky130_fd_sc_hd__dfxtp_1
X_5911_ _4760_/X _6870_/Q _5911_/S vssd1 vssd1 vccd1 vccd1 _5911_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6891_ _6891_/CLK _6891_/D vssd1 vssd1 vccd1 vccd1 _6891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4724_ _4724_/A vssd1 vssd1 vccd1 vccd1 _4904_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__2522_ _5182_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2522_/X sky130_fd_sc_hd__clkbuf_16
X_4655_ _4655_/A vssd1 vssd1 vccd1 vccd1 _6473_/D sky130_fd_sc_hd__clkbuf_1
X_4586_ _4496_/X _6503_/Q _4588_/S vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__2453_ _5027_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2453_/X sky130_fd_sc_hd__clkbuf_16
Xinput60 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 _4682_/A sky130_fd_sc_hd__clkbuf_1
Xinput82 wbs_data_i[21] vssd1 vssd1 vccd1 vccd1 _7146_/A sky130_fd_sc_hd__buf_4
Xinput71 wbs_data_i[11] vssd1 vssd1 vccd1 vccd1 _7136_/A sky130_fd_sc_hd__buf_4
X_3606_ _6927_/Q _3605_/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__mux2_1
X_5806__497 _5806__497/A vssd1 vssd1 vccd1 vccd1 _6803_/CLK sky130_fd_sc_hd__inv_2
Xinput93 wbs_data_i[31] vssd1 vssd1 vccd1 vccd1 _7156_/A sky130_fd_sc_hd__buf_4
X_3537_ _3537_/A vssd1 vssd1 vccd1 vccd1 _6956_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6256_ _7007_/Q _6249_/X _6255_/Y _6238_/A vssd1 vssd1 vccd1 vccd1 _7007_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3468_ _3357_/X _6985_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3469_/A sky130_fd_sc_hd__mux2_1
X_5207_ _5213_/A vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__buf_1
X_6187_ _6245_/B _6187_/B _6187_/C vssd1 vssd1 vccd1 vccd1 _6188_/C sky130_fd_sc_hd__or3_1
X_3399_ _3708_/A _4167_/A _4167_/B vssd1 vssd1 vccd1 vccd1 _4626_/A sky130_fd_sc_hd__or3b_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5138_ _5138_/A vssd1 vssd1 vccd1 vccd1 _5138_/X sky130_fd_sc_hd__buf_1
Xclkbuf_0__3005_ _6066_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3005_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5069_ _6452_/Q _7106_/A _5071_/S vssd1 vssd1 vccd1 vccd1 _5070_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5139__205 _5140__206/A vssd1 vssd1 vccd1 vccd1 _6487_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5562__385 _5564__387/A vssd1 vssd1 vccd1 vccd1 _6675_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _4502_/A _4608_/B vssd1 vssd1 vccd1 vccd1 _4456_/S sky130_fd_sc_hd__or2_2
X_4371_ _4371_/A vssd1 vssd1 vccd1 vccd1 _6605_/D sky130_fd_sc_hd__clkbuf_1
X_7090_ _7096_/CLK _7090_/D vssd1 vssd1 vccd1 vccd1 _7090_/Q sky130_fd_sc_hd__dfxtp_4
X_3322_ _7127_/A _3242_/X _5047_/A vssd1 vssd1 vccd1 vccd1 _3936_/A sky130_fd_sc_hd__a21o_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6047_/A vssd1 vssd1 vccd1 vccd1 _6041_/X sky130_fd_sc_hd__buf_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3253_/A vssd1 vssd1 vccd1 vccd1 _7077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5771__471 _5773__473/A vssd1 vssd1 vccd1 vccd1 _6775_/CLK sky130_fd_sc_hd__inv_2
X_6943_ _6943_/CLK _6943_/D vssd1 vssd1 vccd1 vccd1 _6943_/Q sky130_fd_sc_hd__dfxtp_1
X_6874_ _7095_/CLK _6874_/D vssd1 vssd1 vccd1 vccd1 _6874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5756_ _5756_/A vssd1 vssd1 vccd1 vccd1 _5756_/X sky130_fd_sc_hd__buf_1
X_4707_ _4878_/S vssd1 vssd1 vccd1 vccd1 _4891_/B sky130_fd_sc_hd__buf_4
X_4638_ _3862_/X _6480_/Q _4642_/S vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4569_ _4569_/A vssd1 vssd1 vccd1 vccd1 _6511_/D sky130_fd_sc_hd__clkbuf_1
X_6308_ _7127_/A _6314_/B _6312_/C vssd1 vssd1 vccd1 vccd1 _6309_/A sky130_fd_sc_hd__and3_1
XFILLER_103_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6239_ _6239_/A vssd1 vssd1 vccd1 vccd1 _7004_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _3990_/C _3937_/Y _4562_/S vssd1 vssd1 vccd1 vccd1 _6776_/D sky130_fd_sc_hd__a21o_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3871_ _6748_/Q vssd1 vssd1 vccd1 vccd1 _3871_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5610_ _7083_/Q _7082_/Q _7081_/Q _5659_/B vssd1 vssd1 vccd1 vccd1 _5610_/X sky130_fd_sc_hd__or4_4
X_6590_ _6590_/CLK _6590_/D vssd1 vssd1 vccd1 vccd1 _6590_/Q sky130_fd_sc_hd__dfxtp_1
X_4423_ _4438_/S vssd1 vssd1 vccd1 vccd1 _4432_/S sky130_fd_sc_hd__buf_2
X_7142_ _7142_/A vssd1 vssd1 vccd1 vccd1 _7142_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4354_ _6612_/Q _3770_/A _4360_/S vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__mux2_1
X_3305_ _6774_/Q _6773_/Q _3315_/D vssd1 vssd1 vccd1 vccd1 _3941_/B sky130_fd_sc_hd__and3_1
XFILLER_59_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7073_ _7073_/CLK _7073_/D vssd1 vssd1 vccd1 vccd1 _7073_/Q sky130_fd_sc_hd__dfxtp_1
X_5209__261 _5210__262/A vssd1 vssd1 vccd1 vccd1 _6543_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6024_ _6023_/Y _6021_/Y _6013_/X vssd1 vssd1 vccd1 vccd1 _6888_/D sky130_fd_sc_hd__a21boi_1
X_4285_ _4285_/A vssd1 vssd1 vccd1 vccd1 _6643_/D sky130_fd_sc_hd__clkbuf_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _6459_/Q _6460_/Q _6461_/Q _6462_/Q vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__or4_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _6926_/CLK _6926_/D vssd1 vssd1 vccd1 vccd1 _6926_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3021_ clkbuf_0__3021_/X vssd1 vssd1 vccd1 vccd1 _6152__9/A sky130_fd_sc_hd__clkbuf_4
X_6857_ _6857_/CLK _6857_/D vssd1 vssd1 vccd1 vccd1 _6857_/Q sky130_fd_sc_hd__dfxtp_1
X_5513__346 _5514__347/A vssd1 vssd1 vccd1 vccd1 _6636_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6788_ _6788_/CLK _6788_/D vssd1 vssd1 vccd1 vccd1 _6788_/Q sky130_fd_sc_hd__dfxtp_1
X_5739_ _6897_/Q _6318_/B _5739_/C _7079_/Q vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__and4b_1
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2736_ clkbuf_0__2736_/X vssd1 vssd1 vccd1 vccd1 _5504__339/A sky130_fd_sc_hd__clkbuf_4
X_5594__407 _5594__407/A vssd1 vssd1 vccd1 vccd1 _6700_/CLK sky130_fd_sc_hd__inv_2
X_5881__77 _5882__78/A vssd1 vssd1 vccd1 vccd1 _6863_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_51 _7056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_40 _5739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6043__96 _6043__96/A vssd1 vssd1 vccd1 vccd1 _6904_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _4070_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__2871_ clkbuf_0__2871_/X vssd1 vssd1 vccd1 vccd1 _5845__529/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4972_ _4888_/X input34/X _4970_/X _5663_/A vssd1 vssd1 vccd1 vccd1 _4972_/X sky130_fd_sc_hd__a22o_2
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6711_ _6711_/CLK _6711_/D vssd1 vssd1 vccd1 vccd1 _6711_/Q sky130_fd_sc_hd__dfxtp_1
X_3923_ _3923_/A vssd1 vssd1 vccd1 vccd1 _6785_/D sky130_fd_sc_hd__clkbuf_1
X_3854_ _6809_/Q _3853_/X _3860_/S vssd1 vssd1 vccd1 vccd1 _3855_/A sky130_fd_sc_hd__mux2_1
X_6642_ _6642_/CLK _6642_/D vssd1 vssd1 vccd1 vccd1 _6642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6573_ _6573_/CLK _6573_/D vssd1 vssd1 vccd1 vccd1 _6573_/Q sky130_fd_sc_hd__dfxtp_1
X_3785_ _3785_/A vssd1 vssd1 vccd1 vccd1 _3785_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5455_ _5461_/A vssd1 vssd1 vccd1 vccd1 _5455_/X sky130_fd_sc_hd__buf_1
X_4406_ _3200_/X _6589_/Q _4414_/S vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__mux2_1
X_7125_ _7125_/A vssd1 vssd1 vccd1 vccd1 _7125_/X sky130_fd_sc_hd__clkbuf_1
X_5386_ _5324_/X _5375_/X _5385_/Y vssd1 vssd1 vccd1 vccd1 _5386_/X sky130_fd_sc_hd__a21o_1
XFILLER_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4337_ _4337_/A vssd1 vssd1 vccd1 vccd1 _6620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2521_ clkbuf_0__2521_/X vssd1 vssd1 vccd1 vccd1 _5179__237/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7056_ _7056_/CLK _7056_/D vssd1 vssd1 vccd1 vccd1 _7056_/Q sky130_fd_sc_hd__dfxtp_1
X_4268_ _4268_/A vssd1 vssd1 vccd1 vccd1 _6650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6007_ _6005_/X _6019_/B _6007_/C vssd1 vssd1 vccd1 vccd1 _6008_/A sky130_fd_sc_hd__and3b_1
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3219_ _3226_/A _3623_/B _4068_/C vssd1 vssd1 vccd1 vccd1 _3227_/B sky130_fd_sc_hd__o21a_1
X_4199_ _4199_/A vssd1 vssd1 vccd1 vccd1 _6680_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6909_ _6909_/CLK _6909_/D vssd1 vssd1 vccd1 vccd1 _6909_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__3004_ clkbuf_0__3004_/X vssd1 vssd1 vccd1 vccd1 _6064__113/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3570_ _3570_/A vssd1 vssd1 vccd1 vccd1 _6942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6334__23 _6334__23/A vssd1 vssd1 vccd1 vccd1 _7043_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _4122_/A vssd1 vssd1 vccd1 vccd1 _6714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4053_ _4053_/A vssd1 vssd1 vccd1 vccd1 _6735_/D sky130_fd_sc_hd__clkbuf_1
Xinput3 caravel_wb_data_i[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6113__153 _6113__153/A vssd1 vssd1 vccd1 vccd1 _6961_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__2854_ clkbuf_0__2854_/X vssd1 vssd1 vccd1 vccd1 _5778_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _6549_/Q _6729_/Q _6867_/Q _6533_/Q _4906_/X _3966_/X vssd1 vssd1 vccd1 vccd1
+ _4955_/X sky130_fd_sc_hd__mux4_1
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3906_ _6792_/Q _3608_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__mux2_1
X_4886_ _4884_/X _4885_/X _4969_/A vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6625_ _6625_/CLK _6625_/D vssd1 vssd1 vccd1 vccd1 _6625_/Q sky130_fd_sc_hd__dfxtp_1
X_3837_ _6815_/Q _3611_/X _3837_/S vssd1 vssd1 vccd1 vccd1 _3838_/A sky130_fd_sc_hd__mux2_1
X_6556_ _6556_/CLK _6556_/D vssd1 vssd1 vccd1 vccd1 _6556_/Q sky130_fd_sc_hd__dfxtp_1
X_3768_ _3764_/X _6843_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3769_/A sky130_fd_sc_hd__mux2_1
X_3699_ _4026_/A vssd1 vssd1 vccd1 vccd1 _3699_/X sky130_fd_sc_hd__buf_2
X_6487_ _6487_/CLK _6487_/D vssd1 vssd1 vccd1 vccd1 _6487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5438_ _6929_/Q _6921_/Q _7038_/Q _7054_/Q _5311_/X _5341_/X vssd1 vssd1 vccd1 vccd1
+ _5438_/X sky130_fd_sc_hd__mux4_2
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5369_ _7075_/Q _6701_/Q _6570_/Q _6848_/Q _5251_/X _5254_/X vssd1 vssd1 vccd1 vccd1
+ _5369_/X sky130_fd_sc_hd__mux4_1
X_7108_ _7108_/A vssd1 vssd1 vccd1 vccd1 _7108_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7039_ _7039_/CLK _7039_/D vssd1 vssd1 vccd1 vccd1 _7039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _4750_/A vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4671_ _4671_/A vssd1 vssd1 vccd1 vccd1 _6440_/D sky130_fd_sc_hd__clkbuf_1
X_6410_ _6427_/A _6427_/C vssd1 vssd1 vccd1 vccd1 _6432_/S sky130_fd_sc_hd__nand2_2
X_3622_ _3622_/A vssd1 vssd1 vccd1 vccd1 _6922_/D sky130_fd_sc_hd__clkbuf_1
X_3553_ _6949_/Q _3453_/X _3553_/S vssd1 vssd1 vccd1 vccd1 _3554_/A sky130_fd_sc_hd__mux2_1
X_6272_ _6272_/A _6272_/B vssd1 vssd1 vccd1 vccd1 _6280_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3484_ _3484_/A vssd1 vssd1 vccd1 vccd1 _3485_/B sky130_fd_sc_hd__inv_2
XFILLER_115_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3021_ _6147_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3021_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4105_ _4590_/A _4123_/B vssd1 vssd1 vccd1 vccd1 _4121_/S sky130_fd_sc_hd__nor2_2
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5085_ _6459_/Q _7113_/A _5093_/S vssd1 vssd1 vccd1 vccd1 _5086_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4036_ _4036_/A vssd1 vssd1 vccd1 vccd1 _6305_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2837_ clkbuf_0__2837_/X vssd1 vssd1 vccd1 vccd1 _5705__435/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5987_ _6879_/Q _5966_/X _5986_/Y _5970_/X vssd1 vssd1 vccd1 vccd1 _5988_/B sky130_fd_sc_hd__a22o_1
X_4938_ _6548_/Q _6728_/Q _6866_/Q _6532_/Q _4906_/X _3966_/X vssd1 vssd1 vccd1 vccd1
+ _4938_/X sky130_fd_sc_hd__mux4_1
X_4869_ _4808_/A _4868_/X _4732_/A vssd1 vssd1 vccd1 vccd1 _4869_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_0__2736_ _5499_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2736_/X sky130_fd_sc_hd__clkbuf_16
X_6608_ _6608_/CLK _6608_/D vssd1 vssd1 vccd1 vccd1 _6608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6539_ _6539_/CLK _6539_/D vssd1 vssd1 vccd1 vccd1 _6539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput170 _7158_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput181 _4983_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput192 _5004_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[24] sky130_fd_sc_hd__buf_2
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6062__111 _6064__113/A vssd1 vssd1 vccd1 vccd1 _6919_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5910_ _5910_/A _6871_/Q vssd1 vssd1 vccd1 vccd1 _5911_/S sky130_fd_sc_hd__xor2_1
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6890_ _6890_/CLK _6890_/D vssd1 vssd1 vccd1 vccd1 _6890_/Q sky130_fd_sc_hd__dfxtp_1
X_4723_ _4826_/A _4720_/X _4722_/X vssd1 vssd1 vccd1 vccd1 _4723_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_0__2521_ _5176_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2521_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4654_ _3859_/X _6473_/Q _4654_/S vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4585_ _4585_/A vssd1 vssd1 vccd1 vccd1 _6504_/D sky130_fd_sc_hd__clkbuf_1
X_3605_ _7028_/Q vssd1 vssd1 vccd1 vccd1 _3605_/X sky130_fd_sc_hd__buf_6
Xinput61 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 _7100_/A sky130_fd_sc_hd__buf_4
Xinput72 wbs_data_i[12] vssd1 vssd1 vccd1 vccd1 _7137_/A sky130_fd_sc_hd__buf_4
Xinput50 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 _7119_/A sky130_fd_sc_hd__buf_4
XFILLER_115_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6324_ _6330_/A vssd1 vssd1 vccd1 vccd1 _6324_/X sky130_fd_sc_hd__buf_1
Xinput94 wbs_data_i[3] vssd1 vssd1 vccd1 vccd1 _7128_/A sky130_fd_sc_hd__buf_8
Xinput83 wbs_data_i[22] vssd1 vssd1 vccd1 vccd1 _7147_/A sky130_fd_sc_hd__buf_4
X_3536_ _6956_/Q _3456_/X _3540_/S vssd1 vssd1 vccd1 vccd1 _3537_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6255_ _6258_/B vssd1 vssd1 vccd1 vccd1 _6255_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5206_ _5206_/A vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__buf_1
X_3467_ _3482_/S vssd1 vssd1 vccd1 vccd1 _3476_/S sky130_fd_sc_hd__buf_2
X_6186_ _6187_/B _6187_/C _6245_/B vssd1 vssd1 vccd1 vccd1 _6188_/B sky130_fd_sc_hd__o21ai_1
X_3398_ _4502_/A vssd1 vssd1 vccd1 vccd1 _4590_/A sky130_fd_sc_hd__buf_4
Xclkbuf_0__3004_ _6060_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3004_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5068_ _5068_/A vssd1 vssd1 vccd1 vccd1 _6451_/D sky130_fd_sc_hd__clkbuf_1
X_4019_ _4019_/A vssd1 vssd1 vccd1 vccd1 _6756_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6126__163 _6127__164/A vssd1 vssd1 vccd1 vccd1 _6971_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _6605_/Q _3764_/A _4378_/S vssd1 vssd1 vccd1 vccd1 _4371_/A sky130_fd_sc_hd__mux2_1
X_3321_ _3948_/A _3948_/B vssd1 vssd1 vccd1 vccd1 _3949_/A sky130_fd_sc_hd__nand2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _7077_/Q _3251_/X _3261_/S vssd1 vssd1 vccd1 vccd1 _3253_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6069__117 _6069__117/A vssd1 vssd1 vccd1 vccd1 _6925_/CLK sky130_fd_sc_hd__inv_2
X_6942_ _6942_/CLK _6942_/D vssd1 vssd1 vccd1 vccd1 _6942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6873_ _7008_/CLK _6873_/D vssd1 vssd1 vccd1 vccd1 _6873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4706_ _4868_/S vssd1 vssd1 vccd1 vccd1 _4878_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_118_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4637_ _4637_/A vssd1 vssd1 vccd1 vccd1 _6481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4568_ _6511_/Q _4029_/A _4570_/S vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4499_ _6741_/Q vssd1 vssd1 vccd1 vccd1 _4499_/X sky130_fd_sc_hd__clkbuf_4
X_6307_ _6307_/A vssd1 vssd1 vccd1 vccd1 _7024_/D sky130_fd_sc_hd__clkbuf_1
X_3519_ _3519_/A vssd1 vssd1 vccd1 vccd1 _6964_/D sky130_fd_sc_hd__clkbuf_1
X_6238_ _6238_/A _6238_/B _6238_/C vssd1 vssd1 vccd1 vccd1 _6239_/A sky130_fd_sc_hd__and3_1
Xclkbuf_1_1_0__3019_ clkbuf_0__3019_/X vssd1 vssd1 vccd1 vccd1 _6145__179/A sky130_fd_sc_hd__clkbuf_4
X_6169_ _6161_/A _6166_/Y _7002_/Q _6167_/Y _6168_/Y vssd1 vssd1 vccd1 vccd1 _6172_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _3870_/A vssd1 vssd1 vccd1 vccd1 _6804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4422_ _4422_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _4438_/S sky130_fd_sc_hd__or2_2
X_7141_ _7141_/A vssd1 vssd1 vccd1 vccd1 _7141_/X sky130_fd_sc_hd__clkbuf_1
X_4353_ _4353_/A vssd1 vssd1 vccd1 vccd1 _6613_/D sky130_fd_sc_hd__clkbuf_1
X_3304_ _3315_/D vssd1 vssd1 vccd1 vccd1 _3948_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4284_ _6643_/Q _4149_/X _4288_/S vssd1 vssd1 vccd1 vccd1 _4285_/A sky130_fd_sc_hd__mux2_1
X_7072_ _7072_/CLK _7072_/D vssd1 vssd1 vccd1 vccd1 _7072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3235_ _6446_/Q _5113_/B _6445_/Q vssd1 vssd1 vccd1 vccd1 _3240_/C sky130_fd_sc_hd__or3b_1
X_6023_ _6888_/Q vssd1 vssd1 vccd1 vccd1 _6023_/Y sky130_fd_sc_hd__inv_2
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _6925_/CLK _6925_/D vssd1 vssd1 vccd1 vccd1 _6925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3020_ clkbuf_0__3020_/X vssd1 vssd1 vccd1 vccd1 _6336_/A sky130_fd_sc_hd__clkbuf_4
X_6856_ _6856_/CLK _6856_/D vssd1 vssd1 vccd1 vccd1 _6856_/Q sky130_fd_sc_hd__dfxtp_1
X_3999_ _3693_/X _6763_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _4000_/A sky130_fd_sc_hd__mux2_1
X_6787_ _6787_/CLK _6787_/D vssd1 vssd1 vccd1 vccd1 _6787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2519_ clkbuf_0__2519_/X vssd1 vssd1 vccd1 vccd1 _5174__234/A sky130_fd_sc_hd__clkbuf_4
X_5738_ _5738_/A vssd1 vssd1 vccd1 vccd1 _6749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5669_ _5669_/A _5669_/B _5669_/C _5668_/X vssd1 vssd1 vccd1 vccd1 _6271_/A sky130_fd_sc_hd__or4b_4
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_30 _3853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_41 _4146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6346__32 _6347__33/A vssd1 vssd1 vccd1 vccd1 _7052_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2870_ clkbuf_0__2870_/X vssd1 vssd1 vccd1 vccd1 _5839__524/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5575__396 _5578__399/A vssd1 vssd1 vccd1 vccd1 _6686_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4971_ _7087_/Q vssd1 vssd1 vccd1 vccd1 _5663_/A sky130_fd_sc_hd__buf_4
X_6710_ _6710_/CLK _6710_/D vssd1 vssd1 vccd1 vccd1 _6710_/Q sky130_fd_sc_hd__dfxtp_1
X_3922_ _6785_/Q _3880_/X _3926_/S vssd1 vssd1 vccd1 vccd1 _3923_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3853_ _6746_/Q vssd1 vssd1 vccd1 vccd1 _3853_/X sky130_fd_sc_hd__buf_4
X_6641_ _6641_/CLK _6641_/D vssd1 vssd1 vccd1 vccd1 _6641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6572_ _6572_/CLK _6572_/D vssd1 vssd1 vccd1 vccd1 _6572_/Q sky130_fd_sc_hd__dfxtp_1
X_3784_ _3784_/A vssd1 vssd1 vccd1 vccd1 _6838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5523_ _5523_/A vssd1 vssd1 vccd1 vccd1 _5523_/X sky130_fd_sc_hd__buf_1
XFILLER_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4405_ _4420_/S vssd1 vssd1 vccd1 vccd1 _4414_/S sky130_fd_sc_hd__clkbuf_2
X_5385_ _5366_/A _5384_/X _5250_/A vssd1 vssd1 vccd1 vccd1 _5385_/Y sky130_fd_sc_hd__o21ai_1
X_7124_ _7124_/A vssd1 vssd1 vccd1 vccd1 _7124_/X sky130_fd_sc_hd__clkbuf_1
X_4336_ _3770_/X _6620_/Q _4342_/S vssd1 vssd1 vccd1 vccd1 _4337_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__2520_ clkbuf_0__2520_/X vssd1 vssd1 vccd1 vccd1 _5188_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7055_ _7055_/CLK _7055_/D vssd1 vssd1 vccd1 vccd1 _7055_/Q sky130_fd_sc_hd__dfxtp_2
X_4267_ _6650_/Q _4152_/X _4269_/S vssd1 vssd1 vccd1 vccd1 _4268_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4198_ _6680_/Q _4158_/X _4202_/S vssd1 vssd1 vccd1 vccd1 _4199_/A sky130_fd_sc_hd__mux2_1
X_6006_ _6882_/Q _5970_/A _6004_/C _6883_/Q vssd1 vssd1 vccd1 vccd1 _6007_/C sky130_fd_sc_hd__a31o_1
X_3218_ _6739_/Q _6734_/Q vssd1 vssd1 vccd1 vccd1 _4068_/C sky130_fd_sc_hd__xor2_2
XFILLER_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__2999_ clkbuf_0__2999_/X vssd1 vssd1 vccd1 vccd1 _6040__94/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6908_ _6908_/CLK _6908_/D vssd1 vssd1 vccd1 vccd1 _6908_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3003_ clkbuf_0__3003_/X vssd1 vssd1 vccd1 vccd1 _6059__109/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6839_ _6839_/CLK _6839_/D vssd1 vssd1 vccd1 vccd1 _6839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5158__220 _5160__222/A vssd1 vssd1 vccd1 vccd1 _6502_/CLK sky130_fd_sc_hd__inv_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5462__305 _5464__307/A vssd1 vssd1 vccd1 vccd1 _6595_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4121_ _6714_/Q _3895_/X _4121_/S vssd1 vssd1 vccd1 vccd1 _4122_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4052_ _6303_/B _4052_/B _4052_/C vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__and3_1
Xinput4 caravel_wb_data_i[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__2853_ clkbuf_0__2853_/X vssd1 vssd1 vccd1 vccd1 _5755__459/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5811__501 _5813__503/A vssd1 vssd1 vccd1 vccd1 _6807_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4954_ _4952_/X _4953_/X _4954_/S vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3905_ _3905_/A vssd1 vssd1 vccd1 vccd1 _6793_/D sky130_fd_sc_hd__clkbuf_1
X_4885_ _7092_/Q vssd1 vssd1 vccd1 vccd1 _4885_/X sky130_fd_sc_hd__clkbuf_4
X_6624_ _6624_/CLK _6624_/D vssd1 vssd1 vccd1 vccd1 _6624_/Q sky130_fd_sc_hd__dfxtp_1
X_3836_ _3836_/A vssd1 vssd1 vccd1 vccd1 _6816_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6555_ _6555_/CLK _6555_/D vssd1 vssd1 vccd1 vccd1 _6555_/Q sky130_fd_sc_hd__dfxtp_1
X_3767_ _3789_/S vssd1 vssd1 vccd1 vccd1 _3780_/S sky130_fd_sc_hd__buf_2
X_6120__158 _6121__159/A vssd1 vssd1 vccd1 vccd1 _6966_/CLK sky130_fd_sc_hd__inv_2
XFILLER_118_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3698_ _3698_/A vssd1 vssd1 vccd1 vccd1 _6892_/D sky130_fd_sc_hd__clkbuf_1
X_6486_ _6486_/CLK _6486_/D vssd1 vssd1 vccd1 vccd1 _6486_/Q sky130_fd_sc_hd__dfxtp_1
X_5437_ _5437_/A _5437_/B vssd1 vssd1 vccd1 vccd1 _5437_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5368_ _6577_/Q _5250_/X _5367_/Y _5298_/X vssd1 vssd1 vccd1 vccd1 _6577_/D sky130_fd_sc_hd__o211a_1
X_7107_ _7107_/A vssd1 vssd1 vccd1 vccd1 _7107_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4319_ _4319_/A vssd1 vssd1 vccd1 vccd1 _6628_/D sky130_fd_sc_hd__clkbuf_1
X_5299_ _6574_/Q _5250_/X _5296_/X _5298_/X vssd1 vssd1 vccd1 vccd1 _6574_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7038_ _7038_/CLK _7038_/D vssd1 vssd1 vccd1 vccd1 _7038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5526__357 _5527__358/A vssd1 vssd1 vccd1 vccd1 _6647_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4670_ _3856_/X _6440_/Q _4672_/S vssd1 vssd1 vccd1 vccd1 _4671_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3621_ _6922_/Q _3620_/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3622_/A sky130_fd_sc_hd__mux2_1
X_3552_ _3552_/A vssd1 vssd1 vccd1 vccd1 _6950_/D sky130_fd_sc_hd__clkbuf_1
X_6271_ _6271_/A _6271_/B vssd1 vssd1 vccd1 vccd1 _6271_/X sky130_fd_sc_hd__and2_1
X_3483_ _3483_/A vssd1 vssd1 vccd1 vccd1 _6978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3020_ _6146_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3020_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4104_ _4104_/A vssd1 vssd1 vccd1 vccd1 _6722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5084_ _5588_/S vssd1 vssd1 vccd1 vccd1 _5093_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4035_ _4051_/B vssd1 vssd1 vccd1 vccd1 _4035_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5986_ _5994_/C _5986_/B vssd1 vssd1 vccd1 vccd1 _5986_/Y sky130_fd_sc_hd__nor2_1
X_4937_ _4774_/X _4936_/X _4905_/A vssd1 vssd1 vccd1 vccd1 _4937_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4868_ _6474_/Q _7059_/Q _4868_/S vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2735_ _5498_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2735_/X sky130_fd_sc_hd__clkbuf_16
X_3819_ _6823_/Q _3611_/X _3819_/S vssd1 vssd1 vccd1 vccd1 _3820_/A sky130_fd_sc_hd__mux2_1
X_6607_ _6607_/CLK _6607_/D vssd1 vssd1 vccd1 vccd1 _6607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4799_ _4765_/Y _4766_/Y _4784_/X _4797_/Y _4798_/Y vssd1 vssd1 vccd1 vccd1 _4799_/X
+ sky130_fd_sc_hd__a221o_1
X_6538_ _6538_/CLK _6538_/D vssd1 vssd1 vccd1 vccd1 _6538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6469_ _6696_/CLK _6469_/D vssd1 vssd1 vccd1 vccd1 _6469_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput160 _7155_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[30] sky130_fd_sc_hd__buf_2
XFILLER_79_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput171 _7159_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[2] sky130_fd_sc_hd__buf_2
Xoutput193 _5007_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput182 _4986_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[15] sky130_fd_sc_hd__buf_2
XFILLER_101_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5818__507 _5820__509/A vssd1 vssd1 vccd1 vccd1 _6813_/CLK sky130_fd_sc_hd__inv_2
XFILLER_102_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5532__361 _5534__363/A vssd1 vssd1 vccd1 vccd1 _6651_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5203__257 _5205__259/A vssd1 vssd1 vccd1 vccd1 _6539_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5840_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5840_/X sky130_fd_sc_hd__buf_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4722_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4722_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__2520_ _5175_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2520_/X sky130_fd_sc_hd__clkbuf_16
X_4653_ _4653_/A vssd1 vssd1 vccd1 vccd1 _6474_/D sky130_fd_sc_hd__clkbuf_1
Xinput40 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 _7110_/A sky130_fd_sc_hd__buf_4
X_4584_ _4493_/X _6504_/Q _4588_/S vssd1 vssd1 vccd1 vccd1 _4585_/A sky130_fd_sc_hd__mux2_1
Xinput62 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 _7101_/A sky130_fd_sc_hd__buf_4
Xinput73 wbs_data_i[13] vssd1 vssd1 vccd1 vccd1 _7138_/A sky130_fd_sc_hd__buf_4
Xinput51 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 _7120_/A sky130_fd_sc_hd__buf_4
X_3604_ _3604_/A vssd1 vssd1 vccd1 vccd1 _6928_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput95 wbs_data_i[4] vssd1 vssd1 vccd1 vccd1 _7129_/A sky130_fd_sc_hd__buf_6
Xinput84 wbs_data_i[23] vssd1 vssd1 vccd1 vccd1 _7148_/A sky130_fd_sc_hd__buf_4
X_3535_ _3535_/A vssd1 vssd1 vccd1 vccd1 _6957_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6254_ _7007_/Q _7006_/Q _6254_/C _6254_/D vssd1 vssd1 vccd1 vccd1 _6258_/B sky130_fd_sc_hd__and4_1
X_3466_ _4404_/A _3898_/B vssd1 vssd1 vccd1 vccd1 _3482_/S sky130_fd_sc_hd__or2_2
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6185_ _6272_/A vssd1 vssd1 vccd1 vccd1 _6245_/B sky130_fd_sc_hd__inv_2
XFILLER_69_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3397_ _3948_/A _3661_/C _3661_/A vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__or3b_4
Xclkbuf_0__3003_ _6054_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3003_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_96_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5067_ _6451_/Q _7105_/A _5071_/S vssd1 vssd1 vccd1 vccd1 _5068_/A sky130_fd_sc_hd__mux2_1
X_4018_ _4017_/X _6756_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4019_/A sky130_fd_sc_hd__mux2_1
X_5475__315 _5479__319/A vssd1 vssd1 vccd1 vccd1 _6605_/CLK sky130_fd_sc_hd__inv_2
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5969_ _5969_/A _5978_/C vssd1 vssd1 vccd1 vccd1 _5969_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5824__511 _5825__512/A vssd1 vssd1 vccd1 vccd1 _6817_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3320_ _3484_/A vssd1 vssd1 vccd1 vccd1 _3948_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3251_ _7029_/Q vssd1 vssd1 vccd1 vccd1 _3251_/X sky130_fd_sc_hd__buf_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6941_ _6941_/CLK _6941_/D vssd1 vssd1 vccd1 vccd1 _6941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5539__367 _5541__369/A vssd1 vssd1 vccd1 vccd1 _6657_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6872_ _7095_/CLK _6872_/D vssd1 vssd1 vccd1 vccd1 _6872_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2535_ clkbuf_0__2535_/X vssd1 vssd1 vccd1 vccd1 _5448__294/A sky130_fd_sc_hd__clkbuf_4
X_5685_ _5685_/A vssd1 vssd1 vccd1 vccd1 _5685_/X sky130_fd_sc_hd__buf_1
X_4705_ _4875_/S vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4636_ _3859_/X _6481_/Q _4636_/S vssd1 vssd1 vccd1 vccd1 _4637_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4567_ _4567_/A vssd1 vssd1 vccd1 vccd1 _6512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6306_ _7126_/A _6314_/B _6312_/C vssd1 vssd1 vccd1 vccd1 _6307_/A sky130_fd_sc_hd__and3_1
X_4498_ _4498_/A vssd1 vssd1 vccd1 vccd1 _6543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2751_ clkbuf_0__2751_/X vssd1 vssd1 vccd1 vccd1 _5590__404/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3518_ _6964_/Q _3456_/X _3522_/S vssd1 vssd1 vccd1 vccd1 _3519_/A sky130_fd_sc_hd__mux2_1
X_6237_ _7004_/Q _6241_/B _6237_/C vssd1 vssd1 vccd1 vccd1 _6238_/C sky130_fd_sc_hd__nand3_1
X_3449_ _3449_/A vssd1 vssd1 vccd1 vccd1 _6991_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3018_ clkbuf_0__3018_/X vssd1 vssd1 vccd1 vccd1 _6137__172/A sky130_fd_sc_hd__clkbuf_4
X_6168_ _6168_/A _6168_/B vssd1 vssd1 vccd1 vccd1 _6168_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5748__453 _5749__454/A vssd1 vssd1 vccd1 vccd1 _6757_/CLK sky130_fd_sc_hd__inv_2
X_5152__215 _5155__218/A vssd1 vssd1 vccd1 vccd1 _6497_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4421_ _4421_/A vssd1 vssd1 vccd1 vccd1 _6582_/D sky130_fd_sc_hd__clkbuf_1
X_7140_ _7140_/A vssd1 vssd1 vccd1 vccd1 _7140_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4352_ _6613_/Q _3764_/A _4360_/S vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__mux2_1
X_6075__122 _6075__122/A vssd1 vssd1 vccd1 vccd1 _6930_/CLK sky130_fd_sc_hd__inv_2
X_3303_ _6772_/Q vssd1 vssd1 vccd1 vccd1 _3315_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4283_ _4283_/A vssd1 vssd1 vccd1 vccd1 _6644_/D sky130_fd_sc_hd__clkbuf_1
X_7071_ _7071_/CLK _7071_/D vssd1 vssd1 vccd1 vccd1 _7071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3234_ _6469_/Q _6468_/Q vssd1 vssd1 vccd1 vccd1 _5113_/B sky130_fd_sc_hd__nor2_2
X_6022_ _6887_/Q _6021_/B _6021_/Y _6013_/X vssd1 vssd1 vccd1 vccd1 _6887_/D sky130_fd_sc_hd__o211a_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6924_ _6924_/CLK _6924_/D vssd1 vssd1 vccd1 vccd1 _6924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6855_ _6855_/CLK _6855_/D vssd1 vssd1 vccd1 vccd1 _6855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3998_ _3998_/A vssd1 vssd1 vccd1 vccd1 _6764_/D sky130_fd_sc_hd__clkbuf_1
X_6786_ _6786_/CLK _6786_/D vssd1 vssd1 vccd1 vccd1 _6786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5737_ _5046_/B _6318_/C _6305_/A _5737_/D vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__and4b_1
X_5216__267 _5216__267/A vssd1 vssd1 vccd1 vccd1 _6549_/CLK sky130_fd_sc_hd__inv_2
X_5668_ _7005_/Q _5623_/X _5662_/X _5666_/X _5667_/Y vssd1 vssd1 vccd1 vccd1 _5668_/X
+ sky130_fd_sc_hd__o2111a_1
X_4619_ _4619_/A vssd1 vssd1 vccd1 vccd1 _6489_/D sky130_fd_sc_hd__clkbuf_1
X_5599_ _5685_/A vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__buf_1
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2734_ clkbuf_0__2734_/X vssd1 vssd1 vccd1 vccd1 _5494__331/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_31 _3856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_20 _7062_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_42 _4146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6139__174 _6139__174/A vssd1 vssd1 vccd1 vccd1 _6982_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4970_ _4970_/A vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3921_ _3921_/A vssd1 vssd1 vccd1 vccd1 _6786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3852_ _3852_/A vssd1 vssd1 vccd1 vccd1 _6810_/D sky130_fd_sc_hd__clkbuf_1
X_6640_ _6640_/CLK _6640_/D vssd1 vssd1 vccd1 vccd1 _6640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6571_ _6571_/CLK _6571_/D vssd1 vssd1 vccd1 vccd1 _6571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3783_ _3782_/X _6838_/Q _3789_/S vssd1 vssd1 vccd1 vccd1 _3784_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4404_ _4404_/A _4404_/B vssd1 vssd1 vccd1 vccd1 _4420_/S sky130_fd_sc_hd__or2_2
X_5384_ _5334_/X _5377_/X _5379_/Y _5381_/X _5383_/Y vssd1 vssd1 vccd1 vccd1 _5384_/X
+ sky130_fd_sc_hd__o32a_2
X_7123_ _7123_/A vssd1 vssd1 vccd1 vccd1 _7123_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4335_ _4335_/A vssd1 vssd1 vccd1 vccd1 _6621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7054_ _7054_/CLK _7054_/D vssd1 vssd1 vccd1 vccd1 _7054_/Q sky130_fd_sc_hd__dfxtp_1
X_4266_ _4266_/A vssd1 vssd1 vccd1 vccd1 _6651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6005_ _5953_/B _6012_/B _5944_/X vssd1 vssd1 vccd1 vccd1 _6005_/X sky130_fd_sc_hd__o21ba_1
X_4197_ _4197_/A vssd1 vssd1 vccd1 vccd1 _6681_/D sky130_fd_sc_hd__clkbuf_1
X_3217_ _4204_/A _6737_/Q vssd1 vssd1 vccd1 vccd1 _3623_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1_0__2998_ clkbuf_0__2998_/X vssd1 vssd1 vccd1 vccd1 _6033__89/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6907_ _6907_/CLK _6907_/D vssd1 vssd1 vccd1 vccd1 _6907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__3002_ clkbuf_0__3002_/X vssd1 vssd1 vccd1 vccd1 _6078_/A sky130_fd_sc_hd__clkbuf_4
X_6838_ _6838_/CLK _6838_/D vssd1 vssd1 vccd1 vccd1 _6838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6769_ _6769_/CLK _6769_/D vssd1 vssd1 vccd1 vccd1 _6769_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_104_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4120_ _4120_/A vssd1 vssd1 vccd1 vccd1 _6715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4051_ _4051_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _4052_/C sky130_fd_sc_hd__or2_1
Xinput5 caravel_wb_data_i[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__2852_ clkbuf_0__2852_/X vssd1 vssd1 vccd1 vccd1 _5749__454/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4953_ _6905_/Q _6565_/Q _6913_/Q _6493_/Q _4906_/X _4772_/S vssd1 vssd1 vccd1 vccd1
+ _4953_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2751_ _5579_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2751_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3904_ _6793_/Q _3605_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3905_/A sky130_fd_sc_hd__mux2_1
X_6623_ _6623_/CLK _6623_/D vssd1 vssd1 vccd1 vccd1 _6623_/Q sky130_fd_sc_hd__dfxtp_1
X_4884_ _4856_/Y _4872_/X _4882_/X _4883_/Y vssd1 vssd1 vccd1 vccd1 _4884_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3835_ _6816_/Q _3608_/X _3837_/S vssd1 vssd1 vccd1 vccd1 _3836_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6554_ _6554_/CLK _6554_/D vssd1 vssd1 vccd1 vccd1 _6554_/Q sky130_fd_sc_hd__dfxtp_1
X_3766_ _4186_/A _4404_/B vssd1 vssd1 vccd1 vccd1 _3789_/S sky130_fd_sc_hd__or2_2
XFILLER_118_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6485_ _6485_/CLK _6485_/D vssd1 vssd1 vccd1 vccd1 _6485_/Q sky130_fd_sc_hd__dfxtp_1
X_5505_ _5523_/A vssd1 vssd1 vccd1 vccd1 _5505_/X sky130_fd_sc_hd__buf_1
XFILLER_106_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3697_ _3696_/X _6892_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3698_/A sky130_fd_sc_hd__mux2_1
X_5436_ _6953_/Q _6685_/Q _6597_/Q _6819_/Q _5337_/X _5338_/X vssd1 vssd1 vccd1 vccd1
+ _5437_/B sky130_fd_sc_hd__mux4_1
X_6340__28 _6341__29/A vssd1 vssd1 vccd1 vccd1 _7048_/CLK sky130_fd_sc_hd__inv_2
X_5367_ _4055_/X _5358_/X _5366_/Y _5321_/X vssd1 vssd1 vccd1 vccd1 _5367_/Y sky130_fd_sc_hd__o211ai_1
X_7106_ _7106_/A vssd1 vssd1 vccd1 vccd1 _7106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4318_ _6628_/Q _3877_/X _4324_/S vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5298_ _6019_/B vssd1 vssd1 vccd1 vccd1 _5298_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7037_ _7037_/CLK _7037_/D vssd1 vssd1 vccd1 vccd1 _7037_/Q sky130_fd_sc_hd__dfxtp_1
X_4249_ _3776_/X _6658_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6088__132 _6088__132/A vssd1 vssd1 vccd1 vccd1 _6940_/CLK sky130_fd_sc_hd__inv_2
XFILLER_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5687__421 _5688__422/A vssd1 vssd1 vccd1 vccd1 _6715_/CLK sky130_fd_sc_hd__inv_2
XFILLER_42_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3620_ _7023_/Q vssd1 vssd1 vccd1 vccd1 _3620_/X sky130_fd_sc_hd__buf_4
X_3551_ _6950_/Q _3450_/X _3553_/S vssd1 vssd1 vccd1 vccd1 _3552_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6270_ _6270_/A _6270_/B vssd1 vssd1 vccd1 vccd1 _7011_/D sky130_fd_sc_hd__nor2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3482_ _3392_/X _6978_/Q _3482_/S vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4103_ _4032_/X _6722_/Q _4103_/S vssd1 vssd1 vccd1 vccd1 _4104_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5083_ _5083_/A vssd1 vssd1 vccd1 vccd1 _6458_/D sky130_fd_sc_hd__clkbuf_1
X_4034_ _4034_/A vssd1 vssd1 vccd1 vccd1 _6751_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__2835_ clkbuf_0__2835_/X vssd1 vssd1 vccd1 vccd1 _5702__434/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5985_ _6879_/Q _5985_/B vssd1 vssd1 vccd1 vccd1 _5986_/B sky130_fd_sc_hd__nor2_1
X_4936_ _6895_/Q _6524_/Q _4936_/S vssd1 vssd1 vccd1 vccd1 _4936_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4867_ _6626_/Q _6784_/Q _4878_/S vssd1 vssd1 vccd1 vccd1 _4867_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_0__2734_ _5492_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2734_/X sky130_fd_sc_hd__clkbuf_16
X_3818_ _3818_/A vssd1 vssd1 vccd1 vccd1 _6824_/D sky130_fd_sc_hd__clkbuf_1
X_6606_ _6606_/CLK _6606_/D vssd1 vssd1 vccd1 vccd1 _6606_/Q sky130_fd_sc_hd__dfxtp_1
X_6537_ _6537_/CLK _6537_/D vssd1 vssd1 vccd1 vccd1 _6537_/Q sky130_fd_sc_hd__dfxtp_1
X_4798_ _4798_/A _4798_/B vssd1 vssd1 vccd1 vccd1 _4798_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3749_ _3749_/A vssd1 vssd1 vccd1 vccd1 _6851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5742__448 _5743__449/A vssd1 vssd1 vccd1 vccd1 _6752_/CLK sky130_fd_sc_hd__inv_2
X_6468_ _7096_/CLK _6468_/D vssd1 vssd1 vccd1 vccd1 _6468_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput150 _7146_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[21] sky130_fd_sc_hd__buf_2
Xoutput161 _7156_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[31] sky130_fd_sc_hd__buf_2
X_6399_ _6408_/A _6399_/B vssd1 vssd1 vccd1 vccd1 _6400_/A sky130_fd_sc_hd__and2_1
X_5419_ _6928_/Q _6920_/Q _7037_/Q _7053_/Q _5311_/X _5341_/X vssd1 vssd1 vccd1 vccd1
+ _5419_/X sky130_fd_sc_hd__mux4_2
Xoutput172 _7160_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[3] sky130_fd_sc_hd__buf_2
XFILLER_87_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput194 _5009_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput183 _4988_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149__6 _6150__7/A vssd1 vssd1 vccd1 vccd1 _6989_/CLK sky130_fd_sc_hd__inv_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4721_ _6770_/Q vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__inv_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4652_ _3856_/X _6474_/Q _4654_/S vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__mux2_1
Xinput30 caravel_wb_data_i[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
X_3603_ _6928_/Q _3602_/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3604_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4583_ _4583_/A vssd1 vssd1 vccd1 vccd1 _6505_/D sky130_fd_sc_hd__clkbuf_1
Xinput41 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 _7111_/A sky130_fd_sc_hd__buf_4
Xinput52 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 _7121_/A sky130_fd_sc_hd__buf_4
Xinput63 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 _7102_/A sky130_fd_sc_hd__buf_4
Xclkbuf_4_5_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _5852_/A sky130_fd_sc_hd__clkbuf_4
Xinput96 wbs_data_i[5] vssd1 vssd1 vccd1 vccd1 _7130_/A sky130_fd_sc_hd__buf_6
Xinput74 wbs_data_i[14] vssd1 vssd1 vccd1 vccd1 _7139_/A sky130_fd_sc_hd__buf_4
Xinput85 wbs_data_i[24] vssd1 vssd1 vccd1 vccd1 _7149_/A sky130_fd_sc_hd__buf_4
X_3534_ _6957_/Q _3453_/X _3534_/S vssd1 vssd1 vccd1 vccd1 _3535_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6253_ _6253_/A vssd1 vssd1 vccd1 vccd1 _7006_/D sky130_fd_sc_hd__clkbuf_1
X_3465_ _4422_/B vssd1 vssd1 vccd1 vccd1 _4404_/A sky130_fd_sc_hd__clkbuf_4
X_6184_ _6272_/B _6184_/B vssd1 vssd1 vccd1 vccd1 _6187_/C sky130_fd_sc_hd__nor2_1
X_3396_ _3948_/B _3947_/A vssd1 vssd1 vccd1 vccd1 _3661_/C sky130_fd_sc_hd__nand2_1
Xclkbuf_0__3002_ _6053_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3002_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_111_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5066_ _5066_/A vssd1 vssd1 vccd1 vccd1 _6450_/D sky130_fd_sc_hd__clkbuf_1
X_4017_ _4017_/A vssd1 vssd1 vccd1 vccd1 _4017_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5968_ _6876_/Q _5968_/B vssd1 vssd1 vccd1 vccd1 _5978_/C sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__2749_ clkbuf_0__2749_/X vssd1 vssd1 vccd1 vccd1 _5569__391/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4919_ _6740_/Q _4766_/Y _4904_/X _4918_/Y _4798_/Y vssd1 vssd1 vccd1 vccd1 _4919_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5899_ _6884_/Q vssd1 vssd1 vccd1 vccd1 _6012_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6133__169 _6133__169/A vssd1 vssd1 vccd1 vccd1 _6977_/CLK sky130_fd_sc_hd__inv_2
XFILLER_48_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5580__400 _5583__403/A vssd1 vssd1 vccd1 vccd1 _6690_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3250_/A vssd1 vssd1 vccd1 vccd1 _7078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6940_ _6940_/CLK _6940_/D vssd1 vssd1 vccd1 vccd1 _6940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6871_ _6888_/CLK _6871_/D vssd1 vssd1 vccd1 vccd1 _6871_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__2757_ clkbuf_0__2757_/X vssd1 vssd1 vccd1 vccd1 _5685_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5822_ _5846_/A vssd1 vssd1 vccd1 vccd1 _5822_/X sky130_fd_sc_hd__buf_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2534_ clkbuf_0__2534_/X vssd1 vssd1 vccd1 vccd1 _5244__289/A sky130_fd_sc_hd__clkbuf_4
X_4704_ _6769_/Q vssd1 vssd1 vccd1 vccd1 _4875_/S sky130_fd_sc_hd__clkbuf_4
X_4635_ _4635_/A vssd1 vssd1 vccd1 vccd1 _6482_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4566_ _6512_/Q _4026_/A _4570_/S vssd1 vssd1 vccd1 vccd1 _4567_/A sky130_fd_sc_hd__mux2_1
X_3517_ _3517_/A vssd1 vssd1 vccd1 vccd1 _6965_/D sky130_fd_sc_hd__clkbuf_1
X_5481__320 _5483__322/A vssd1 vssd1 vccd1 vccd1 _6610_/CLK sky130_fd_sc_hd__inv_2
X_6305_ _6305_/A vssd1 vssd1 vccd1 vccd1 _6314_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4497_ _4496_/X _6543_/Q _4500_/S vssd1 vssd1 vccd1 vccd1 _4498_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__3017_ clkbuf_0__3017_/X vssd1 vssd1 vccd1 vccd1 _6133__169/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0_0__2750_ clkbuf_0__2750_/X vssd1 vssd1 vccd1 vccd1 _5577__398/A sky130_fd_sc_hd__clkbuf_4
X_6236_ _6241_/B _6241_/C _6228_/B _7004_/Q vssd1 vssd1 vccd1 vccd1 _6238_/B sky130_fd_sc_hd__a31o_1
X_3448_ _6991_/Q _3447_/X _3454_/S vssd1 vssd1 vccd1 vccd1 _3449_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6167_ _6167_/A vssd1 vssd1 vccd1 vccd1 _6167_/Y sky130_fd_sc_hd__inv_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _7026_/Q vssd1 vssd1 vccd1 vccd1 _3779_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5049_ _6377_/A _4798_/A _5046_/X _5025_/A _6430_/A vssd1 vssd1 vccd1 vccd1 _6444_/D
+ sky130_fd_sc_hd__a221oi_1
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6358__42 _6358__42/A vssd1 vssd1 vccd1 vccd1 _7062_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2879_ clkbuf_0__2879_/X vssd1 vssd1 vccd1 vccd1 _5883__79/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4420_ _3269_/X _6582_/Q _4420_/S vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__mux2_1
X_4351_ _4366_/S vssd1 vssd1 vccd1 vccd1 _4360_/S sky130_fd_sc_hd__clkbuf_2
X_5545__372 _5547__374/A vssd1 vssd1 vccd1 vccd1 _6662_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3302_ _6773_/Q vssd1 vssd1 vccd1 vccd1 _3661_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7070_ _7070_/CLK _7070_/D vssd1 vssd1 vccd1 vccd1 _7070_/Q sky130_fd_sc_hd__dfxtp_1
X_4282_ _6644_/Q _4146_/X _4288_/S vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3233_ _4693_/A _4766_/B vssd1 vssd1 vccd1 vccd1 _3241_/C sky130_fd_sc_hd__nand2_1
X_6021_ _6887_/Q _6021_/B vssd1 vssd1 vccd1 vccd1 _6021_/Y sky130_fd_sc_hd__nand2_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6923_ _6923_/CLK _6923_/D vssd1 vssd1 vccd1 vccd1 _6923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6854_ _6854_/CLK _6854_/D vssd1 vssd1 vccd1 vccd1 _6854_/Q sky130_fd_sc_hd__dfxtp_1
X_3997_ _3690_/X _6764_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _3998_/A sky130_fd_sc_hd__mux2_1
X_6785_ _6785_/CLK _6785_/D vssd1 vssd1 vccd1 vccd1 _6785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__2517_ clkbuf_0__2517_/X vssd1 vssd1 vccd1 vccd1 _5162__224/A sky130_fd_sc_hd__clkbuf_4
X_5736_ _6427_/A _5736_/B vssd1 vssd1 vccd1 vccd1 _5737_/D sky130_fd_sc_hd__and2_1
XFILLER_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5667_ _7007_/Q _5902_/B vssd1 vssd1 vccd1 vccd1 _5667_/Y sky130_fd_sc_hd__nand2_1
X_4618_ _3859_/X _6489_/Q _4618_/S vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__mux2_1
X_5598_ _5756_/A vssd1 vssd1 vccd1 vccd1 _5598_/X sky130_fd_sc_hd__buf_1
XFILLER_116_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4549_ _4549_/A vssd1 vssd1 vccd1 vccd1 _6521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2733_ clkbuf_0__2733_/X vssd1 vssd1 vccd1 vccd1 _5491__329/A sky130_fd_sc_hd__clkbuf_4
X_5446__292 _5447__293/A vssd1 vssd1 vccd1 vccd1 _6582_/CLK sky130_fd_sc_hd__inv_2
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6219_ _6229_/C vssd1 vssd1 vccd1 vccd1 _6267_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_10 _4155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_43 _4490_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_32 _3859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_21 _6705_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5488__326 _5488__326/A vssd1 vssd1 vccd1 vccd1 _6616_/CLK sky130_fd_sc_hd__inv_2
X_5681__416 _5684__419/A vssd1 vssd1 vccd1 vccd1 _6710_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5837__522 _5839__524/A vssd1 vssd1 vccd1 vccd1 _6828_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _6786_/Q _3877_/X _3926_/S vssd1 vssd1 vccd1 vccd1 _3921_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3851_ _6810_/Q _3850_/X _3860_/S vssd1 vssd1 vccd1 vccd1 _3852_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3782_ _3782_/A vssd1 vssd1 vccd1 vccd1 _3782_/X sky130_fd_sc_hd__clkbuf_2
X_6570_ _6570_/CLK _6570_/D vssd1 vssd1 vccd1 vccd1 _6570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6352__37 _6352__37/A vssd1 vssd1 vccd1 vccd1 _7057_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4403_ _4403_/A vssd1 vssd1 vccd1 vccd1 _6590_/D sky130_fd_sc_hd__clkbuf_1
X_5383_ _5289_/X _5382_/X _5292_/X vssd1 vssd1 vccd1 vccd1 _5383_/Y sky130_fd_sc_hd__o21ai_1
X_7122_ _7122_/A vssd1 vssd1 vccd1 vccd1 _7122_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4334_ _3764_/X _6621_/Q _4342_/S vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7053_ _7053_/CLK _7053_/D vssd1 vssd1 vccd1 vccd1 _7053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6004_ _6883_/Q _6882_/Q _6004_/C vssd1 vssd1 vccd1 vccd1 _6012_/B sky130_fd_sc_hd__and3_1
X_4265_ _6651_/Q _4149_/X _4269_/S vssd1 vssd1 vccd1 vccd1 _4266_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4196_ _6681_/Q _4155_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4197_/A sky130_fd_sc_hd__mux2_1
X_3216_ _6736_/Q _6735_/Q vssd1 vssd1 vccd1 vccd1 _3226_/A sky130_fd_sc_hd__nand2_1
X_5222__272 _5224__274/A vssd1 vssd1 vccd1 vccd1 _6554_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ _6906_/CLK _6906_/D vssd1 vssd1 vccd1 vccd1 _6906_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3001_ clkbuf_0__3001_/X vssd1 vssd1 vccd1 vccd1 _6049__101/A sky130_fd_sc_hd__clkbuf_4
X_6837_ _6837_/CLK _6837_/D vssd1 vssd1 vccd1 vccd1 _6837_/Q sky130_fd_sc_hd__dfxtp_1
X_6768_ _6768_/CLK _6768_/D vssd1 vssd1 vccd1 vccd1 _6768_/Q sky130_fd_sc_hd__dfxtp_2
X_5719_ _7015_/Q _5723_/B vssd1 vssd1 vccd1 vccd1 _5720_/A sky130_fd_sc_hd__and2_1
X_6699_ _6699_/CLK _6699_/D vssd1 vssd1 vccd1 vccd1 _6699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5123__192 _5123__192/A vssd1 vssd1 vccd1 vccd1 _6474_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5165__226 _5166__227/A vssd1 vssd1 vccd1 vccd1 _6508_/CLK sky130_fd_sc_hd__inv_2
XFILLER_110_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4050_ _4050_/A vssd1 vssd1 vccd1 vccd1 _6736_/D sky130_fd_sc_hd__clkbuf_1
Xinput6 caravel_wb_data_i[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
XFILLER_83_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _6485_/Q _6557_/Q _7046_/Q _6977_/Q _4923_/X _4914_/X vssd1 vssd1 vccd1 vccd1
+ _4952_/X sky130_fd_sc_hd__mux4_1
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2750_ _5573_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2750_/X sky130_fd_sc_hd__clkbuf_16
X_4883_ _5043_/B _4883_/B vssd1 vssd1 vccd1 vccd1 _4883_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3903_ _3903_/A vssd1 vssd1 vccd1 vccd1 _6794_/D sky130_fd_sc_hd__clkbuf_1
X_6622_ _6622_/CLK _6622_/D vssd1 vssd1 vccd1 vccd1 _6622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3834_ _3834_/A vssd1 vssd1 vccd1 vccd1 _6817_/D sky130_fd_sc_hd__clkbuf_1
X_6553_ _6553_/CLK _6553_/D vssd1 vssd1 vccd1 vccd1 _6553_/Q sky130_fd_sc_hd__dfxtp_1
X_3765_ _4277_/A _4277_/B _4044_/A vssd1 vssd1 vccd1 vccd1 _4404_/B sky130_fd_sc_hd__nand3_2
X_3696_ _4023_/A vssd1 vssd1 vccd1 vccd1 _3696_/X sky130_fd_sc_hd__clkbuf_4
X_6484_ _6484_/CLK _6484_/D vssd1 vssd1 vccd1 vccd1 _6484_/Q sky130_fd_sc_hd__dfxtp_1
X_6325__15 _6328__18/A vssd1 vssd1 vccd1 vccd1 _7035_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5435_ _5434_/X _5435_/B vssd1 vssd1 vccd1 vccd1 _5435_/X sky130_fd_sc_hd__and2b_1
XFILLER_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5366_ _5366_/A _5366_/B vssd1 vssd1 vccd1 vccd1 _5366_/Y sky130_fd_sc_hd__nand2_1
X_7105_ _7105_/A vssd1 vssd1 vccd1 vccd1 _7105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4317_ _4317_/A vssd1 vssd1 vccd1 vccd1 _6629_/D sky130_fd_sc_hd__clkbuf_1
X_5297_ _6013_/A vssd1 vssd1 vccd1 vccd1 _6019_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7036_ _7036_/CLK _7036_/D vssd1 vssd1 vccd1 vccd1 _7036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4248_ _4248_/A vssd1 vssd1 vccd1 vccd1 _6659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6375__3 _6376__4/A vssd1 vssd1 vccd1 vccd1 _7077_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4179_ _4179_/A vssd1 vssd1 vccd1 vccd1 _6689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2879_ _5878_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2879_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5229__278 _5229__278/A vssd1 vssd1 vccd1 vccd1 _6560_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3550_ _3550_/A vssd1 vssd1 vccd1 vccd1 _6951_/D sky130_fd_sc_hd__clkbuf_1
X_3481_ _3481_/A vssd1 vssd1 vccd1 vccd1 _6979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5151_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__buf_1
XFILLER_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4102_ _4102_/A vssd1 vssd1 vccd1 vccd1 _6723_/D sky130_fd_sc_hd__clkbuf_1
X_5082_ _6458_/Q _7112_/A _5082_/S vssd1 vssd1 vccd1 vccd1 _5083_/A sky130_fd_sc_hd__mux2_1
X_4033_ _4032_/X _6751_/Q _4033_/S vssd1 vssd1 vccd1 vccd1 _4034_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__2834_ clkbuf_0__2834_/X vssd1 vssd1 vccd1 vccd1 _5694__427/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5984_ _6879_/Q _5985_/B vssd1 vssd1 vccd1 vccd1 _5994_/C sky130_fd_sc_hd__and2_1
X_4935_ _3986_/X _6516_/Q _4934_/X _4806_/X vssd1 vssd1 vccd1 vccd1 _4935_/X sky130_fd_sc_hd__o211a_1
X_4866_ _6763_/Q _6755_/Q _6718_/Q _6710_/Q _4957_/S _4914_/A vssd1 vssd1 vccd1 vccd1
+ _4866_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_0__2733_ _5486_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2733_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4797_ _3971_/X _4793_/X _4918_/A vssd1 vssd1 vccd1 vccd1 _4797_/Y sky130_fd_sc_hd__a21oi_1
X_3817_ _6824_/Q _3608_/X _3819_/S vssd1 vssd1 vccd1 vccd1 _3818_/A sky130_fd_sc_hd__mux2_1
X_6605_ _6605_/CLK _6605_/D vssd1 vssd1 vccd1 vccd1 _6605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6536_ _6536_/CLK _6536_/D vssd1 vssd1 vccd1 vccd1 _6536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3748_ _6851_/Q _3597_/X _3756_/S vssd1 vssd1 vccd1 vccd1 _3749_/A sky130_fd_sc_hd__mux2_1
X_6467_ _7019_/CLK _6467_/D vssd1 vssd1 vccd1 vccd1 _6467_/Q sky130_fd_sc_hd__dfxtp_1
X_3679_ _3679_/A vssd1 vssd1 vccd1 vccd1 _6898_/D sky130_fd_sc_hd__clkbuf_1
Xoutput151 _7147_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput140 _7137_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[12] sky130_fd_sc_hd__buf_2
X_6398_ _7136_/A _5892_/A _6401_/S vssd1 vssd1 vccd1 vccd1 _6399_/B sky130_fd_sc_hd__mux2_1
X_5418_ _5437_/A _5418_/B vssd1 vssd1 vccd1 vccd1 _5418_/Y sky130_fd_sc_hd__nor2_1
Xoutput173 _4687_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_stb_o sky130_fd_sc_hd__buf_2
Xoutput162 _7128_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput195 _5011_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput184 _4989_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5349_ _6576_/Q _5250_/X _5348_/X _5298_/X vssd1 vssd1 vccd1 vccd1 _6576_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7019_ _7019_/CLK _7019_/D vssd1 vssd1 vccd1 vccd1 _7019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _6852_/Q _6828_/Q _6804_/Q _6796_/Q _4891_/B _4719_/X vssd1 vssd1 vccd1 vccd1
+ _4720_/X sky130_fd_sc_hd__mux4_2
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4651_ _4651_/A vssd1 vssd1 vccd1 vccd1 _6475_/D sky130_fd_sc_hd__clkbuf_1
Xinput20 caravel_wb_data_i[25] vssd1 vssd1 vccd1 vccd1 _5006_/B sky130_fd_sc_hd__buf_4
Xinput31 caravel_wb_data_i[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_2
X_3602_ _7029_/Q vssd1 vssd1 vccd1 vccd1 _3602_/X sky130_fd_sc_hd__buf_6
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4582_ _4490_/X _6505_/Q _4582_/S vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__mux2_1
Xinput42 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 _7112_/A sky130_fd_sc_hd__buf_4
Xinput53 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 _7122_/A sky130_fd_sc_hd__buf_4
Xinput64 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 _7103_/A sky130_fd_sc_hd__buf_4
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3533_ _3533_/A vssd1 vssd1 vccd1 vccd1 _6958_/D sky130_fd_sc_hd__clkbuf_1
Xinput97 wbs_data_i[6] vssd1 vssd1 vccd1 vccd1 _7131_/A sky130_fd_sc_hd__clkbuf_8
Xinput75 wbs_data_i[15] vssd1 vssd1 vccd1 vccd1 _7140_/A sky130_fd_sc_hd__buf_4
Xinput86 wbs_data_i[25] vssd1 vssd1 vccd1 vccd1 _7150_/A sky130_fd_sc_hd__buf_4
X_5509__343 _5510__344/A vssd1 vssd1 vccd1 vccd1 _6633_/CLK sky130_fd_sc_hd__inv_2
X_6252_ _6249_/X _6267_/A _6252_/C vssd1 vssd1 vccd1 vccd1 _6253_/A sky130_fd_sc_hd__and3b_1
X_3464_ _3464_/A vssd1 vssd1 vccd1 vccd1 _6986_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6183_ _6245_/A _6272_/A input1/X vssd1 vssd1 vccd1 vccd1 _6184_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_0__3001_ _6047_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3001_/X sky130_fd_sc_hd__clkbuf_16
X_3395_ _7127_/A _3242_/A _5047_/A vssd1 vssd1 vccd1 vccd1 _3947_/A sky130_fd_sc_hd__a21oi_4
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5065_ _6450_/Q _7104_/A _5071_/S vssd1 vssd1 vccd1 vccd1 _5066_/A sky130_fd_sc_hd__mux2_1
X_4016_ _4016_/A vssd1 vssd1 vccd1 vccd1 _6757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5178__236 _5181__239/A vssd1 vssd1 vccd1 vccd1 _6518_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5967_ _6876_/Q _5968_/B vssd1 vssd1 vccd1 vccd1 _5969_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1_0__2748_ clkbuf_0__2748_/X vssd1 vssd1 vccd1 vccd1 _5564__387/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4918_ _4918_/A _4918_/B vssd1 vssd1 vccd1 vccd1 _4918_/Y sky130_fd_sc_hd__nor2_1
X_5898_ _6880_/Q _5898_/B _5898_/C vssd1 vssd1 vccd1 vccd1 _5898_/X sky130_fd_sc_hd__and3_1
XFILLER_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4849_ _4876_/A _6625_/Q vssd1 vssd1 vccd1 vccd1 _4849_/X sky130_fd_sc_hd__or2_1
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6519_ _6519_/CLK _6519_/D vssd1 vssd1 vccd1 vccd1 _6519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5831__517 _5831__517/A vssd1 vssd1 vccd1 vccd1 _6823_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6151__8 _6152__9/A vssd1 vssd1 vccd1 vccd1 _6991_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6870_ _7095_/CLK _6870_/D vssd1 vssd1 vccd1 vccd1 _6870_/Q sky130_fd_sc_hd__dfxtp_1
X_5821_ _5821_/A vssd1 vssd1 vccd1 vccd1 _5821_/X sky130_fd_sc_hd__buf_1
XFILLER_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0__2533_ clkbuf_0__2533_/X vssd1 vssd1 vccd1 vccd1 _5449_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4703_ _4954_/S _4703_/B vssd1 vssd1 vccd1 vccd1 _4703_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4634_ _3856_/X _6482_/Q _4636_/S vssd1 vssd1 vccd1 vccd1 _4635_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4565_ _4565_/A vssd1 vssd1 vccd1 vccd1 _6513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3516_ _6965_/Q _3453_/X _3516_/S vssd1 vssd1 vccd1 vccd1 _3517_/A sky130_fd_sc_hd__mux2_1
X_6304_ _6304_/A vssd1 vssd1 vccd1 vccd1 _7023_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4496_ _6742_/Q vssd1 vssd1 vccd1 vccd1 _4496_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0__3016_ clkbuf_0__3016_/X vssd1 vssd1 vccd1 vccd1 _6127__164/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6235_ _6235_/A vssd1 vssd1 vccd1 vccd1 _7003_/D sky130_fd_sc_hd__clkbuf_1
X_3447_ _3773_/A vssd1 vssd1 vccd1 vccd1 _3447_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6166_ _7010_/Q vssd1 vssd1 vccd1 vccd1 _6166_/Y sky130_fd_sc_hd__inv_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _3378_/A vssd1 vssd1 vccd1 vccd1 _7051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5117_/A vssd1 vssd1 vccd1 vccd1 _6469_/D sky130_fd_sc_hd__clkbuf_1
X_6097_ _6097_/A vssd1 vssd1 vccd1 vccd1 _6097_/X sky130_fd_sc_hd__buf_1
X_5048_ _6433_/A vssd1 vssd1 vccd1 vccd1 _6430_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6999_ _7093_/CLK _6999_/D vssd1 vssd1 vccd1 vccd1 _6999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5787__482 _5789__484/A vssd1 vssd1 vccd1 vccd1 _6788_/CLK sky130_fd_sc_hd__inv_2
X_5709__439 _5709__439/A vssd1 vssd1 vccd1 vccd1 _6733_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2878_ clkbuf_0__2878_/X vssd1 vssd1 vccd1 vccd1 _5877__74/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5755__459 _5755__459/A vssd1 vssd1 vccd1 vccd1 _6763_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4350_ _4350_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4366_/S sky130_fd_sc_hd__nor2_2
X_3301_ _3990_/C _3990_/B _3727_/B vssd1 vssd1 vccd1 vccd1 _4644_/A sky130_fd_sc_hd__nand3_4
XFILLER_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4281_ _4281_/A vssd1 vssd1 vccd1 vccd1 _6645_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3232_ _6447_/Q _6448_/Q _4741_/B vssd1 vssd1 vccd1 vccd1 _4766_/B sky130_fd_sc_hd__or3_1
X_6020_ _6020_/A vssd1 vssd1 vccd1 vccd1 _6886_/D sky130_fd_sc_hd__clkbuf_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6922_ _6922_/CLK _6922_/D vssd1 vssd1 vccd1 vccd1 _6922_/Q sky130_fd_sc_hd__dfxtp_1
X_6853_ _6853_/CLK _6853_/D vssd1 vssd1 vccd1 vccd1 _6853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6082__128 _6082__128/A vssd1 vssd1 vccd1 vccd1 _6936_/CLK sky130_fd_sc_hd__inv_2
X_3996_ _3996_/A vssd1 vssd1 vccd1 vccd1 _6765_/D sky130_fd_sc_hd__clkbuf_1
X_6784_ _6784_/CLK _6784_/D vssd1 vssd1 vccd1 vccd1 _6784_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__2516_ clkbuf_0__2516_/X vssd1 vssd1 vccd1 vccd1 _5155__218/A sky130_fd_sc_hd__clkbuf_4
X_5735_ _5735_/A vssd1 vssd1 vccd1 vccd1 _6748_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5666_ _7007_/Q _5902_/B vssd1 vssd1 vccd1 vccd1 _5666_/X sky130_fd_sc_hd__or2_1
XFILLER_108_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4617_ _4617_/A vssd1 vssd1 vccd1 vccd1 _6490_/D sky130_fd_sc_hd__clkbuf_1
X_5597_ _5597_/A vssd1 vssd1 vccd1 vccd1 _5597_/X sky130_fd_sc_hd__buf_1
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4548_ _4490_/X _6521_/Q _4548_/S vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__mux2_1
X_4479_ _4476_/X _6549_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2732_ clkbuf_0__2732_/X vssd1 vssd1 vccd1 vccd1 _5483__322/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6218_ _6249_/C _6250_/C vssd1 vssd1 vccd1 vccd1 _6224_/B sky130_fd_sc_hd__and2_1
XFILLER_100_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_33 _3859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_22 _7136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_11 _4164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_44 _4701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5761__463 _5762__464/A vssd1 vssd1 vccd1 vccd1 _6767_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3850_ _6747_/Q vssd1 vssd1 vccd1 vccd1 _3850_/X sky130_fd_sc_hd__buf_6
X_3781_ _3781_/A vssd1 vssd1 vccd1 vccd1 _6839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5382_ _6958_/Q _6942_/Q _7067_/Q _6934_/Q _5266_/X _5268_/X vssd1 vssd1 vccd1 vccd1
+ _5382_/X sky130_fd_sc_hd__mux4_2
X_4402_ _3269_/X _6590_/Q _4402_/S vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__mux2_1
X_7121_ _7121_/A vssd1 vssd1 vccd1 vccd1 _7121_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4333_ _4348_/S vssd1 vssd1 vccd1 vccd1 _4342_/S sky130_fd_sc_hd__buf_2
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7052_ _7052_/CLK _7052_/D vssd1 vssd1 vccd1 vccd1 _7052_/Q sky130_fd_sc_hd__dfxtp_1
X_4264_ _4264_/A vssd1 vssd1 vccd1 vccd1 _6652_/D sky130_fd_sc_hd__clkbuf_1
X_3215_ _4048_/A _5258_/A _4068_/A _3214_/X vssd1 vssd1 vccd1 vccd1 _3227_/A sky130_fd_sc_hd__a211oi_1
X_6003_ _6003_/A vssd1 vssd1 vccd1 vccd1 _6882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4195_ _4195_/A vssd1 vssd1 vccd1 vccd1 _6682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6905_ _6905_/CLK _6905_/D vssd1 vssd1 vccd1 vccd1 _6905_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3000_ clkbuf_0__3000_/X vssd1 vssd1 vccd1 vccd1 _6046__99/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6836_ _6836_/CLK _6836_/D vssd1 vssd1 vccd1 vccd1 _6836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6767_ _6767_/CLK _6767_/D vssd1 vssd1 vccd1 vccd1 _6767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3979_ _3968_/A _3981_/A _3978_/Y vssd1 vssd1 vccd1 vccd1 _6769_/D sky130_fd_sc_hd__o21a_1
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6698_ _6698_/CLK _6698_/D vssd1 vssd1 vccd1 vccd1 _6698_/Q sky130_fd_sc_hd__dfxtp_1
X_5649_ _6996_/Q _5648_/A vssd1 vssd1 vccd1 vccd1 _5649_/X sky130_fd_sc_hd__or2b_1
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5494__331 _5494__331/A vssd1 vssd1 vccd1 vccd1 _6621_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5503__338 _5504__339/A vssd1 vssd1 vccd1 vccd1 _6628_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput7 caravel_wb_data_i[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_2
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _4944_/X _4946_/X _4948_/X _4950_/X _3951_/Y vssd1 vssd1 vccd1 vccd1 _4951_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4882_ _4802_/X _4875_/X _4881_/X _4724_/A vssd1 vssd1 vccd1 vccd1 _4882_/X sky130_fd_sc_hd__a211o_1
X_3902_ _6794_/Q _3602_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6621_ _6621_/CLK _6621_/D vssd1 vssd1 vccd1 vccd1 _6621_/Q sky130_fd_sc_hd__dfxtp_1
X_3833_ _6817_/Q _3605_/X _3837_/S vssd1 vssd1 vccd1 vccd1 _3834_/A sky130_fd_sc_hd__mux2_1
X_5768__469 _5768__469/A vssd1 vssd1 vccd1 vccd1 _6773_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6552_ _6552_/CLK _6552_/D vssd1 vssd1 vccd1 vccd1 _6552_/Q sky130_fd_sc_hd__dfxtp_1
X_3764_ _3764_/A vssd1 vssd1 vccd1 vccd1 _3764_/X sky130_fd_sc_hd__clkbuf_2
X_3695_ _3695_/A vssd1 vssd1 vccd1 vccd1 _6893_/D sky130_fd_sc_hd__clkbuf_1
X_6483_ _6483_/CLK _6483_/D vssd1 vssd1 vccd1 vccd1 _6483_/Q sky130_fd_sc_hd__dfxtp_1
X_5434_ _6795_/Q _6985_/Q _6993_/Q _6969_/Q _5341_/A _5251_/X vssd1 vssd1 vccd1 vccd1
+ _5434_/X sky130_fd_sc_hd__mux4_2
X_7104_ _7104_/A vssd1 vssd1 vccd1 vccd1 _7104_/X sky130_fd_sc_hd__clkbuf_1
X_5365_ _5361_/X _5364_/X _5433_/S vssd1 vssd1 vccd1 vccd1 _5366_/B sky130_fd_sc_hd__mux2_1
X_4316_ _6629_/Q _3871_/X _4324_/S vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__mux2_1
X_5296_ _4055_/X _5273_/X _5295_/Y vssd1 vssd1 vccd1 vccd1 _5296_/X sky130_fd_sc_hd__a21o_1
X_7035_ _7035_/CLK _7035_/D vssd1 vssd1 vccd1 vccd1 _7035_/Q sky130_fd_sc_hd__dfxtp_1
X_4247_ _3773_/X _6659_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4248_/A sky130_fd_sc_hd__mux2_1
X_4178_ _4023_/X _6689_/Q _4178_/S vssd1 vssd1 vccd1 vccd1 _4179_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5558__383 _5559__384/A vssd1 vssd1 vccd1 vccd1 _6673_/CLK sky130_fd_sc_hd__inv_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_6819_ _6819_/CLK _6819_/D vssd1 vssd1 vccd1 vccd1 _6819_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2878_ _5872_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2878_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6095__138 _6096__139/A vssd1 vssd1 vccd1 vccd1 _6946_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5171__231 _5174__234/A vssd1 vssd1 vccd1 vccd1 _6513_/CLK sky130_fd_sc_hd__inv_2
X_3480_ _3388_/X _6979_/Q _3482_/S vssd1 vssd1 vccd1 vccd1 _3481_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4101_ _4029_/X _6723_/Q _4103_/S vssd1 vssd1 vccd1 vccd1 _4102_/A sky130_fd_sc_hd__mux2_1
X_5694__427 _5694__427/A vssd1 vssd1 vccd1 vccd1 _6721_/CLK sky130_fd_sc_hd__inv_2
XFILLER_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5081_ _5081_/A vssd1 vssd1 vccd1 vccd1 _6457_/D sky130_fd_sc_hd__clkbuf_1
X_4032_ _4032_/A vssd1 vssd1 vccd1 vccd1 _4032_/X sky130_fd_sc_hd__buf_4
XFILLER_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2833_ clkbuf_0__2833_/X vssd1 vssd1 vccd1 vccd1 _5690__424/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5983_ _5983_/A vssd1 vssd1 vccd1 vccd1 _6878_/D sky130_fd_sc_hd__clkbuf_1
X_4934_ _4956_/S _6500_/Q vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__or2_1
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4865_ _4865_/A _4865_/B vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__or2_1
Xclkbuf_0__2732_ _5480_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2732_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4796_ _4856_/A _5776_/B vssd1 vssd1 vccd1 vccd1 _4918_/A sky130_fd_sc_hd__or2_1
X_3816_ _3816_/A vssd1 vssd1 vccd1 vccd1 _6825_/D sky130_fd_sc_hd__clkbuf_1
X_6604_ _6604_/CLK _6604_/D vssd1 vssd1 vccd1 vccd1 _6604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6535_ _6535_/CLK _6535_/D vssd1 vssd1 vccd1 vccd1 _6535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3747_ _3762_/S vssd1 vssd1 vccd1 vccd1 _3756_/S sky130_fd_sc_hd__clkbuf_2
X_5781__477 _5783__479/A vssd1 vssd1 vccd1 vccd1 _6783_/CLK sky130_fd_sc_hd__inv_2
XFILLER_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3678_ _3353_/X _6898_/Q _3678_/S vssd1 vssd1 vccd1 vccd1 _3679_/A sky130_fd_sc_hd__mux2_1
X_6466_ _6897_/CLK _6466_/D vssd1 vssd1 vccd1 vccd1 _6466_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput152 _7148_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput130 _7101_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[4] sky130_fd_sc_hd__buf_2
Xoutput141 _7138_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[13] sky130_fd_sc_hd__buf_2
X_6397_ _6397_/A vssd1 vssd1 vccd1 vccd1 _7084_/D sky130_fd_sc_hd__clkbuf_1
X_5417_ _6952_/Q _6684_/Q _6596_/Q _6818_/Q _5337_/X _5338_/X vssd1 vssd1 vccd1 vccd1
+ _5418_/B sky130_fd_sc_hd__mux4_2
Xoutput163 _7129_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[4] sky130_fd_sc_hd__buf_2
Xoutput174 _7161_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_we_o sky130_fd_sc_hd__buf_2
XFILLER_102_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput185 _4991_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5348_ _5324_/X _5333_/X _5347_/Y vssd1 vssd1 vccd1 vccd1 _5348_/X sky130_fd_sc_hd__a21o_1
XFILLER_101_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput196 _5013_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[28] sky130_fd_sc_hd__buf_2
X_7018_ _7022_/CLK _7018_/D vssd1 vssd1 vccd1 vccd1 _7018_/Q sky130_fd_sc_hd__dfxtp_1
X_5279_ _5277_/X _5364_/S vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__and2b_1
XFILLER_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5235__283 _5235__283/A vssd1 vssd1 vccd1 vccd1 _6565_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5242__287 _5242__287/A vssd1 vssd1 vccd1 vccd1 _6569_/CLK sky130_fd_sc_hd__inv_2
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ _3853_/X _6475_/Q _4654_/S vssd1 vssd1 vccd1 vccd1 _4651_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput21 caravel_wb_data_i[26] vssd1 vssd1 vccd1 vccd1 _5008_/B sky130_fd_sc_hd__buf_4
Xinput10 caravel_wb_data_i[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_2
X_3601_ _3601_/A vssd1 vssd1 vccd1 vccd1 _6929_/D sky130_fd_sc_hd__clkbuf_1
Xinput32 caravel_wb_data_i[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_2
X_4581_ _4581_/A vssd1 vssd1 vccd1 vccd1 _6506_/D sky130_fd_sc_hd__clkbuf_1
Xinput43 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 _7113_/A sky130_fd_sc_hd__buf_4
Xinput54 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 _7123_/A sky130_fd_sc_hd__buf_4
X_3532_ _6958_/Q _3450_/X _3534_/S vssd1 vssd1 vccd1 vccd1 _3533_/A sky130_fd_sc_hd__mux2_1
Xinput65 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 _7104_/A sky130_fd_sc_hd__buf_4
Xinput98 wbs_data_i[7] vssd1 vssd1 vccd1 vccd1 _7132_/A sky130_fd_sc_hd__buf_6
Xinput76 wbs_data_i[16] vssd1 vssd1 vccd1 vccd1 _7141_/A sky130_fd_sc_hd__buf_4
Xinput87 wbs_data_i[26] vssd1 vssd1 vccd1 vccd1 _7151_/A sky130_fd_sc_hd__buf_4
XFILLER_107_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6251_ _6249_/C _6254_/D _7006_/Q vssd1 vssd1 vccd1 vccd1 _6252_/C sky130_fd_sc_hd__a21o_1
X_3463_ _6986_/Q _3462_/X _3463_/S vssd1 vssd1 vccd1 vccd1 _3464_/A sky130_fd_sc_hd__mux2_1
X_5702__434 _5702__434/A vssd1 vssd1 vccd1 vccd1 _6728_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6182_ _6994_/Q vssd1 vssd1 vccd1 vccd1 _6272_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3000_ _6041_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3000_/X sky130_fd_sc_hd__clkbuf_16
X_3394_ _3394_/A vssd1 vssd1 vccd1 vccd1 _7047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5064_ _5064_/A vssd1 vssd1 vccd1 vccd1 _6449_/D sky130_fd_sc_hd__clkbuf_1
X_4015_ _4014_/X _6757_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__2747_ clkbuf_0__2747_/X vssd1 vssd1 vccd1 vccd1 _5591_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5966_ _5966_/A vssd1 vssd1 vccd1 vccd1 _5966_/X sky130_fd_sc_hd__clkbuf_2
X_4917_ _4908_/Y _4911_/Y _4913_/Y _4916_/Y _4904_/A vssd1 vssd1 vccd1 vccd1 _4918_/B
+ sky130_fd_sc_hd__o221a_2
X_5897_ _6882_/Q _5897_/B vssd1 vssd1 vccd1 vccd1 _5897_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4848_ _4846_/X _4847_/X _4875_/S vssd1 vssd1 vccd1 vccd1 _4848_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4779_ _6890_/Q _6519_/Q _6495_/Q _6511_/Q _4778_/X _3959_/A vssd1 vssd1 vccd1 vccd1
+ _4779_/X sky130_fd_sc_hd__mux4_1
XFILLER_107_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6518_ _6518_/CLK _6518_/D vssd1 vssd1 vccd1 vccd1 _6518_/Q sky130_fd_sc_hd__dfxtp_1
X_6449_ _6750_/CLK _6449_/D vssd1 vssd1 vccd1 vccd1 _6449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4702_ _6470_/Q _6622_/Q _7055_/Q _6780_/Q _4914_/A _4701_/X vssd1 vssd1 vccd1 vccd1
+ _4703_/B sky130_fd_sc_hd__mux4_1
XFILLER_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _4633_/A vssd1 vssd1 vccd1 vccd1 _6483_/D sky130_fd_sc_hd__clkbuf_1
X_4564_ _6513_/Q _4023_/A _4570_/S vssd1 vssd1 vccd1 vccd1 _4565_/A sky130_fd_sc_hd__mux2_1
X_6303_ _7125_/A _6303_/B _6312_/C vssd1 vssd1 vccd1 vccd1 _6304_/A sky130_fd_sc_hd__and3_1
X_3515_ _3515_/A vssd1 vssd1 vccd1 vccd1 _6966_/D sky130_fd_sc_hd__clkbuf_1
X_4495_ _4495_/A vssd1 vssd1 vccd1 vccd1 _6544_/D sky130_fd_sc_hd__clkbuf_1
X_6234_ _6238_/A _6234_/B _6234_/C vssd1 vssd1 vccd1 vccd1 _6235_/A sky130_fd_sc_hd__and3_1
Xclkbuf_1_1_0__3015_ clkbuf_0__3015_/X vssd1 vssd1 vccd1 vccd1 _6119__157/A sky130_fd_sc_hd__clkbuf_4
X_5184__241 _5186__243/A vssd1 vssd1 vccd1 vccd1 _6523_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3446_ _3446_/A vssd1 vssd1 vccd1 vccd1 _6992_/D sky130_fd_sc_hd__clkbuf_1
X_6165_ _6161_/Y _6266_/A _6162_/Y _4974_/X _6164_/X vssd1 vssd1 vccd1 vccd1 _6172_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _3376_/X _7051_/Q _3381_/S vssd1 vssd1 vccd1 vccd1 _3378_/A sky130_fd_sc_hd__mux2_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _7161_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5117_/A sky130_fd_sc_hd__and2b_1
X_5047_ _5047_/A vssd1 vssd1 vccd1 vccd1 _6433_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6998_ _7093_/CLK _6998_/D vssd1 vssd1 vccd1 vccd1 _6998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5949_ _5972_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5950_/A sky130_fd_sc_hd__and2_1
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2877_ clkbuf_0__2877_/X vssd1 vssd1 vccd1 vccd1 _5870__68/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5458__302 _5458__302/A vssd1 vssd1 vccd1 vccd1 _6592_/CLK sky130_fd_sc_hd__inv_2
X_5794__487 _5795__488/A vssd1 vssd1 vccd1 vccd1 _6793_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6364__47 _6366__49/A vssd1 vssd1 vccd1 vccd1 _7067_/CLK sky130_fd_sc_hd__inv_2
X_3300_ _4167_/B vssd1 vssd1 vccd1 vccd1 _3727_/B sky130_fd_sc_hd__clkbuf_4
X_4280_ _6645_/Q _4141_/X _4288_/S vssd1 vssd1 vccd1 vccd1 _4281_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3231_ _6449_/Q _6450_/Q _6451_/Q _6452_/Q vssd1 vssd1 vccd1 vccd1 _4741_/B sky130_fd_sc_hd__or4_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6921_ _6921_/CLK _6921_/D vssd1 vssd1 vccd1 vccd1 _6921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6852_ _6852_/CLK _6852_/D vssd1 vssd1 vccd1 vccd1 _6852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5803_ _5809_/A vssd1 vssd1 vccd1 vccd1 _5803_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__2515_ clkbuf_0__2515_/X vssd1 vssd1 vccd1 vccd1 _5150__214/A sky130_fd_sc_hd__clkbuf_4
X_3995_ _3687_/X _6765_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__mux2_1
X_6783_ _6783_/CLK _6783_/D vssd1 vssd1 vccd1 vccd1 _6783_/Q sky130_fd_sc_hd__dfxtp_1
X_5552__378 _5553__379/A vssd1 vssd1 vccd1 vccd1 _6668_/CLK sky130_fd_sc_hd__inv_2
X_5734_ _7022_/Q _5734_/B vssd1 vssd1 vccd1 vccd1 _5735_/A sky130_fd_sc_hd__and2_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5665_ _4978_/X _5898_/B _5659_/B vssd1 vssd1 vccd1 vccd1 _5902_/B sky130_fd_sc_hd__a21boi_2
X_4616_ _3856_/X _6490_/Q _4618_/S vssd1 vssd1 vccd1 vccd1 _4617_/A sky130_fd_sc_hd__mux2_1
X_4547_ _4547_/A vssd1 vssd1 vccd1 vccd1 _6522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4478_ _4500_/S vssd1 vssd1 vccd1 vccd1 _4491_/S sky130_fd_sc_hd__buf_2
XFILLER_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2731_ clkbuf_0__2731_/X vssd1 vssd1 vccd1 vccd1 _5479__319/A sky130_fd_sc_hd__clkbuf_4
X_6217_ _7000_/Q _6217_/B _6217_/C vssd1 vssd1 vccd1 vccd1 _6250_/C sky130_fd_sc_hd__and3_1
X_3429_ _3380_/X _7034_/Q _3429_/S vssd1 vssd1 vccd1 vccd1 _3430_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_12 _4662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_34 _3859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_23 _7136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_45 _7055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5715__444 _5715__444/A vssd1 vssd1 vccd1 vccd1 _6738_/CLK sky130_fd_sc_hd__inv_2
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5453__298 _5453__298/A vssd1 vssd1 vccd1 vccd1 _6588_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6059__109 _6059__109/A vssd1 vssd1 vccd1 vccd1 _6917_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5802__494 _5802__494/A vssd1 vssd1 vccd1 vccd1 _6800_/CLK sky130_fd_sc_hd__inv_2
X_5857__57 _5857__57/A vssd1 vssd1 vccd1 vccd1 _6843_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2875_ clkbuf_0__2875_/X vssd1 vssd1 vccd1 vccd1 _5859__59/A sky130_fd_sc_hd__clkbuf_16
XFILLER_95_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5135__202 _5136__203/A vssd1 vssd1 vccd1 vccd1 _6484_/CLK sky130_fd_sc_hd__inv_2
X_3780_ _3779_/X _6839_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3781_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0__f__2454_ clkbuf_0__2454_/X vssd1 vssd1 vccd1 vccd1 _5206_/A sky130_fd_sc_hd__clkbuf_16
X_5844__528 _5845__529/A vssd1 vssd1 vccd1 vccd1 _6834_/CLK sky130_fd_sc_hd__inv_2
X_6337__25 _6338__26/A vssd1 vssd1 vccd1 vccd1 _7045_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4401_ _4401_/A vssd1 vssd1 vccd1 vccd1 _6591_/D sky130_fd_sc_hd__clkbuf_1
X_5381_ _5380_/X _5432_/S vssd1 vssd1 vccd1 vccd1 _5381_/X sky130_fd_sc_hd__and2b_1
X_7120_ _7120_/A vssd1 vssd1 vccd1 vccd1 _7120_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
X_4332_ _4404_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4348_/S sky130_fd_sc_hd__or2_2
XFILLER_113_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7051_ _7051_/CLK _7051_/D vssd1 vssd1 vccd1 vccd1 _7051_/Q sky130_fd_sc_hd__dfxtp_1
X_4263_ _6652_/Q _4146_/X _4269_/S vssd1 vssd1 vccd1 vccd1 _4264_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3214_ _5302_/A _3221_/A _3221_/B _3213_/Y _3361_/A vssd1 vssd1 vccd1 vccd1 _3214_/X
+ sky130_fd_sc_hd__o2111a_1
X_6002_ _6002_/A _6002_/B vssd1 vssd1 vccd1 vccd1 _6003_/A sky130_fd_sc_hd__and2_1
XFILLER_67_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4194_ _6682_/Q _4152_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6904_ _6904_/CLK _6904_/D vssd1 vssd1 vccd1 vccd1 _6904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6835_ _6835_/CLK _6835_/D vssd1 vssd1 vccd1 vccd1 _6835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6766_ _6766_/CLK _6766_/D vssd1 vssd1 vccd1 vccd1 _6766_/Q sky130_fd_sc_hd__dfxtp_1
X_3978_ _5776_/A _3978_/B vssd1 vssd1 vccd1 vccd1 _3978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6697_ _6697_/CLK _6697_/D vssd1 vssd1 vccd1 vccd1 _6697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _5648_/A _6216_/C vssd1 vssd1 vccd1 vccd1 _5648_/X sky130_fd_sc_hd__or2b_1
XFILLER_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5579_ _5591_/A vssd1 vssd1 vccd1 vccd1 _5579_/X sky130_fd_sc_hd__buf_1
XFILLER_116_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5130__198 _5130__198/A vssd1 vssd1 vccd1 vccd1 _6480_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 caravel_wb_data_i[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4950_ _4944_/A _4949_/X _4782_/X vssd1 vssd1 vccd1 vccd1 _4950_/X sky130_fd_sc_hd__o21a_1
XFILLER_17_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4881_ _4877_/X _4879_/X _4880_/X _4804_/A _3953_/A vssd1 vssd1 vccd1 vccd1 _4881_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3901_ _3901_/A vssd1 vssd1 vccd1 vccd1 _6795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6620_ _6620_/CLK _6620_/D vssd1 vssd1 vccd1 vccd1 _6620_/Q sky130_fd_sc_hd__dfxtp_1
X_3832_ _3832_/A vssd1 vssd1 vccd1 vccd1 _6818_/D sky130_fd_sc_hd__clkbuf_1
X_6551_ _6551_/CLK _6551_/D vssd1 vssd1 vccd1 vccd1 _6551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3763_ _3763_/A vssd1 vssd1 vccd1 vccd1 _6844_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3694_ _3693_/X _6893_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3695_/A sky130_fd_sc_hd__mux2_1
X_6482_ _6482_/CLK _6482_/D vssd1 vssd1 vccd1 vccd1 _6482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5433_ _5429_/X _5432_/X _5433_/S vssd1 vssd1 vccd1 vccd1 _5433_/X sky130_fd_sc_hd__mux2_1
X_5364_ _5362_/X _5363_/X _5364_/S vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__mux2_1
X_7103_ _7103_/A vssd1 vssd1 vccd1 vccd1 _7103_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4315_ _4330_/S vssd1 vssd1 vccd1 vccd1 _4324_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5295_ _5366_/A _5294_/X _5250_/A vssd1 vssd1 vccd1 vccd1 _5295_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4246_ _4246_/A vssd1 vssd1 vccd1 vccd1 _6660_/D sky130_fd_sc_hd__clkbuf_1
X_7034_ _7034_/CLK _7034_/D vssd1 vssd1 vccd1 vccd1 _7034_/Q sky130_fd_sc_hd__dfxtp_1
X_4177_ _4177_/A vssd1 vssd1 vccd1 vccd1 _6690_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6129__165 _6132__168/A vssd1 vssd1 vccd1 vccd1 _6973_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6818_ _6818_/CLK _6818_/D vssd1 vssd1 vccd1 vccd1 _6818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__2877_ _5866_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2877_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6749_ _7096_/CLK _6749_/D vssd1 vssd1 vccd1 vccd1 _6749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5565__388 _5566__389/A vssd1 vssd1 vccd1 vccd1 _6678_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4100_ _4100_/A vssd1 vssd1 vccd1 vccd1 _6724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5080_ _6457_/Q _7111_/A _5082_/S vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__mux2_1
X_4031_ _4031_/A vssd1 vssd1 vccd1 vccd1 _6752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__2832_ clkbuf_0__2832_/X vssd1 vssd1 vccd1 vccd1 _5684__419/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5590__404 _5590__404/A vssd1 vssd1 vccd1 vccd1 _6697_/CLK sky130_fd_sc_hd__inv_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5982_ _6002_/A _5982_/B vssd1 vssd1 vccd1 vccd1 _5983_/A sky130_fd_sc_hd__and2_1
X_4933_ _4931_/X _4932_/X _4933_/S vssd1 vssd1 vccd1 vccd1 _4933_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2731_ _5474_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2731_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_33_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4864_ _6856_/Q _6832_/Q _6808_/Q _6800_/Q _4814_/A _4845_/X vssd1 vssd1 vccd1 vccd1
+ _4865_/B sky130_fd_sc_hd__mux4_2
X_4795_ _4795_/A _4795_/B _4794_/X vssd1 vssd1 vccd1 vccd1 _5776_/B sky130_fd_sc_hd__or3b_1
X_3815_ _6825_/Q _3605_/X _3819_/S vssd1 vssd1 vccd1 vccd1 _3816_/A sky130_fd_sc_hd__mux2_1
X_6603_ _6603_/CLK _6603_/D vssd1 vssd1 vccd1 vccd1 _6603_/Q sky130_fd_sc_hd__dfxtp_1
X_6534_ _6534_/CLK _6534_/D vssd1 vssd1 vccd1 vccd1 _6534_/Q sky130_fd_sc_hd__dfxtp_1
X_3746_ _4422_/A _3827_/A vssd1 vssd1 vccd1 vccd1 _3762_/S sky130_fd_sc_hd__nor2_2
X_6465_ _6888_/CLK _6465_/D vssd1 vssd1 vccd1 vccd1 _6465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3677_ _3677_/A vssd1 vssd1 vccd1 vccd1 _6899_/D sky130_fd_sc_hd__clkbuf_1
X_5416_ _5415_/X _5435_/B vssd1 vssd1 vccd1 vccd1 _5416_/X sky130_fd_sc_hd__and2b_1
Xoutput120 _7117_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput142 _7139_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput131 _7102_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[5] sky130_fd_sc_hd__buf_2
X_6396_ _6430_/A _6396_/B vssd1 vssd1 vccd1 vccd1 _6397_/A sky130_fd_sc_hd__or2_1
Xoutput153 _7149_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[24] sky130_fd_sc_hd__buf_2
Xoutput164 _7130_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_114_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5148__212 _5150__214/A vssd1 vssd1 vccd1 vccd1 _6494_/CLK sky130_fd_sc_hd__inv_2
Xoutput175 _4689_/X vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
Xoutput186 _4993_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[19] sky130_fd_sc_hd__buf_2
X_5347_ _5366_/A _5346_/X _5250_/A vssd1 vssd1 vccd1 vccd1 _5347_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput197 _5015_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[29] sky130_fd_sc_hd__buf_2
X_5278_ _5302_/A vssd1 vssd1 vccd1 vccd1 _5364_/S sky130_fd_sc_hd__clkbuf_4
X_7017_ _7022_/CLK _7017_/D vssd1 vssd1 vccd1 vccd1 _7017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4229_ _3773_/X _6667_/Q _4233_/S vssd1 vssd1 vccd1 vccd1 _4230_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput22 caravel_wb_data_i[27] vssd1 vssd1 vccd1 vccd1 _5010_/B sky130_fd_sc_hd__buf_4
Xinput11 caravel_wb_data_i[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_2
X_4580_ _4487_/X _6506_/Q _4582_/S vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__mux2_1
X_3600_ _6929_/Q _3597_/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3601_/A sky130_fd_sc_hd__mux2_1
Xinput33 caravel_wb_data_i[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_2
X_3531_ _3531_/A vssd1 vssd1 vccd1 vccd1 _6959_/D sky130_fd_sc_hd__clkbuf_1
Xinput44 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 _7114_/A sky130_fd_sc_hd__buf_4
Xinput55 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 _7124_/A sky130_fd_sc_hd__buf_4
XFILLER_115_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput66 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 _7105_/A sky130_fd_sc_hd__buf_4
Xinput77 wbs_data_i[17] vssd1 vssd1 vccd1 vccd1 _7142_/A sky130_fd_sc_hd__buf_4
Xinput88 wbs_data_i[27] vssd1 vssd1 vccd1 vccd1 _7152_/A sky130_fd_sc_hd__buf_4
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6250_ _6250_/A _7001_/Q _6250_/C _6250_/D vssd1 vssd1 vccd1 vccd1 _6254_/D sky130_fd_sc_hd__and4_1
Xinput99 wbs_data_i[8] vssd1 vssd1 vccd1 vccd1 _7133_/A sky130_fd_sc_hd__clkbuf_8
X_3462_ _3788_/A vssd1 vssd1 vccd1 vccd1 _3462_/X sky130_fd_sc_hd__clkbuf_2
X_6181_ _6271_/A _6271_/B _6179_/X _6245_/A vssd1 vssd1 vccd1 vccd1 _6187_/B sky130_fd_sc_hd__a22o_1
X_3393_ _3392_/X _7047_/Q _3393_/S vssd1 vssd1 vccd1 vccd1 _3394_/A sky130_fd_sc_hd__mux2_1
X_5132_ _5138_/A vssd1 vssd1 vccd1 vccd1 _5132_/X sky130_fd_sc_hd__buf_1
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5063_ _6449_/Q _7103_/A _5071_/S vssd1 vssd1 vccd1 vccd1 _5064_/A sky130_fd_sc_hd__mux2_1
X_4014_ _4014_/A vssd1 vssd1 vccd1 vccd1 _4014_/X sky130_fd_sc_hd__buf_4
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2746_ clkbuf_0__2746_/X vssd1 vssd1 vccd1 vccd1 _5559__384/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5965_ _5965_/A vssd1 vssd1 vccd1 vccd1 _6875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5516__349 _5516__349/A vssd1 vssd1 vccd1 vccd1 _6639_/CLK sky130_fd_sc_hd__inv_2
X_4916_ _4944_/A _4915_/X _4802_/X vssd1 vssd1 vccd1 vccd1 _4916_/Y sky130_fd_sc_hd__o21ai_1
X_5896_ _6883_/Q _5609_/Y _5891_/Y _5894_/X _5895_/X vssd1 vssd1 vccd1 vccd1 _5922_/B
+ sky130_fd_sc_hd__o2111ai_1
X_4847_ _6855_/Q _6831_/Q _6807_/Q _6799_/Q _4814_/A _4845_/X vssd1 vssd1 vccd1 vccd1
+ _4847_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4778_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4778_/X sky130_fd_sc_hd__buf_6
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6517_ _6517_/CLK _6517_/D vssd1 vssd1 vccd1 vccd1 _6517_/Q sky130_fd_sc_hd__dfxtp_1
X_3729_ _3744_/S vssd1 vssd1 vccd1 vccd1 _3738_/S sky130_fd_sc_hd__buf_2
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6448_ _6696_/CLK _6448_/D vssd1 vssd1 vccd1 vccd1 _6448_/Q sky130_fd_sc_hd__dfxtp_1
X_6379_ _6696_/Q _6427_/C _7079_/Q vssd1 vssd1 vccd1 vccd1 _6379_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5750_ _5750_/A vssd1 vssd1 vccd1 vccd1 _5750_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__2531_ clkbuf_0__2531_/X vssd1 vssd1 vccd1 vccd1 _5235__283/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4701_ _4701_/A vssd1 vssd1 vccd1 vccd1 _4701_/X sky130_fd_sc_hd__buf_4
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4632_ _3853_/X _6483_/Q _4636_/S vssd1 vssd1 vccd1 vccd1 _4633_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4563_ _4563_/A vssd1 vssd1 vccd1 vccd1 _6514_/D sky130_fd_sc_hd__clkbuf_1
X_4494_ _4493_/X _6544_/Q _4500_/S vssd1 vssd1 vccd1 vccd1 _4495_/A sky130_fd_sc_hd__mux2_1
X_3514_ _6966_/Q _3450_/X _3516_/S vssd1 vssd1 vccd1 vccd1 _3515_/A sky130_fd_sc_hd__mux2_1
X_6302_ _6302_/A vssd1 vssd1 vccd1 vccd1 _6312_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6233_ _6241_/B _6237_/C vssd1 vssd1 vccd1 vccd1 _6234_/C sky130_fd_sc_hd__or2_1
Xclkbuf_1_1_0__3014_ clkbuf_0__3014_/X vssd1 vssd1 vccd1 vccd1 _6128_/A sky130_fd_sc_hd__clkbuf_4
X_3445_ _6992_/Q _3444_/X _3454_/S vssd1 vssd1 vccd1 vccd1 _3446_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6052__104 _6052__104/A vssd1 vssd1 vccd1 vccd1 _6912_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6164_ _4885_/X _6156_/Y _6163_/Y _4978_/X vssd1 vssd1 vccd1 vccd1 _6164_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3776_/A vssd1 vssd1 vccd1 vccd1 _3376_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5046_/X _5113_/X _6389_/A vssd1 vssd1 vccd1 vccd1 _6468_/D sky130_fd_sc_hd__o21a_1
X_5046_ _7079_/Q _5046_/B _6318_/C vssd1 vssd1 vccd1 vccd1 _5046_/X sky130_fd_sc_hd__and3_1
XFILLER_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6997_ _7093_/CLK _6997_/D vssd1 vssd1 vccd1 vccd1 _6997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5948_ _5951_/B _5944_/X _5947_/Y _5936_/X vssd1 vssd1 vccd1 vccd1 _5949_/B sky130_fd_sc_hd__a22o_1
Xclkbuf_1_1_0__2729_ clkbuf_0__2729_/X vssd1 vssd1 vccd1 vccd1 _5486_/A sky130_fd_sc_hd__clkbuf_4
X_5039__186 _5040__187/A vssd1 vssd1 vccd1 vccd1 _6442_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2876_ clkbuf_0__2876_/X vssd1 vssd1 vccd1 vccd1 _5862__61/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_4_0_wb_clk_i clkbuf_4_5_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6696_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6046__99 _6046__99/A vssd1 vssd1 vccd1 vccd1 _6907_/CLK sky130_fd_sc_hd__inv_2
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3230_ _6469_/Q _6468_/Q vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__or2_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6920_ _6920_/CLK _6920_/D vssd1 vssd1 vccd1 vccd1 _6920_/Q sky130_fd_sc_hd__dfxtp_1
X_6851_ _6851_/CLK _6851_/D vssd1 vssd1 vccd1 vccd1 _6851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2514_ clkbuf_0__2514_/X vssd1 vssd1 vccd1 vccd1 _5163_/A sky130_fd_sc_hd__clkbuf_4
X_3994_ _3994_/A vssd1 vssd1 vccd1 vccd1 _6766_/D sky130_fd_sc_hd__clkbuf_1
X_6782_ _6782_/CLK _6782_/D vssd1 vssd1 vccd1 vccd1 _6782_/Q sky130_fd_sc_hd__dfxtp_1
X_5733_ _5733_/A vssd1 vssd1 vccd1 vccd1 _6747_/D sky130_fd_sc_hd__clkbuf_1
X_5664_ _5664_/A _5913_/B _5664_/C _5664_/D vssd1 vssd1 vccd1 vccd1 _5898_/B sky130_fd_sc_hd__or4_2
X_4615_ _4615_/A vssd1 vssd1 vccd1 vccd1 _6491_/D sky130_fd_sc_hd__clkbuf_1
X_4546_ _4487_/X _6522_/Q _4548_/S vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__mux2_1
X_4477_ _4572_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4500_/S sky130_fd_sc_hd__or2_2
XFILLER_89_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2730_ clkbuf_0__2730_/X vssd1 vssd1 vccd1 vccd1 _5473__314/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6216_ _6216_/A _6216_/B _6216_/C vssd1 vssd1 vccd1 vccd1 _6217_/C sky130_fd_sc_hd__and3_1
X_3428_ _3428_/A vssd1 vssd1 vccd1 vccd1 _7035_/D sky130_fd_sc_hd__clkbuf_1
X_6147_ _6336_/A vssd1 vssd1 vccd1 vccd1 _6147_/X sky130_fd_sc_hd__buf_1
X_3359_ _4277_/A vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__clkbuf_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_24 _7131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_13 _4760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_35 _3862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_46 _7056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6078_ _6078_/A vssd1 vssd1 vccd1 vccd1 _6078_/X sky130_fd_sc_hd__buf_1
XFILLER_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5029_ _5175_/A vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__buf_1
XFILLER_81_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2859_ clkbuf_0__2859_/X vssd1 vssd1 vccd1 vccd1 _5780__476/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4400_ _3266_/X _6591_/Q _4402_/S vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__mux2_1
X_5380_ _6926_/Q _6918_/Q _7035_/Q _7051_/Q _4066_/A _5341_/X vssd1 vssd1 vccd1 vccd1
+ _5380_/X sky130_fd_sc_hd__mux4_2
X_4331_ _4331_/A vssd1 vssd1 vccd1 vccd1 _6622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7050_ _7050_/CLK _7050_/D vssd1 vssd1 vccd1 vccd1 _7050_/Q sky130_fd_sc_hd__dfxtp_1
X_4262_ _4262_/A vssd1 vssd1 vccd1 vccd1 _6653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3213_ _6731_/Q vssd1 vssd1 vccd1 vccd1 _3213_/Y sky130_fd_sc_hd__inv_2
X_6001_ _6882_/Q _5966_/A _6000_/X _5970_/A vssd1 vssd1 vccd1 vccd1 _6002_/B sky130_fd_sc_hd__a22o_1
X_4193_ _4193_/A vssd1 vssd1 vccd1 vccd1 _6683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6903_ _6903_/CLK _6903_/D vssd1 vssd1 vccd1 vccd1 _6903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6834_ _6834_/CLK _6834_/D vssd1 vssd1 vccd1 vccd1 _6834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6765_ _6765_/CLK _6765_/D vssd1 vssd1 vccd1 vccd1 _6765_/Q sky130_fd_sc_hd__dfxtp_1
X_3977_ _3977_/A _3977_/B vssd1 vssd1 vccd1 vccd1 _3981_/A sky130_fd_sc_hd__and2_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5716_ _5716_/A vssd1 vssd1 vccd1 vccd1 _5716_/X sky130_fd_sc_hd__buf_1
X_6696_ _6696_/CLK _6696_/D vssd1 vssd1 vccd1 vccd1 _6696_/Q sky130_fd_sc_hd__dfxtp_2
X_5647_ _6996_/Q vssd1 vssd1 vccd1 vccd1 _6216_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4529_ _4529_/A vssd1 vssd1 vccd1 vccd1 _6530_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5862__61 _5862__61/A vssd1 vssd1 vccd1 vccd1 _6847_/CLK sky130_fd_sc_hd__inv_2
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5197__252 _5199__254/A vssd1 vssd1 vccd1 vccd1 _6534_/CLK sky130_fd_sc_hd__inv_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6065__114 _6065__114/A vssd1 vssd1 vccd1 vccd1 _6922_/CLK sky130_fd_sc_hd__inv_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 caravel_wb_data_i[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_92_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5850__533 _5851__534/A vssd1 vssd1 vccd1 vccd1 _6839_/CLK sky130_fd_sc_hd__inv_2
X_4880_ _6546_/Q _6726_/Q _6864_/Q _6530_/Q _4906_/A _4898_/A vssd1 vssd1 vccd1 vccd1
+ _4880_/X sky130_fd_sc_hd__mux4_2
X_3900_ _6795_/Q _3597_/X _3908_/S vssd1 vssd1 vccd1 vccd1 _3901_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _6818_/Q _3602_/X _3837_/S vssd1 vssd1 vccd1 vccd1 _3832_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6550_ _6550_/CLK _6550_/D vssd1 vssd1 vccd1 vccd1 _6550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3762_ _6844_/Q _3620_/X _3762_/S vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3693_ _4020_/A vssd1 vssd1 vccd1 vccd1 _3693_/X sky130_fd_sc_hd__buf_2
X_6481_ _6481_/CLK _6481_/D vssd1 vssd1 vccd1 vccd1 _6481_/Q sky130_fd_sc_hd__dfxtp_1
X_5432_ _5430_/X _5431_/X _5432_/S vssd1 vssd1 vccd1 vccd1 _5432_/X sky130_fd_sc_hd__mux2_1
X_5363_ _6601_/Q _6585_/Q _6839_/Q _6823_/Q _5338_/A _5281_/X vssd1 vssd1 vccd1 vccd1
+ _5363_/X sky130_fd_sc_hd__mux4_1
X_7102_ _7102_/A vssd1 vssd1 vccd1 vccd1 _7102_/X sky130_fd_sc_hd__clkbuf_1
X_4314_ _4644_/A _4590_/A vssd1 vssd1 vccd1 vccd1 _4330_/S sky130_fd_sc_hd__nor2_2
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5294_ _5433_/S _5279_/X _5284_/Y _5287_/X _5293_/Y vssd1 vssd1 vccd1 vccd1 _5294_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_101_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4245_ _3770_/X _6660_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__mux2_1
X_7033_ _7033_/CLK _7033_/D vssd1 vssd1 vccd1 vccd1 _7033_/Q sky130_fd_sc_hd__dfxtp_1
X_4176_ _4020_/X _6690_/Q _4178_/S vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6817_ _6817_/CLK _6817_/D vssd1 vssd1 vccd1 vccd1 _6817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2876_ _5860_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2876_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6748_ _7022_/CLK _6748_/D vssd1 vssd1 vccd1 vccd1 _6748_/Q sky130_fd_sc_hd__dfxtp_2
X_6679_ _6679_/CLK _6679_/D vssd1 vssd1 vccd1 vccd1 _6679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4030_ _4029_/X _6752_/Q _4033_/S vssd1 vssd1 vccd1 vccd1 _4031_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5981_ _6878_/Q _5966_/X _5980_/Y _5970_/X vssd1 vssd1 vccd1 vccd1 _5982_/B sky130_fd_sc_hd__a22o_1
X_4932_ _6484_/Q _6556_/Q _7045_/Q _6976_/Q _4778_/X _4914_/X vssd1 vssd1 vccd1 vccd1
+ _4932_/X sky130_fd_sc_hd__mux4_1
XFILLER_18_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2730_ _5468_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2730_/X sky130_fd_sc_hd__clkbuf_16
X_4863_ _4909_/A _4863_/B vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__or2_1
X_6602_ _6602_/CLK _6602_/D vssd1 vssd1 vccd1 vccd1 _6602_/Q sky130_fd_sc_hd__dfxtp_1
X_4794_ _6447_/Q _4794_/B _4794_/C vssd1 vssd1 vccd1 vccd1 _4794_/X sky130_fd_sc_hd__and3_1
X_3814_ _3814_/A vssd1 vssd1 vccd1 vccd1 _6826_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6533_ _6533_/CLK _6533_/D vssd1 vssd1 vccd1 vccd1 _6533_/Q sky130_fd_sc_hd__dfxtp_1
X_3745_ _3745_/A vssd1 vssd1 vccd1 vccd1 _6852_/D sky130_fd_sc_hd__clkbuf_1
X_6464_ _7095_/CLK _6464_/D vssd1 vssd1 vccd1 vccd1 _6464_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput110 _7108_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[11] sky130_fd_sc_hd__buf_2
XFILLER_118_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3676_ _3349_/X _6899_/Q _3678_/S vssd1 vssd1 vccd1 vccd1 _3677_/A sky130_fd_sc_hd__mux2_1
X_5415_ _6794_/Q _6984_/Q _6992_/Q _6968_/Q _5341_/A _5276_/X vssd1 vssd1 vccd1 vccd1
+ _5415_/X sky130_fd_sc_hd__mux4_2
Xoutput121 _7118_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput143 _7140_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput132 _7103_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[6] sky130_fd_sc_hd__buf_2
X_6395_ _7137_/A _4978_/X _6407_/S vssd1 vssd1 vccd1 vccd1 _6396_/B sky130_fd_sc_hd__mux2_1
Xoutput154 _7150_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput165 _7131_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput176 _4758_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[0] sky130_fd_sc_hd__buf_2
X_5346_ _5334_/X _5336_/X _5340_/Y _5343_/X _5345_/Y vssd1 vssd1 vccd1 vccd1 _5346_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput187 _4800_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput198 _4833_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[2] sky130_fd_sc_hd__buf_2
X_5277_ _6788_/Q _6978_/Q _6986_/Q _6962_/Q _5264_/A _5276_/X vssd1 vssd1 vccd1 vccd1
+ _5277_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7016_ _7022_/CLK _7016_/D vssd1 vssd1 vccd1 vccd1 _7016_/Q sky130_fd_sc_hd__dfxtp_1
X_4228_ _4228_/A vssd1 vssd1 vccd1 vccd1 _6668_/D sky130_fd_sc_hd__clkbuf_1
X_6135__170 _6137__172/A vssd1 vssd1 vccd1 vccd1 _6978_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4159_ _6699_/Q _4158_/X _4165_/S vssd1 vssd1 vccd1 vccd1 _4160_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5571__393 _5572__394/A vssd1 vssd1 vccd1 vccd1 _6683_/CLK sky130_fd_sc_hd__inv_2
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2859_ _5778_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2859_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 caravel_wb_data_i[18] vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__buf_2
Xinput23 caravel_wb_data_i[28] vssd1 vssd1 vccd1 vccd1 _5012_/B sky130_fd_sc_hd__buf_4
Xinput34 caravel_wb_data_i[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_2
Xinput45 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 _7115_/A sky130_fd_sc_hd__buf_4
X_3530_ _6959_/Q _3447_/X _3534_/S vssd1 vssd1 vccd1 vccd1 _3531_/A sky130_fd_sc_hd__mux2_1
Xinput67 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 _7106_/A sky130_fd_sc_hd__buf_4
Xinput78 wbs_data_i[18] vssd1 vssd1 vccd1 vccd1 _7143_/A sky130_fd_sc_hd__buf_4
Xinput89 wbs_data_i[28] vssd1 vssd1 vccd1 vccd1 _7153_/A sky130_fd_sc_hd__buf_4
Xinput56 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 _4683_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3461_ _3461_/A vssd1 vssd1 vccd1 vccd1 _6987_/D sky130_fd_sc_hd__clkbuf_1
X_5200_ _5200_/A vssd1 vssd1 vccd1 vccd1 _5200_/X sky130_fd_sc_hd__buf_1
X_5032__181 _5033__182/A vssd1 vssd1 vccd1 vccd1 _6437_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6180_ _6180_/A vssd1 vssd1 vccd1 vccd1 _6245_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3392_ _3788_/A vssd1 vssd1 vccd1 vccd1 _3392_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5062_ _5588_/S vssd1 vssd1 vccd1 vccd1 _5071_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4013_ _4013_/A vssd1 vssd1 vccd1 vccd1 _6758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2745_ clkbuf_0__2745_/X vssd1 vssd1 vccd1 vccd1 _5553__379/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5964_ _5972_/A _5964_/B vssd1 vssd1 vccd1 vccd1 _5965_/A sky130_fd_sc_hd__and2_1
X_4915_ _6507_/Q _6441_/Q _6539_/Q _6691_/Q _4778_/X _4914_/X vssd1 vssd1 vccd1 vccd1
+ _4915_/X sky130_fd_sc_hd__mux4_2
X_5895_ _6877_/Q _5895_/B vssd1 vssd1 vccd1 vccd1 _5895_/X sky130_fd_sc_hd__xor2_1
X_4846_ _6505_/Q _6439_/Q _6537_/Q _6689_/Q _4814_/A _4845_/X vssd1 vssd1 vccd1 vccd1
+ _4846_/X sky130_fd_sc_hd__mux4_2
XFILLER_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6516_ _6516_/CLK _6516_/D vssd1 vssd1 vccd1 vccd1 _6516_/Q sky130_fd_sc_hd__dfxtp_1
X_4777_ _3977_/A _4772_/X _4776_/X vssd1 vssd1 vccd1 vccd1 _4777_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3728_ _4572_/A _3873_/B vssd1 vssd1 vccd1 vccd1 _3744_/S sky130_fd_sc_hd__or2_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3659_ _3353_/X _6906_/Q _3659_/S vssd1 vssd1 vccd1 vccd1 _3660_/A sky130_fd_sc_hd__mux2_1
X_6447_ _6696_/CLK _6447_/D vssd1 vssd1 vccd1 vccd1 _6447_/Q sky130_fd_sc_hd__dfxtp_1
X_6378_ _6696_/Q _6427_/C vssd1 vssd1 vccd1 vccd1 _6381_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1_0__3159_ clkbuf_0__3159_/X vssd1 vssd1 vccd1 vccd1 _6372__54/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5329_ _5329_/A vssd1 vssd1 vccd1 vccd1 _5329_/X sky130_fd_sc_hd__buf_2
XFILLER_87_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5677__413 _5678__414/A vssd1 vssd1 vccd1 vccd1 _6707_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5578__399 _5578__399/A vssd1 vssd1 vccd1 vccd1 _6689_/CLK sky130_fd_sc_hd__inv_2
XFILLER_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2530_ clkbuf_0__2530_/X vssd1 vssd1 vccd1 vccd1 _5230__279/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4700_ _4851_/S vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__buf_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4631_ _4631_/A vssd1 vssd1 vccd1 vccd1 _6484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4562_ _6514_/Q _4020_/A _4562_/S vssd1 vssd1 vccd1 vccd1 _4563_/A sky130_fd_sc_hd__mux2_1
X_6301_ input1/X _6284_/A _6300_/X _6247_/A vssd1 vssd1 vccd1 vccd1 _7022_/D sky130_fd_sc_hd__o211a_1
X_4493_ _6743_/Q vssd1 vssd1 vccd1 vccd1 _4493_/X sky130_fd_sc_hd__buf_2
X_3513_ _3513_/A vssd1 vssd1 vccd1 vccd1 _6967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6232_ _6241_/B _6237_/C vssd1 vssd1 vccd1 vccd1 _6234_/B sky130_fd_sc_hd__nand2_1
X_3444_ _3770_/A vssd1 vssd1 vccd1 vccd1 _3444_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__3013_ clkbuf_0__3013_/X vssd1 vssd1 vccd1 vccd1 _6114__154/A sky130_fd_sc_hd__clkbuf_4
X_6163_ _7007_/Q vssd1 vssd1 vccd1 vccd1 _6163_/Y sky130_fd_sc_hd__inv_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _7027_/Q vssd1 vssd1 vccd1 vccd1 _3776_/A sky130_fd_sc_hd__clkbuf_4
X_5522__354 _5522__354/A vssd1 vssd1 vccd1 vccd1 _6644_/CLK sky130_fd_sc_hd__inv_2
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _6391_/A vssd1 vssd1 vccd1 vccd1 _6389_/A sky130_fd_sc_hd__clkbuf_2
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _6302_/A vssd1 vssd1 vccd1 vccd1 _6318_/C sky130_fd_sc_hd__buf_2
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6996_ _7093_/CLK _6996_/D vssd1 vssd1 vccd1 vccd1 _6996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5947_ _5952_/B _5947_/B vssd1 vssd1 vccd1 vccd1 _5947_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1_0__2728_ clkbuf_0__2728_/X vssd1 vssd1 vccd1 vccd1 _5466__309/A sky130_fd_sc_hd__clkbuf_4
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5191__247 _5193__249/A vssd1 vssd1 vccd1 vccd1 _6529_/CLK sky130_fd_sc_hd__inv_2
X_5878_ _5878_/A vssd1 vssd1 vccd1 vccd1 _5878_/X sky130_fd_sc_hd__buf_1
X_4829_ _4822_/Y _4824_/Y _4826_/Y _4828_/Y _4724_/A vssd1 vssd1 vccd1 vccd1 _4830_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5869__67 _5871__69/A vssd1 vssd1 vccd1 vccd1 _6853_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5465__308 _5466__309/A vssd1 vssd1 vccd1 vccd1 _6598_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5814__504 _5814__504/A vssd1 vssd1 vccd1 vccd1 _6810_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6850_ _6850_/CLK _6850_/D vssd1 vssd1 vccd1 vccd1 _6850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6781_ _6781_/CLK _6781_/D vssd1 vssd1 vccd1 vccd1 _6781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5732_ _7021_/Q _5734_/B vssd1 vssd1 vccd1 vccd1 _5733_/A sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__2513_ clkbuf_0__2513_/X vssd1 vssd1 vccd1 vccd1 _5143__209/A sky130_fd_sc_hd__clkbuf_4
X_3993_ _3680_/X _6766_/Q _4001_/S vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5663_ _5663_/A _7086_/Q _5892_/A vssd1 vssd1 vccd1 vccd1 _5664_/D sky130_fd_sc_hd__or3_1
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4614_ _3853_/X _6491_/Q _4618_/S vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _6523_/D sky130_fd_sc_hd__clkbuf_1
X_4476_ _6748_/Q vssd1 vssd1 vccd1 vccd1 _4476_/X sky130_fd_sc_hd__buf_2
X_6215_ _6215_/A vssd1 vssd1 vccd1 vccd1 _6999_/D sky130_fd_sc_hd__clkbuf_1
X_3427_ _3376_/X _7035_/Q _3429_/S vssd1 vssd1 vccd1 vccd1 _3428_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6146_ _6342_/A vssd1 vssd1 vccd1 vccd1 _6146_/X sky130_fd_sc_hd__buf_1
XFILLER_58_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3358_ _6739_/Q vssd1 vssd1 vccd1 vccd1 _4277_/A sky130_fd_sc_hd__clkbuf_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_25 _4502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_14 _4760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XINSDIODE2_36 _3862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_47 _7130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3289_ _7064_/Q _3266_/X _3291_/S vssd1 vssd1 vccd1 vccd1 _3290_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5028_ _5597_/A vssd1 vssd1 vccd1 vccd1 _5028_/X sky130_fd_sc_hd__buf_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6979_ _6979_/CLK _6979_/D vssd1 vssd1 vccd1 vccd1 _6979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5471__312 _5473__314/A vssd1 vssd1 vccd1 vccd1 _6602_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ _6622_/Q _3895_/X _4330_/S vssd1 vssd1 vccd1 vccd1 _4331_/A sky130_fd_sc_hd__mux2_1
X_4261_ _6653_/Q _4141_/X _4269_/S vssd1 vssd1 vccd1 vccd1 _4262_/A sky130_fd_sc_hd__mux2_1
X_3212_ _6737_/Q _6732_/Q vssd1 vssd1 vccd1 vccd1 _3221_/B sky130_fd_sc_hd__xor2_1
X_6000_ _6882_/Q _6004_/C vssd1 vssd1 vccd1 vccd1 _6000_/X sky130_fd_sc_hd__xor2_1
X_5142__208 _5143__209/A vssd1 vssd1 vccd1 vccd1 _6490_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4192_ _6683_/Q _4149_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4193_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6902_ _6902_/CLK _6902_/D vssd1 vssd1 vccd1 vccd1 _6902_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6833_ _6833_/CLK _6833_/D vssd1 vssd1 vccd1 vccd1 _6833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6764_ _6764_/CLK _6764_/D vssd1 vssd1 vccd1 vccd1 _6764_/Q sky130_fd_sc_hd__dfxtp_1
X_3976_ _3976_/A vssd1 vssd1 vccd1 vccd1 _6770_/D sky130_fd_sc_hd__clkbuf_1
X_6695_ _5852_/A _6695_/D vssd1 vssd1 vccd1 vccd1 _6695_/Q sky130_fd_sc_hd__dfxtp_2
X_5646_ _7091_/Q _5664_/A _5652_/C vssd1 vssd1 vccd1 vccd1 _5653_/A sky130_fd_sc_hd__o21ba_1
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4528_ _4487_/X _6530_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4529_/A sky130_fd_sc_hd__mux2_1
X_4459_ _4474_/S vssd1 vssd1 vccd1 vccd1 _4468_/S sky130_fd_sc_hd__buf_2
XFILLER_105_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5535__364 _5535__364/A vssd1 vssd1 vccd1 vccd1 _6654_/CLK sky130_fd_sc_hd__inv_2
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _3830_/A vssd1 vssd1 vccd1 vccd1 _6819_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3761_ _3761_/A vssd1 vssd1 vccd1 vccd1 _6845_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3692_ _3692_/A vssd1 vssd1 vccd1 vccd1 _6894_/D sky130_fd_sc_hd__clkbuf_1
X_6480_ _6480_/CLK _6480_/D vssd1 vssd1 vccd1 vccd1 _6480_/Q sky130_fd_sc_hd__dfxtp_1
X_5431_ _6605_/Q _6589_/Q _6843_/Q _6827_/Q _5329_/X _5330_/X vssd1 vssd1 vccd1 vccd1
+ _5431_/X sky130_fd_sc_hd__mux4_1
X_5362_ _6641_/Q _6633_/Q _6617_/Q _6609_/Q _5330_/A _5290_/X vssd1 vssd1 vccd1 vccd1
+ _5362_/X sky130_fd_sc_hd__mux4_1
X_7101_ _7101_/A vssd1 vssd1 vccd1 vccd1 _7101_/X sky130_fd_sc_hd__clkbuf_1
X_4313_ _4313_/A vssd1 vssd1 vccd1 vccd1 _6630_/D sky130_fd_sc_hd__clkbuf_1
X_5293_ _5289_/X _5291_/X _5292_/X vssd1 vssd1 vccd1 vccd1 _5293_/Y sky130_fd_sc_hd__o21ai_1
X_7032_ _7032_/CLK _7032_/D vssd1 vssd1 vccd1 vccd1 _7032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4244_ _4244_/A vssd1 vssd1 vccd1 vccd1 _6661_/D sky130_fd_sc_hd__clkbuf_1
X_4175_ _4175_/A vssd1 vssd1 vccd1 vccd1 _6691_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5478__318 _5478__318/A vssd1 vssd1 vccd1 vccd1 _6608_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6816_ _6816_/CLK _6816_/D vssd1 vssd1 vccd1 vccd1 _6816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__2875_ _5854_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2875_/X sky130_fd_sc_hd__clkbuf_16
X_6747_ _7022_/CLK _6747_/D vssd1 vssd1 vccd1 vccd1 _6747_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3959_ _3959_/A vssd1 vssd1 vccd1 vccd1 _3977_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5827__514 _5827__514/A vssd1 vssd1 vccd1 vccd1 _6820_/CLK sky130_fd_sc_hd__inv_2
X_6678_ _6678_/CLK _6678_/D vssd1 vssd1 vccd1 vccd1 _6678_/Q sky130_fd_sc_hd__dfxtp_1
X_5629_ _5892_/B _6175_/A vssd1 vssd1 vccd1 vccd1 _5642_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5212__264 _5212__264/A vssd1 vssd1 vccd1 vccd1 _6546_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _5985_/B _5980_/B vssd1 vssd1 vccd1 vccd1 _5980_/Y sky130_fd_sc_hd__nor2_1
X_4931_ _6904_/Q _6564_/Q _6912_/Q _6492_/Q _4906_/X _3966_/X vssd1 vssd1 vccd1 vccd1
+ _4931_/X sky130_fd_sc_hd__mux4_1
XFILLER_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4862_ _6506_/Q _6440_/Q _6538_/Q _6690_/Q _4814_/A _4845_/X vssd1 vssd1 vccd1 vccd1
+ _4863_/B sky130_fd_sc_hd__mux4_2
XFILLER_60_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3813_ _6826_/Q _3602_/X _3819_/S vssd1 vssd1 vccd1 vccd1 _3814_/A sky130_fd_sc_hd__mux2_1
X_6601_ _6601_/CLK _6601_/D vssd1 vssd1 vccd1 vccd1 _6601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4793_ _4726_/X _4788_/X _4790_/Y _4792_/Y vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6532_ _6532_/CLK _6532_/D vssd1 vssd1 vccd1 vccd1 _6532_/Q sky130_fd_sc_hd__dfxtp_1
X_3744_ _3705_/X _6852_/Q _3744_/S vssd1 vssd1 vccd1 vccd1 _3745_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3675_ _3675_/A vssd1 vssd1 vccd1 vccd1 _6900_/D sky130_fd_sc_hd__clkbuf_1
X_6463_ _6897_/CLK _6463_/D vssd1 vssd1 vccd1 vccd1 _6463_/Q sky130_fd_sc_hd__dfxtp_1
X_5414_ _5410_/X _5413_/X _5433_/S vssd1 vssd1 vccd1 vccd1 _5414_/X sky130_fd_sc_hd__mux2_1
Xoutput122 _7119_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput111 _7109_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[12] sky130_fd_sc_hd__buf_2
Xoutput133 _7104_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[7] sky130_fd_sc_hd__buf_2
XFILLER_114_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6394_ _6394_/A vssd1 vssd1 vccd1 vccd1 _7083_/D sky130_fd_sc_hd__clkbuf_1
Xoutput155 _7151_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput144 _7141_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[16] sky130_fd_sc_hd__buf_2
Xoutput166 _7132_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_114_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput177 _4975_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[10] sky130_fd_sc_hd__buf_2
X_5345_ _5289_/X _5344_/X _5292_/X vssd1 vssd1 vccd1 vccd1 _5345_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput188 _4996_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[20] sky130_fd_sc_hd__buf_2
Xoutput199 _5017_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[30] sky130_fd_sc_hd__buf_2
X_5276_ _5281_/A vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__buf_2
X_7015_ _7019_/CLK _7015_/D vssd1 vssd1 vccd1 vccd1 _7015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4227_ _3770_/X _6668_/Q _4233_/S vssd1 vssd1 vccd1 vccd1 _4228_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4158_ _7025_/Q vssd1 vssd1 vccd1 vccd1 _4158_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4089_ _4009_/X _6729_/Q _4097_/S vssd1 vssd1 vccd1 vccd1 _4090_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5155__218 _5155__218/A vssd1 vssd1 vccd1 vccd1 _6500_/CLK sky130_fd_sc_hd__inv_2
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 caravel_wb_data_i[19] vssd1 vssd1 vccd1 vccd1 _4992_/B sky130_fd_sc_hd__buf_2
Xinput24 caravel_wb_data_i[29] vssd1 vssd1 vccd1 vccd1 _5014_/B sky130_fd_sc_hd__buf_4
Xinput35 wb_rst_i vssd1 vssd1 vccd1 vccd1 _5047_/A sky130_fd_sc_hd__buf_6
Xinput46 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 _7116_/A sky130_fd_sc_hd__buf_4
Xinput68 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 _5050_/B sky130_fd_sc_hd__clkbuf_2
Xinput79 wbs_data_i[19] vssd1 vssd1 vccd1 vccd1 _7144_/A sky130_fd_sc_hd__buf_4
Xinput57 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 _4683_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3460_ _6987_/Q _3459_/X _3463_/S vssd1 vssd1 vccd1 vccd1 _3461_/A sky130_fd_sc_hd__mux2_1
X_3391_ _7023_/Q vssd1 vssd1 vccd1 vccd1 _3788_/A sky130_fd_sc_hd__buf_4
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5061_ _5061_/A vssd1 vssd1 vccd1 vccd1 _5588_/S sky130_fd_sc_hd__buf_2
X_4012_ _4009_/X _6758_/Q _4024_/S vssd1 vssd1 vccd1 vccd1 _4013_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5963_ _6875_/Q _5944_/X _5962_/Y _5936_/X vssd1 vssd1 vccd1 vccd1 _5964_/B sky130_fd_sc_hd__a22o_1
XFILLER_25_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2744_ clkbuf_0__2744_/X vssd1 vssd1 vccd1 vccd1 _5544__371/A sky130_fd_sc_hd__clkbuf_4
X_4914_ _4914_/A vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__buf_4
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5894_ _5898_/B _5898_/C _5994_/B vssd1 vssd1 vccd1 vccd1 _5894_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4845_ _4845_/A vssd1 vssd1 vccd1 vccd1 _4845_/X sky130_fd_sc_hd__buf_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4776_ _4774_/X _4775_/X _4826_/A vssd1 vssd1 vccd1 vccd1 _4776_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6515_ _6515_/CLK _6515_/D vssd1 vssd1 vccd1 vccd1 _6515_/Q sky130_fd_sc_hd__dfxtp_1
X_3727_ _3990_/B _3727_/B _3990_/C vssd1 vssd1 vccd1 vccd1 _3873_/B sky130_fd_sc_hd__nand3b_4
X_3658_ _3658_/A vssd1 vssd1 vccd1 vccd1 _6907_/D sky130_fd_sc_hd__clkbuf_1
X_6446_ _5852_/A _6446_/D vssd1 vssd1 vccd1 vccd1 _6446_/Q sky130_fd_sc_hd__dfxtp_1
X_6377_ _6377_/A _6377_/B vssd1 vssd1 vccd1 vccd1 _6427_/C sky130_fd_sc_hd__nor2_2
X_3589_ _6933_/Q _3453_/X _3589_/S vssd1 vssd1 vccd1 vccd1 _3590_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3158_ clkbuf_0__3158_/X vssd1 vssd1 vccd1 vccd1 _6363__46/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5328_ _6640_/Q _6632_/Q _6616_/Q _6608_/Q _5263_/X _5264_/X vssd1 vssd1 vccd1 vccd1
+ _5328_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5259_ _5264_/A vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__buf_2
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _3850_/X _6484_/Q _4636_/S vssd1 vssd1 vccd1 vccd1 _4631_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4561_ _4561_/A vssd1 vssd1 vccd1 vccd1 _6515_/D sky130_fd_sc_hd__clkbuf_1
X_6300_ _7022_/Q _6300_/B vssd1 vssd1 vccd1 vccd1 _6300_/X sky130_fd_sc_hd__or2_1
XFILLER_116_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4492_ _4492_/A vssd1 vssd1 vccd1 vccd1 _6545_/D sky130_fd_sc_hd__clkbuf_1
X_3512_ _6967_/Q _3447_/X _3516_/S vssd1 vssd1 vccd1 vccd1 _3513_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6231_ _7003_/Q vssd1 vssd1 vccd1 vccd1 _6241_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3443_ _3443_/A vssd1 vssd1 vccd1 vccd1 _6993_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3012_ clkbuf_0__3012_/X vssd1 vssd1 vccd1 vccd1 _6104__145/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6162_ _7005_/Q vssd1 vssd1 vccd1 vccd1 _6162_/Y sky130_fd_sc_hd__inv_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _7161_/A _5113_/B _5113_/C vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__and3_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3374_/A vssd1 vssd1 vccd1 vccd1 _7052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A _5044_/B _5044_/C vssd1 vssd1 vccd1 vccd1 _6302_/A sky130_fd_sc_hd__and3_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6995_ _7022_/CLK _6995_/D vssd1 vssd1 vccd1 vccd1 _6995_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5946_ _5951_/C _5945_/C _5951_/B vssd1 vssd1 vccd1 vccd1 _5947_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_1_1_0__2727_ clkbuf_0__2727_/X vssd1 vssd1 vccd1 vccd1 _5458__302/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4828_ _4716_/A _4827_/X _4802_/A vssd1 vssd1 vccd1 vccd1 _4828_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4759_ _7095_/Q vssd1 vssd1 vccd1 vccd1 _5648_/A sky130_fd_sc_hd__clkbuf_2
X_6429_ _7126_/A _4760_/X _6432_/S vssd1 vssd1 vccd1 vccd1 _6430_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2874_ clkbuf_0__2874_/X vssd1 vssd1 vccd1 vccd1 _5866_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _4007_/S vssd1 vssd1 vccd1 vccd1 _4001_/S sky130_fd_sc_hd__buf_2
X_6780_ _6780_/CLK _6780_/D vssd1 vssd1 vccd1 vccd1 _6780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__2735_ clkbuf_0__2735_/X vssd1 vssd1 vccd1 vccd1 _5523_/A sky130_fd_sc_hd__clkbuf_16
X_5731_ _5731_/A vssd1 vssd1 vccd1 vccd1 _6746_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__2512_ clkbuf_0__2512_/X vssd1 vssd1 vccd1 vccd1 _5137__204/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5662_ _5888_/C _5610_/X _6266_/A vssd1 vssd1 vccd1 vccd1 _5662_/X sky130_fd_sc_hd__a21o_1
X_4613_ _4613_/A vssd1 vssd1 vccd1 vccd1 _6492_/D sky130_fd_sc_hd__clkbuf_1
X_4544_ _4484_/X _6523_/Q _4548_/S vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4475_ _4475_/A vssd1 vssd1 vccd1 vccd1 _6550_/D sky130_fd_sc_hd__clkbuf_1
X_6214_ _6238_/A _6214_/B _6214_/C vssd1 vssd1 vccd1 vccd1 _6215_/A sky130_fd_sc_hd__and3_1
X_3426_ _3426_/A vssd1 vssd1 vccd1 vccd1 _7036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3357_ _3764_/A vssd1 vssd1 vccd1 vccd1 _3357_/X sky130_fd_sc_hd__buf_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5874__71 _5877__74/A vssd1 vssd1 vccd1 vccd1 _6857_/CLK sky130_fd_sc_hd__inv_2
XINSDIODE2_15 _4863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XINSDIODE2_48 _3868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_37 _3868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5027_ _5852_/A vssd1 vssd1 vccd1 vccd1 _5027_/X sky130_fd_sc_hd__buf_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_26 _3597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3288_ _3288_/A vssd1 vssd1 vccd1 vccd1 _7065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6036__90 _6038__92/A vssd1 vssd1 vccd1 vccd1 _6898_/CLK sky130_fd_sc_hd__inv_2
X_6978_ _6978_/CLK _6978_/D vssd1 vssd1 vccd1 vccd1 _6978_/Q sky130_fd_sc_hd__dfxtp_1
X_5929_ _5929_/A _5929_/B _6017_/A vssd1 vssd1 vccd1 vccd1 _5966_/A sky130_fd_sc_hd__nor3_2
XFILLER_119_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2857_ clkbuf_0__2857_/X vssd1 vssd1 vccd1 vccd1 _5773__473/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4260_ _4275_/S vssd1 vssd1 vccd1 vccd1 _4269_/S sky130_fd_sc_hd__buf_2
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4191_ _4191_/A vssd1 vssd1 vccd1 vccd1 _6684_/D sky130_fd_sc_hd__clkbuf_1
X_3211_ _6738_/Q _6733_/Q vssd1 vssd1 vccd1 vccd1 _3221_/A sky130_fd_sc_hd__xor2_1
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5777__474 _5777__474/A vssd1 vssd1 vccd1 vccd1 _6780_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6901_ _6901_/CLK _6901_/D vssd1 vssd1 vccd1 vccd1 _6901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6832_ _6832_/CLK _6832_/D vssd1 vssd1 vccd1 vccd1 _6832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6763_ _6763_/CLK _6763_/D vssd1 vssd1 vccd1 vccd1 _6763_/Q sky130_fd_sc_hd__dfxtp_1
X_3975_ _5774_/C _3975_/B _3975_/C vssd1 vssd1 vccd1 vccd1 _3976_/A sky130_fd_sc_hd__and3_1
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6694_ _5852_/A _6694_/D vssd1 vssd1 vccd1 vccd1 _6694_/Q sky130_fd_sc_hd__dfxtp_1
X_5645_ _7090_/Q _7001_/Q vssd1 vssd1 vccd1 vccd1 _5652_/C sky130_fd_sc_hd__xnor2_1
XFILLER_108_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4527_ _4527_/A vssd1 vssd1 vccd1 vccd1 _6531_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4458_ _4458_/A _4626_/A vssd1 vssd1 vccd1 vccd1 _4474_/S sky130_fd_sc_hd__or2_2
XFILLER_104_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3409_ _3409_/A vssd1 vssd1 vccd1 vccd1 _7043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6128_ _6128_/A vssd1 vssd1 vccd1 vccd1 _6128_/X sky130_fd_sc_hd__buf_1
X_4389_ _4389_/A vssd1 vssd1 vccd1 vccd1 _6597_/D sky130_fd_sc_hd__clkbuf_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3760_ _6845_/Q _3617_/X _3762_/S vssd1 vssd1 vccd1 vccd1 _3761_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3691_ _3690_/X _6894_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3692_/A sky130_fd_sc_hd__mux2_1
X_5430_ _6645_/Q _6637_/Q _6621_/Q _6613_/Q _4083_/A _4063_/A vssd1 vssd1 vccd1 vccd1
+ _5430_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5705__435 _5705__435/A vssd1 vssd1 vccd1 vccd1 _6729_/CLK sky130_fd_sc_hd__inv_2
X_5361_ _5359_/X _5360_/X _5364_/S vssd1 vssd1 vccd1 vccd1 _5361_/X sky130_fd_sc_hd__mux2_1
X_7100_ _7100_/A vssd1 vssd1 vccd1 vccd1 _7100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4312_ _3788_/X _6630_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__mux2_1
X_5292_ _6733_/Q vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4243_ _3764_/X _6661_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__mux2_1
X_7031_ _7031_/CLK _7031_/D vssd1 vssd1 vccd1 vccd1 _7031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5601__411 _5601__411/A vssd1 vssd1 vccd1 vccd1 _6704_/CLK sky130_fd_sc_hd__inv_2
X_4174_ _4017_/X _6691_/Q _4178_/S vssd1 vssd1 vccd1 vccd1 _4175_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5751__455 _5752__456/A vssd1 vssd1 vccd1 vccd1 _6759_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2874_ _5853_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2874_/X sky130_fd_sc_hd__clkbuf_16
X_6815_ _6815_/CLK _6815_/D vssd1 vssd1 vccd1 vccd1 _6815_/Q sky130_fd_sc_hd__dfxtp_1
X_6746_ _7022_/CLK _6746_/D vssd1 vssd1 vccd1 vccd1 _6746_/Q sky130_fd_sc_hd__dfxtp_2
X_3958_ _3958_/A vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3889_ _6743_/Q vssd1 vssd1 vccd1 vccd1 _3889_/X sky130_fd_sc_hd__clkbuf_4
X_6677_ _6677_/CLK _6677_/D vssd1 vssd1 vccd1 vccd1 _6677_/Q sky130_fd_sc_hd__dfxtp_1
X_5628_ _5892_/B _6175_/A vssd1 vssd1 vccd1 vccd1 _5642_/A sky130_fd_sc_hd__and2_1
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5583__403 _5583__403/A vssd1 vssd1 vccd1 vccd1 _6693_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6048__100 _6049__101/A vssd1 vssd1 vccd1 vccd1 _6908_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4930_ _4922_/X _4925_/X _4927_/X _4929_/X _3951_/Y vssd1 vssd1 vccd1 vccd1 _4930_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4861_ _4691_/X input28/X _4695_/X _4860_/X vssd1 vssd1 vccd1 vccd1 _4861_/X sky130_fd_sc_hd__a22o_2
XFILLER_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3812_ _3812_/A vssd1 vssd1 vccd1 vccd1 _6827_/D sky130_fd_sc_hd__clkbuf_1
X_6600_ _6600_/CLK _6600_/D vssd1 vssd1 vccd1 vccd1 _6600_/Q sky130_fd_sc_hd__dfxtp_1
X_4792_ _4933_/S _4791_/X _4711_/X vssd1 vssd1 vccd1 vccd1 _4792_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6531_ _6531_/CLK _6531_/D vssd1 vssd1 vccd1 vccd1 _6531_/Q sky130_fd_sc_hd__dfxtp_1
X_3743_ _3743_/A vssd1 vssd1 vccd1 vccd1 _6853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3674_ _3345_/X _6900_/Q _3678_/S vssd1 vssd1 vccd1 vccd1 _3675_/A sky130_fd_sc_hd__mux2_1
X_6462_ _7089_/CLK _6462_/D vssd1 vssd1 vccd1 vccd1 _6462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6393_ _6408_/A _6393_/B vssd1 vssd1 vccd1 vccd1 _6394_/A sky130_fd_sc_hd__and2_1
X_5413_ _5411_/X _5412_/X _5432_/S vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__mux2_1
X_5484__323 _5485__324/A vssd1 vssd1 vccd1 vccd1 _6613_/CLK sky130_fd_sc_hd__inv_2
Xoutput123 _7120_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput112 _7110_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[13] sky130_fd_sc_hd__buf_2
Xoutput134 _7105_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[8] sky130_fd_sc_hd__buf_2
X_5344_ _6956_/Q _6940_/Q _7065_/Q _6932_/Q _5290_/X _4069_/A vssd1 vssd1 vccd1 vccd1
+ _5344_/X sky130_fd_sc_hd__mux4_1
Xoutput156 _7152_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput145 _7142_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[17] sky130_fd_sc_hd__buf_2
Xoutput167 _7133_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[8] sky130_fd_sc_hd__buf_2
X_6321__12 _6323__14/A vssd1 vssd1 vccd1 vccd1 _7032_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput189 _4998_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[21] sky130_fd_sc_hd__buf_2
Xoutput178 _4977_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[11] sky130_fd_sc_hd__buf_2
X_5275_ _5334_/A vssd1 vssd1 vccd1 vccd1 _5433_/S sky130_fd_sc_hd__clkbuf_4
X_7014_ _7019_/CLK _7014_/D vssd1 vssd1 vccd1 vccd1 _7014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4226_ _4226_/A vssd1 vssd1 vccd1 vccd1 _6669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4157_ _4157_/A vssd1 vssd1 vccd1 vccd1 _6700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4088_ _4103_/S vssd1 vssd1 vccd1 vccd1 _4097_/S sky130_fd_sc_hd__buf_2
XFILLER_102_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2857_ _5769_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2857_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6729_ _6729_/CLK _6729_/D vssd1 vssd1 vccd1 vccd1 _6729_/Q sky130_fd_sc_hd__dfxtp_1
X_6142__176 _6143__177/A vssd1 vssd1 vccd1 vccd1 _6984_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput25 caravel_wb_data_i[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_2
Xinput14 caravel_wb_data_i[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_2
Xinput36 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 _7097_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_116_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 _7098_/A sky130_fd_sc_hd__clkbuf_1
Xinput58 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 _7099_/A sky130_fd_sc_hd__buf_4
Xinput69 wbs_data_i[0] vssd1 vssd1 vccd1 vccd1 _7125_/A sky130_fd_sc_hd__buf_8
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3390_ _3390_/A vssd1 vssd1 vccd1 vccd1 _7048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5060_ _5060_/A vssd1 vssd1 vccd1 vccd1 _6448_/D sky130_fd_sc_hd__clkbuf_1
X_4011_ _4033_/S vssd1 vssd1 vccd1 vccd1 _4024_/S sky130_fd_sc_hd__buf_2
XFILLER_96_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5962_ _5962_/A _5968_/B vssd1 vssd1 vccd1 vccd1 _5962_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1_0__2743_ clkbuf_0__2743_/X vssd1 vssd1 vccd1 vccd1 _5541__369/A sky130_fd_sc_hd__clkbuf_4
X_4913_ _4927_/A _4913_/B vssd1 vssd1 vccd1 vccd1 _4913_/Y sky130_fd_sc_hd__nor2_1
X_5893_ _6880_/Q vssd1 vssd1 vccd1 vccd1 _5994_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4844_ _4722_/X _4836_/X _4841_/X _4843_/X _4724_/A vssd1 vssd1 vccd1 vccd1 _4844_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4775_ _6479_/Q _6551_/Q _4936_/S vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6514_ _6514_/CLK _6514_/D vssd1 vssd1 vccd1 vccd1 _6514_/Q sky130_fd_sc_hd__dfxtp_1
X_3726_ _3726_/A vssd1 vssd1 vccd1 vccd1 _6860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3657_ _3349_/X _6907_/Q _3659_/S vssd1 vssd1 vccd1 vccd1 _3658_/A sky130_fd_sc_hd__mux2_1
X_6445_ _5852_/A _6445_/D vssd1 vssd1 vccd1 vccd1 _6445_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__3157_ clkbuf_0__3157_/X vssd1 vssd1 vccd1 vccd1 _6358__42/A sky130_fd_sc_hd__clkbuf_4
X_3588_ _3588_/A vssd1 vssd1 vccd1 vccd1 _6934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5327_ _5325_/X _5326_/X _5410_/S vssd1 vssd1 vccd1 vccd1 _5327_/X sky130_fd_sc_hd__mux2_1
XFILLER_114_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5258_ _5258_/A vssd1 vssd1 vccd1 vccd1 _5264_/A sky130_fd_sc_hd__buf_4
X_5161__223 _5162__224/A vssd1 vssd1 vccd1 vccd1 _6505_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4209_ _6676_/Q _4146_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5684__419 _5684__419/A vssd1 vssd1 vccd1 vccd1 _6713_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5764__465 _5766__467/A vssd1 vssd1 vccd1 vccd1 _6769_/CLK sky130_fd_sc_hd__inv_2
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4560_ _6515_/Q _4017_/A _4562_/S vssd1 vssd1 vccd1 vccd1 _4561_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4491_ _4490_/X _6545_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4492_/A sky130_fd_sc_hd__mux2_1
X_3511_ _3511_/A vssd1 vssd1 vccd1 vccd1 _6968_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3011_ clkbuf_0__3011_/X vssd1 vssd1 vccd1 vccd1 _6099__141/A sky130_fd_sc_hd__clkbuf_4
X_6230_ _6230_/A vssd1 vssd1 vccd1 vccd1 _7002_/D sky130_fd_sc_hd__clkbuf_1
X_3442_ _6993_/Q _3437_/X _3454_/S vssd1 vssd1 vccd1 vccd1 _3443_/A sky130_fd_sc_hd__mux2_1
X_6161_ _6161_/A vssd1 vssd1 vccd1 vccd1 _6161_/Y sky130_fd_sc_hd__inv_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _3372_/X _7052_/Q _3381_/S vssd1 vssd1 vccd1 vccd1 _3374_/A sky130_fd_sc_hd__mux2_1
X_5886__80 _5887__81/A vssd1 vssd1 vccd1 vccd1 _6866_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5924_/D _5929_/B _5972_/A _5111_/X vssd1 vssd1 vccd1 vccd1 _6467_/D sky130_fd_sc_hd__o211a_2
XFILLER_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _6381_/A _5043_/B vssd1 vssd1 vccd1 vccd1 _5046_/B sky130_fd_sc_hd__nor2_1
XFILLER_65_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6994_ _7093_/CLK _6994_/D vssd1 vssd1 vccd1 vccd1 _6994_/Q sky130_fd_sc_hd__dfxtp_1
X_5945_ _5951_/B _5951_/C _5945_/C vssd1 vssd1 vccd1 vccd1 _5952_/B sky130_fd_sc_hd__and3_1
Xclkbuf_1_1_0__2726_ clkbuf_0__2726_/X vssd1 vssd1 vccd1 vccd1 _5454__299/A sky130_fd_sc_hd__clkbuf_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4827_ _6504_/Q _6438_/Q _6536_/Q _6688_/Q _4701_/A _4806_/A vssd1 vssd1 vccd1 vccd1
+ _4827_/X sky130_fd_sc_hd__mux4_2
XFILLER_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4758_ _4691_/X input3/X _4695_/X _4757_/X vssd1 vssd1 vccd1 vccd1 _4758_/X sky130_fd_sc_hd__a22o_2
XFILLER_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3709_ _4458_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _3725_/S sky130_fd_sc_hd__or2_2
X_4689_ _4689_/A vssd1 vssd1 vccd1 vccd1 _4689_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6428_ _5910_/A _6424_/S _6427_/X _6430_/A vssd1 vssd1 vccd1 vccd1 _7094_/D sky130_fd_sc_hd__a211o_1
Xclkbuf_1_0_0__2873_ clkbuf_0__2873_/X vssd1 vssd1 vccd1 vccd1 _6084_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5168__229 _5168__229/A vssd1 vssd1 vccd1 vccd1 _6511_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3991_ _4572_/A _4123_/B vssd1 vssd1 vccd1 vccd1 _4007_/S sky130_fd_sc_hd__or2_2
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5730_ _7020_/Q _5734_/B vssd1 vssd1 vccd1 vccd1 _5731_/A sky130_fd_sc_hd__and2_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2511_ clkbuf_0__2511_/X vssd1 vssd1 vccd1 vccd1 _5130__198/A sky130_fd_sc_hd__clkbuf_4
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5661_ _7009_/Q _5609_/Y _5660_/X vssd1 vssd1 vccd1 vccd1 _5669_/C sky130_fd_sc_hd__o21ai_1
X_4612_ _3850_/X _6492_/Q _4618_/S vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__mux2_1
X_4543_ _4543_/A vssd1 vssd1 vccd1 vccd1 _6524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4474_ _4032_/X _6550_/Q _4474_/S vssd1 vssd1 vccd1 vccd1 _4475_/A sky130_fd_sc_hd__mux2_1
X_6213_ _6216_/A _6213_/B vssd1 vssd1 vccd1 vccd1 _6214_/C sky130_fd_sc_hd__or2_1
X_3425_ _3372_/X _7036_/Q _3429_/S vssd1 vssd1 vccd1 vccd1 _3426_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3356_ _7030_/Q vssd1 vssd1 vccd1 vccd1 _3764_/A sky130_fd_sc_hd__clkbuf_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_16 _4900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3287_ _7065_/Q _3263_/X _3291_/S vssd1 vssd1 vccd1 vccd1 _3288_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_38 _3877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_27 _3850_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_49 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _6435_/D sky130_fd_sc_hd__clkbuf_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6977_ _6977_/CLK _6977_/D vssd1 vssd1 vccd1 vccd1 _6977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5928_ _5929_/B _5926_/B _5927_/X _5406_/X vssd1 vssd1 vccd1 vccd1 _6868_/D sky130_fd_sc_hd__o211a_1
XFILLER_110_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2856_ clkbuf_0__2856_/X vssd1 vssd1 vccd1 vccd1 _5768__469/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4190_ _6684_/Q _4146_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4191_/A sky130_fd_sc_hd__mux2_1
X_3210_ _6732_/Q vssd1 vssd1 vccd1 vccd1 _5302_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6900_ _6900_/CLK _6900_/D vssd1 vssd1 vccd1 vccd1 _6900_/Q sky130_fd_sc_hd__dfxtp_1
X_6831_ _6831_/CLK _6831_/D vssd1 vssd1 vccd1 vccd1 _6831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6762_ _6762_/CLK _6762_/D vssd1 vssd1 vccd1 vccd1 _6762_/Q sky130_fd_sc_hd__dfxtp_1
X_3974_ _3974_/A _3978_/B vssd1 vssd1 vccd1 vccd1 _3975_/C sky130_fd_sc_hd__or2_1
XFILLER_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6693_ _6693_/CLK _6693_/D vssd1 vssd1 vccd1 vccd1 _6693_/Q sky130_fd_sc_hd__dfxtp_1
X_5644_ _5917_/B _5917_/C _7002_/Q vssd1 vssd1 vccd1 vccd1 _5657_/A sky130_fd_sc_hd__a21oi_1
X_6328__18 _6328__18/A vssd1 vssd1 vccd1 vccd1 _7038_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7089_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4526_ _4484_/X _6531_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4457_ _4457_/A vssd1 vssd1 vccd1 vccd1 _6558_/D sky130_fd_sc_hd__clkbuf_1
X_3408_ _3337_/X _7043_/Q _3410_/S vssd1 vssd1 vccd1 vccd1 _3409_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4388_ _3200_/X _6597_/Q _4396_/S vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__mux2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3339_/A vssd1 vssd1 vccd1 vccd1 _7059_/D sky130_fd_sc_hd__clkbuf_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5009_ _5009_/A vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6106__147 _6108__149/A vssd1 vssd1 vccd1 vccd1 _6955_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2839_ clkbuf_0__2839_/X vssd1 vssd1 vccd1 vccd1 _5718__446/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ _4017_/A vssd1 vssd1 vccd1 vccd1 _3690_/X sky130_fd_sc_hd__clkbuf_4
X_6030__86 _6033__89/A vssd1 vssd1 vccd1 vccd1 _6893_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5360_ _6673_/Q _6665_/Q _6657_/Q _6649_/Q _5330_/A _5312_/X vssd1 vssd1 vccd1 vccd1
+ _5360_/X sky130_fd_sc_hd__mux4_2
XFILLER_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5291_ _6954_/Q _6938_/Q _7063_/Q _6930_/Q _5290_/X _4069_/A vssd1 vssd1 vccd1 vccd1
+ _5291_/X sky130_fd_sc_hd__mux4_1
X_4311_ _4311_/A vssd1 vssd1 vccd1 vccd1 _6631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7030_ _7030_/CLK _7030_/D vssd1 vssd1 vccd1 vccd1 _7030_/Q sky130_fd_sc_hd__dfxtp_1
X_4242_ _4257_/S vssd1 vssd1 vccd1 vccd1 _4251_/S sky130_fd_sc_hd__buf_2
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4173_ _4173_/A vssd1 vssd1 vccd1 vccd1 _6692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6814_ _6814_/CLK _6814_/D vssd1 vssd1 vccd1 vccd1 _6814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2873_ _5852_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2873_/X sky130_fd_sc_hd__clkbuf_16
X_6745_ _7022_/CLK _6745_/D vssd1 vssd1 vccd1 vccd1 _6745_/Q sky130_fd_sc_hd__dfxtp_1
X_3957_ _4845_/A vssd1 vssd1 vccd1 vccd1 _3958_/A sky130_fd_sc_hd__buf_4
X_3888_ _3888_/A vssd1 vssd1 vccd1 vccd1 _6799_/D sky130_fd_sc_hd__clkbuf_1
X_6676_ _6676_/CLK _6676_/D vssd1 vssd1 vccd1 vccd1 _6676_/Q sky130_fd_sc_hd__dfxtp_1
X_5627_ _5892_/A _7006_/Q vssd1 vssd1 vccd1 vccd1 _6175_/A sky130_fd_sc_hd__xor2_2
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4509_ _4509_/A vssd1 vssd1 vccd1 vccd1 _6539_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7159_ _7159_/A vssd1 vssd1 vccd1 vccd1 _7159_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5518__350 _5519__351/A vssd1 vssd1 vccd1 vccd1 _6640_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4858_/X _6173_/A _4969_/A vssd1 vssd1 vccd1 vccd1 _4860_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3811_ _6827_/Q _3597_/X _3819_/S vssd1 vssd1 vccd1 vccd1 _3812_/A sky130_fd_sc_hd__mux2_1
X_5711__440 _5713__442/A vssd1 vssd1 vccd1 vccd1 _6734_/CLK sky130_fd_sc_hd__inv_2
X_6530_ _6530_/CLK _6530_/D vssd1 vssd1 vccd1 vccd1 _6530_/Q sky130_fd_sc_hd__dfxtp_1
X_4791_ _6760_/Q _6752_/Q _6715_/Q _6707_/Q _4807_/S _3959_/A vssd1 vssd1 vccd1 vccd1
+ _4791_/X sky130_fd_sc_hd__mux4_2
X_3742_ _3702_/X _6853_/Q _3744_/S vssd1 vssd1 vccd1 vccd1 _3743_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3673_ _3673_/A vssd1 vssd1 vccd1 vccd1 _6901_/D sky130_fd_sc_hd__clkbuf_1
X_6461_ _7089_/CLK _6461_/D vssd1 vssd1 vccd1 vccd1 _6461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6392_ _7138_/A _6170_/A _6401_/S vssd1 vssd1 vccd1 vccd1 _6393_/B sky130_fd_sc_hd__mux2_1
X_5412_ _6604_/Q _6588_/Q _6842_/Q _6826_/Q _5329_/X _5330_/X vssd1 vssd1 vccd1 vccd1
+ _5412_/X sky130_fd_sc_hd__mux4_1
Xoutput124 _7121_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[24] sky130_fd_sc_hd__buf_2
Xoutput113 _7111_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[14] sky130_fd_sc_hd__buf_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _5342_/X _5432_/S vssd1 vssd1 vccd1 vccd1 _5343_/X sky130_fd_sc_hd__and2b_1
Xoutput157 _7153_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[28] sky130_fd_sc_hd__buf_2
Xoutput146 _7143_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[18] sky130_fd_sc_hd__buf_2
Xoutput168 _7134_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[9] sky130_fd_sc_hd__buf_2
Xoutput135 _7106_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[9] sky130_fd_sc_hd__buf_2
X_6055__105 _6055__105/A vssd1 vssd1 vccd1 vccd1 _6913_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput179 _4979_/X vssd1 vssd1 vccd1 vccd1 wbs_data_o[12] sky130_fd_sc_hd__buf_2
X_5274_ _6734_/Q vssd1 vssd1 vccd1 vccd1 _5366_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_7013_ _7019_/CLK _7013_/D vssd1 vssd1 vccd1 vccd1 _7013_/Q sky130_fd_sc_hd__dfxtp_1
X_4225_ _3764_/X _6669_/Q _4233_/S vssd1 vssd1 vccd1 vccd1 _4226_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4156_ _6700_/Q _4155_/X _4156_/S vssd1 vssd1 vccd1 vccd1 _4157_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4087_ _4502_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4103_/S sky130_fd_sc_hd__or2_2
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2856_ _5763_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2856_/X sky130_fd_sc_hd__clkbuf_16
X_4989_ _4992_/A input11/X _4987_/X _7079_/Q vssd1 vssd1 vccd1 vccd1 _4989_/X sky130_fd_sc_hd__a22o_2
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6728_ _6728_/CLK _6728_/D vssd1 vssd1 vccd1 vccd1 _6728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6659_ _6659_/CLK _6659_/D vssd1 vssd1 vccd1 vccd1 _6659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput26 caravel_wb_data_i[30] vssd1 vssd1 vccd1 vccd1 _5016_/B sky130_fd_sc_hd__clkbuf_2
Xinput15 caravel_wb_data_i[20] vssd1 vssd1 vccd1 vccd1 _4995_/B sky130_fd_sc_hd__buf_4
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 _7107_/A sky130_fd_sc_hd__buf_4
Xinput59 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 _4682_/B sky130_fd_sc_hd__clkbuf_1
Xinput48 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 _7117_/A sky130_fd_sc_hd__buf_4
XFILLER_115_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6119__157 _6119__157/A vssd1 vssd1 vccd1 vccd1 _6965_/CLK sky130_fd_sc_hd__inv_2
XFILLER_96_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4010_ _4458_/A _4123_/B vssd1 vssd1 vccd1 vccd1 _4033_/S sky130_fd_sc_hd__or2_2
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5961_ _6875_/Q _6874_/Q _5961_/C vssd1 vssd1 vccd1 vccd1 _5968_/B sky130_fd_sc_hd__and3_1
XFILLER_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2742_ clkbuf_0__2742_/X vssd1 vssd1 vccd1 vccd1 _5534__363/A sky130_fd_sc_hd__clkbuf_4
X_4912_ _6857_/Q _6833_/Q _6809_/Q _6801_/Q _4701_/X _4806_/X vssd1 vssd1 vccd1 vccd1
+ _4913_/B sky130_fd_sc_hd__mux4_1
X_5892_ _5892_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5898_/C sky130_fd_sc_hd__nand2_1
X_4843_ _4804_/A _4842_/X _3953_/A vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4774_ _4808_/A vssd1 vssd1 vccd1 vccd1 _4774_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6513_ _6513_/CLK _6513_/D vssd1 vssd1 vccd1 vccd1 _6513_/Q sky130_fd_sc_hd__dfxtp_1
X_3725_ _3705_/X _6860_/Q _3725_/S vssd1 vssd1 vccd1 vccd1 _3726_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6444_ _7096_/CLK _6444_/D vssd1 vssd1 vccd1 vccd1 _6444_/Q sky130_fd_sc_hd__dfxtp_2
X_3656_ _3656_/A vssd1 vssd1 vccd1 vccd1 _6908_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3156_ clkbuf_0__3156_/X vssd1 vssd1 vccd1 vccd1 _6354__39/A sky130_fd_sc_hd__clkbuf_4
X_3587_ _6934_/Q _3450_/X _3589_/S vssd1 vssd1 vccd1 vccd1 _3588_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5326_ _6672_/Q _6664_/Q _6656_/Q _6648_/Q _5257_/X _5259_/X vssd1 vssd1 vccd1 vccd1
+ _5326_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5257_ _5337_/A vssd1 vssd1 vccd1 vccd1 _5257_/X sky130_fd_sc_hd__clkbuf_4
X_4208_ _4208_/A vssd1 vssd1 vccd1 vccd1 _6677_/D sky130_fd_sc_hd__clkbuf_1
X_5188_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__buf_1
XFILLER_68_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4139_ _6706_/Q _3895_/X _4139_/S vssd1 vssd1 vccd1 vccd1 _4140_/A sky130_fd_sc_hd__mux2_1
X_5718__446 _5718__446/A vssd1 vssd1 vccd1 vccd1 _6740_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2839_ _5716_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2839_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_22_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5805__496 _5806__497/A vssd1 vssd1 vccd1 vccd1 _6802_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3510_ _6968_/Q _3444_/X _3516_/S vssd1 vssd1 vccd1 vccd1 _3511_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4490_ _6744_/Q vssd1 vssd1 vccd1 vccd1 _4490_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__3010_ clkbuf_0__3010_/X vssd1 vssd1 vccd1 vccd1 _6096__139/A sky130_fd_sc_hd__clkbuf_4
XFILLER_109_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3441_ _3463_/S vssd1 vssd1 vccd1 vccd1 _3454_/S sky130_fd_sc_hd__buf_2
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6160_ _6155_/Y _7009_/Q _6156_/Y _4885_/X _6159_/X vssd1 vssd1 vccd1 vccd1 _6172_/A
+ sky130_fd_sc_hd__a221o_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3773_/A vssd1 vssd1 vccd1 vccd1 _3372_/X sky130_fd_sc_hd__buf_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _5929_/A _6868_/Q _5111_/C vssd1 vssd1 vccd1 vccd1 _5111_/X sky130_fd_sc_hd__or3_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6091_/X sky130_fd_sc_hd__buf_1
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5042_ _7080_/Q vssd1 vssd1 vccd1 vccd1 _6381_/A sky130_fd_sc_hd__inv_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6993_ _6993_/CLK _6993_/D vssd1 vssd1 vccd1 vccd1 _6993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5944_ _5966_/A vssd1 vssd1 vccd1 vccd1 _5944_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4826_ _4826_/A _4826_/B vssd1 vssd1 vccd1 vccd1 _4826_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4757_ _4856_/A _4753_/X _4987_/C _7096_/Q vssd1 vssd1 vccd1 vccd1 _4757_/X sky130_fd_sc_hd__a2bb2o_1
X_3708_ _3708_/A _4167_/B _4167_/A vssd1 vssd1 vccd1 vccd1 _4520_/B sky130_fd_sc_hd__or3b_4
X_4688_ input2/X _6444_/Q _4987_/A vssd1 vssd1 vccd1 vccd1 _4689_/A sky130_fd_sc_hd__mux2_2
X_6427_ _6427_/A _7127_/A _6427_/C vssd1 vssd1 vccd1 vccd1 _6427_/X sky130_fd_sc_hd__and3_1
Xclkbuf_1_0_0__2872_ clkbuf_0__2872_/X vssd1 vssd1 vccd1 vccd1 _5851__534/A sky130_fd_sc_hd__clkbuf_4
X_3639_ _3392_/X _6914_/Q _3639_/S vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5309_ _4071_/B _5308_/X _4071_/A vssd1 vssd1 vccd1 vccd1 _5309_/Y sky130_fd_sc_hd__o21ai_1
X_6289_ _7017_/Q _6292_/B vssd1 vssd1 vccd1 vccd1 _6289_/X sky130_fd_sc_hd__or2_1
XFILLER_102_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5497__334 _5497__334/A vssd1 vssd1 vccd1 vccd1 _6624_/CLK sky130_fd_sc_hd__inv_2
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5690__424 _5690__424/A vssd1 vssd1 vccd1 vccd1 _6718_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5770__470 _5773__473/A vssd1 vssd1 vccd1 vccd1 _6774_/CLK sky130_fd_sc_hd__inv_2
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3990_ _3727_/B _3990_/B _3990_/C vssd1 vssd1 vccd1 vccd1 _4123_/B sky130_fd_sc_hd__nand3b_4
Xclkbuf_1_1_0__2510_ clkbuf_0__2510_/X vssd1 vssd1 vccd1 vccd1 _5125__194/A sky130_fd_sc_hd__clkbuf_4
XFILLER_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5660_ _7008_/Q _5897_/B vssd1 vssd1 vccd1 vccd1 _5660_/X sky130_fd_sc_hd__xor2_1
XFILLER_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4611_ _4611_/A vssd1 vssd1 vccd1 vccd1 _6493_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5591_ _5591_/A vssd1 vssd1 vccd1 vccd1 _5591_/X sky130_fd_sc_hd__buf_1
X_4542_ _4481_/X _6524_/Q _4548_/S vssd1 vssd1 vccd1 vccd1 _4543_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4473_ _4473_/A vssd1 vssd1 vccd1 vccd1 _6551_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6212_ _6216_/A _6213_/B vssd1 vssd1 vccd1 vccd1 _6214_/B sky130_fd_sc_hd__nand2_1
X_3424_ _3424_/A vssd1 vssd1 vccd1 vccd1 _7037_/D sky130_fd_sc_hd__clkbuf_1
X_3355_ _3355_/A vssd1 vssd1 vccd1 vccd1 _7055_/D sky130_fd_sc_hd__clkbuf_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3286_ _3286_/A vssd1 vssd1 vccd1 vccd1 _7066_/D sky130_fd_sc_hd__clkbuf_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_39 _5723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XINSDIODE2_28 _3850_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5025_ _5025_/A _6425_/A _5025_/C vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__and3_1
XINSDIODE2_17 _5342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6976_ _6976_/CLK _6976_/D vssd1 vssd1 vccd1 vccd1 _6976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5927_ _6015_/B _5953_/B _6868_/Q _5250_/A vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4809_ _4851_/S vssd1 vssd1 vccd1 vccd1 _4957_/S sky130_fd_sc_hd__buf_4
XFILLER_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2855_ clkbuf_0__2855_/X vssd1 vssd1 vccd1 vccd1 _5762__464/A sky130_fd_sc_hd__clkbuf_4
X_5208__260 _5210__262/A vssd1 vssd1 vccd1 vccd1 _6542_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5880__76 _5883__79/A vssd1 vssd1 vccd1 vccd1 _6862_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5174__234 _5174__234/A vssd1 vssd1 vccd1 vccd1 _6516_/CLK sky130_fd_sc_hd__inv_2
X_6042__95 _6043__96/A vssd1 vssd1 vccd1 vccd1 _6903_/CLK sky130_fd_sc_hd__inv_2
X_5512__345 _5514__347/A vssd1 vssd1 vccd1 vccd1 _6635_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6360__44 _6360__44/A vssd1 vssd1 vccd1 vccd1 _7064_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5593__406 _5596__409/A vssd1 vssd1 vccd1 vccd1 _6699_/CLK sky130_fd_sc_hd__inv_2
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6830_ _6830_/CLK _6830_/D vssd1 vssd1 vccd1 vccd1 _6830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6761_ _6761_/CLK _6761_/D vssd1 vssd1 vccd1 vccd1 _6761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _3951_/Y _3975_/B _3972_/X vssd1 vssd1 vccd1 vccd1 _6771_/D sky130_fd_sc_hd__a21oi_1
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6692_ _6692_/CLK _6692_/D vssd1 vssd1 vccd1 vccd1 _6692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5643_ _5913_/A _5913_/B _6167_/A vssd1 vssd1 vccd1 vccd1 _5917_/C sky130_fd_sc_hd__o21ai_2
XFILLER_117_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4525_ _4525_/A vssd1 vssd1 vccd1 vccd1 _6532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4456_ _4032_/X _6558_/Q _4456_/S vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__mux2_1
X_3407_ _3407_/A vssd1 vssd1 vccd1 vccd1 _7044_/D sky130_fd_sc_hd__clkbuf_1
X_4387_ _4402_/S vssd1 vssd1 vccd1 vccd1 _4396_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3338_ _3337_/X _7059_/Q _3342_/S vssd1 vssd1 vccd1 vccd1 _3339_/A sky130_fd_sc_hd__mux2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3269_ _7023_/Q vssd1 vssd1 vccd1 vccd1 _3269_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5008_ _5014_/A _5008_/B vssd1 vssd1 vccd1 vccd1 _5009_/A sky130_fd_sc_hd__and2_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6959_ _6959_/CLK _6959_/D vssd1 vssd1 vccd1 vccd1 _6959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2838_ clkbuf_0__2838_/X vssd1 vssd1 vccd1 vccd1 _5715__444/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6333__22 _6335__24/A vssd1 vssd1 vccd1 vccd1 _7042_/CLK sky130_fd_sc_hd__inv_2
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5290_ _5329_/A vssd1 vssd1 vccd1 vccd1 _5290_/X sky130_fd_sc_hd__clkbuf_8
X_4310_ _3785_/X _6631_/Q _4312_/S vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4241_ _4404_/A _4259_/B vssd1 vssd1 vccd1 vccd1 _4257_/S sky130_fd_sc_hd__or2_2
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4172_ _4014_/X _6692_/Q _4178_/S vssd1 vssd1 vccd1 vccd1 _4173_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2872_ _5846_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2872_/X sky130_fd_sc_hd__clkbuf_16
X_6813_ _6813_/CLK _6813_/D vssd1 vssd1 vccd1 vccd1 _6813_/Q sky130_fd_sc_hd__dfxtp_1
X_6744_ _7022_/CLK _6744_/D vssd1 vssd1 vccd1 vccd1 _6744_/Q sky130_fd_sc_hd__dfxtp_1
X_3956_ _6768_/Q vssd1 vssd1 vccd1 vccd1 _4845_/A sky130_fd_sc_hd__buf_4
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6675_ _6675_/CLK _6675_/D vssd1 vssd1 vccd1 vccd1 _6675_/Q sky130_fd_sc_hd__dfxtp_1
X_3887_ _6799_/Q _3886_/X _3887_/S vssd1 vssd1 vccd1 vccd1 _3888_/A sky130_fd_sc_hd__mux2_1
X_5626_ _7003_/Q _5895_/B vssd1 vssd1 vccd1 vccd1 _5626_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4508_ _4484_/X _6539_/Q _4512_/S vssd1 vssd1 vccd1 vccd1 _4509_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4439_ _4439_/A vssd1 vssd1 vccd1 vccd1 _6566_/D sky130_fd_sc_hd__clkbuf_1
X_7158_ _7158_/A vssd1 vssd1 vccd1 vccd1 _7158_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7089_ _7089_/CLK _7089_/D vssd1 vssd1 vccd1 vccd1 _7089_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6109_/X sky130_fd_sc_hd__buf_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6112__152 _6113__153/A vssd1 vssd1 vccd1 vccd1 _6960_/CLK sky130_fd_sc_hd__inv_2
XFILLER_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2836_ clkbuf_0__2836_/X vssd1 vssd1 vccd1 vccd1 _5750_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_2_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4790_ _4954_/S _4790_/B vssd1 vssd1 vccd1 vccd1 _4790_/Y sky130_fd_sc_hd__nor2_1
X_3810_ _3825_/S vssd1 vssd1 vccd1 vccd1 _3819_/S sky130_fd_sc_hd__buf_2
XFILLER_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3741_ _3741_/A vssd1 vssd1 vccd1 vccd1 _6854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _3341_/X _6901_/Q _3672_/S vssd1 vssd1 vccd1 vccd1 _3673_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6460_ _7089_/CLK _6460_/D vssd1 vssd1 vccd1 vccd1 _6460_/Q sky130_fd_sc_hd__dfxtp_1
X_6391_ _6391_/A vssd1 vssd1 vccd1 vccd1 _6408_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5411_ _6644_/Q _6636_/Q _6620_/Q _6612_/Q _4083_/A _4063_/A vssd1 vssd1 vccd1 vccd1
+ _5411_/X sky130_fd_sc_hd__mux4_1
Xoutput125 _7122_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput114 _7112_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[15] sky130_fd_sc_hd__buf_2
X_5342_ _6924_/Q _6916_/Q _7033_/Q _7049_/Q _4066_/A _5341_/X vssd1 vssd1 vccd1 vccd1
+ _5342_/X sky130_fd_sc_hd__mux4_2
X_5187__244 _5187__244/A vssd1 vssd1 vccd1 vccd1 _6526_/CLK sky130_fd_sc_hd__inv_2
Xoutput136 _4685_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_cyc_o sky130_fd_sc_hd__buf_2
Xoutput158 _7154_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[29] sky130_fd_sc_hd__buf_2
Xoutput147 _7144_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput169 _7157_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_sel_o[0] sky130_fd_sc_hd__buf_2
XFILLER_114_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7012_ _7019_/CLK _7012_/D vssd1 vssd1 vccd1 vccd1 _7012_/Q sky130_fd_sc_hd__dfxtp_1
X_5273_ _5262_/X _5271_/X _5394_/S vssd1 vssd1 vccd1 vccd1 _5273_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4224_ _4239_/S vssd1 vssd1 vccd1 vccd1 _4233_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4155_ _7026_/Q vssd1 vssd1 vccd1 vccd1 _4155_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4086_ _4086_/A vssd1 vssd1 vccd1 vccd1 _6730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5491__329 _5491__329/A vssd1 vssd1 vccd1 vccd1 _6619_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__2855_ _5757_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2855_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4988_ _4992_/A input10/X _4987_/X _7080_/Q vssd1 vssd1 vccd1 vccd1 _4988_/X sky130_fd_sc_hd__a22o_2
XFILLER_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6727_ _6727_/CLK _6727_/D vssd1 vssd1 vccd1 vccd1 _6727_/Q sky130_fd_sc_hd__dfxtp_1
X_3939_ _4570_/S vssd1 vssd1 vccd1 vccd1 _4562_/S sky130_fd_sc_hd__buf_2
X_6658_ _6658_/CLK _6658_/D vssd1 vssd1 vccd1 vccd1 _6658_/Q sky130_fd_sc_hd__dfxtp_1
X_5609_ _6155_/A _5609_/B vssd1 vssd1 vccd1 vccd1 _5609_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_117_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6589_ _6589_/CLK _6589_/D vssd1 vssd1 vccd1 vccd1 _6589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 caravel_wb_data_i[31] vssd1 vssd1 vccd1 vccd1 _5018_/B sky130_fd_sc_hd__buf_2
Xinput16 caravel_wb_data_i[21] vssd1 vssd1 vccd1 vccd1 _4997_/B sky130_fd_sc_hd__buf_4
Xinput38 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 _7108_/A sky130_fd_sc_hd__buf_4
Xinput49 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 _7118_/A sky130_fd_sc_hd__buf_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5960_ _6874_/Q _5961_/C _6875_/Q vssd1 vssd1 vccd1 vccd1 _5962_/A sky130_fd_sc_hd__a21oi_1
XFILLER_18_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2741_ clkbuf_0__2741_/X vssd1 vssd1 vccd1 vccd1 _5554_/A sky130_fd_sc_hd__clkbuf_4
X_4911_ _4944_/A _4910_/X _4782_/X vssd1 vssd1 vccd1 vccd1 _4911_/Y sky130_fd_sc_hd__o21ai_1
X_5891_ _6878_/Q _5891_/B vssd1 vssd1 vccd1 vccd1 _5891_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4842_ _6545_/Q _6725_/Q _6863_/Q _6529_/Q _4719_/A _4898_/A vssd1 vssd1 vccd1 vccd1
+ _4842_/X sky130_fd_sc_hd__mux4_2
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ _6768_/Q vssd1 vssd1 vccd1 vccd1 _4808_/A sky130_fd_sc_hd__inv_2
X_6061__110 _6064__113/A vssd1 vssd1 vccd1 vccd1 _6918_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ _3724_/A vssd1 vssd1 vccd1 vccd1 _6861_/D sky130_fd_sc_hd__clkbuf_1
X_6512_ _6512_/CLK _6512_/D vssd1 vssd1 vccd1 vccd1 _6512_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6443_ _6443_/CLK _6443_/D vssd1 vssd1 vccd1 vccd1 _6443_/Q sky130_fd_sc_hd__dfxtp_1
X_3655_ _3345_/X _6908_/Q _3659_/S vssd1 vssd1 vccd1 vccd1 _3656_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0__3155_ clkbuf_0__3155_/X vssd1 vssd1 vccd1 vccd1 _6348__34/A sky130_fd_sc_hd__clkbuf_4
X_3586_ _3586_/A vssd1 vssd1 vccd1 vccd1 _6935_/D sky130_fd_sc_hd__clkbuf_1
X_5325_ _7073_/Q _6699_/Q _6568_/Q _6846_/Q _5251_/X _5254_/X vssd1 vssd1 vccd1 vccd1
+ _5325_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5256_ _6730_/Q vssd1 vssd1 vccd1 vccd1 _5337_/A sky130_fd_sc_hd__clkbuf_4
X_4207_ _6677_/Q _4141_/X _4215_/S vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4138_ _4138_/A vssd1 vssd1 vccd1 vccd1 _6707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4069_ _4069_/A _6750_/Q _5739_/C vssd1 vssd1 vccd1 vccd1 _4070_/B sky130_fd_sc_hd__and3_1
XFILLER_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2838_ _5710_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2838_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125__162 _6127__164/A vssd1 vssd1 vccd1 vccd1 _6970_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3440_ _4186_/A _3898_/B vssd1 vssd1 vccd1 vccd1 _3463_/S sky130_fd_sc_hd__nor2_4
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3371_ _7028_/Q vssd1 vssd1 vccd1 vccd1 _3773_/A sky130_fd_sc_hd__clkbuf_4
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5110_ _5108_/X _5109_/X _6888_/Q vssd1 vssd1 vccd1 vccd1 _5111_/C sky130_fd_sc_hd__mux2_1
XFILLER_57_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5041_ _6469_/Q _6468_/Q vssd1 vssd1 vccd1 vccd1 _6377_/A sky130_fd_sc_hd__or2b_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6992_ _6992_/CLK _6992_/D vssd1 vssd1 vccd1 vccd1 _6992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5943_ _5941_/Y _5938_/X _5942_/X _5972_/A vssd1 vssd1 vccd1 vccd1 _6871_/D sky130_fd_sc_hd__o211a_1
XFILLER_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4825_ _6854_/Q _6830_/Q _6806_/Q _6798_/Q _4891_/B _4709_/X vssd1 vssd1 vccd1 vccd1
+ _4826_/B sky130_fd_sc_hd__mux4_2
XFILLER_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4756_ _4969_/A vssd1 vssd1 vccd1 vccd1 _4987_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4687_ _4687_/A vssd1 vssd1 vccd1 vccd1 _4687_/X sky130_fd_sc_hd__clkbuf_1
X_3707_ _3707_/A vssd1 vssd1 vccd1 vccd1 _6889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2871_ clkbuf_0__2871_/X vssd1 vssd1 vccd1 vccd1 _5843__527/A sky130_fd_sc_hd__clkbuf_4
X_6426_ _6426_/A vssd1 vssd1 vccd1 vccd1 _7093_/D sky130_fd_sc_hd__clkbuf_1
X_3638_ _3638_/A vssd1 vssd1 vccd1 vccd1 _6915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3569_ _3376_/X _6942_/Q _3571_/S vssd1 vssd1 vccd1 vccd1 _3570_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5308_ _6955_/Q _6939_/Q _7064_/Q _6931_/Q _5282_/X _4083_/X vssd1 vssd1 vccd1 vccd1
+ _5308_/X sky130_fd_sc_hd__mux4_1
X_6288_ _7017_/Q _6284_/X _6287_/X _6192_/X vssd1 vssd1 vccd1 vccd1 _7016_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5239_ _5449_/A vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__buf_1
XFILLER_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6068__116 _6069__117/A vssd1 vssd1 vccd1 vccd1 _6924_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2518_ clkbuf_0__2518_/X vssd1 vssd1 vccd1 vccd1 _5166__227/A sky130_fd_sc_hd__clkbuf_16
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4610_ _3845_/X _6493_/Q _4618_/S vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4541_ _4541_/A vssd1 vssd1 vccd1 vccd1 _6525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4472_ _4029_/X _6551_/Q _4474_/S vssd1 vssd1 vccd1 vccd1 _4473_/A sky130_fd_sc_hd__mux2_1
X_6211_ _6211_/A vssd1 vssd1 vccd1 vccd1 _6998_/D sky130_fd_sc_hd__clkbuf_1
X_3423_ _3368_/X _7037_/Q _3429_/S vssd1 vssd1 vccd1 vccd1 _3424_/A sky130_fd_sc_hd__mux2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3354_ _3353_/X _7055_/Q _3354_/S vssd1 vssd1 vccd1 vccd1 _3355_/A sky130_fd_sc_hd__mux2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _7066_/Q _3260_/X _3285_/S vssd1 vssd1 vccd1 vccd1 _3286_/A sky130_fd_sc_hd__mux2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XINSDIODE2_29 _3853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XINSDIODE2_18 _5434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5024_ _4683_/B _4683_/C _4683_/D _5023_/X _4987_/A vssd1 vssd1 vccd1 vccd1 _5025_/C
+ sky130_fd_sc_hd__a41o_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6975_ _6975_/CLK _6975_/D vssd1 vssd1 vccd1 vccd1 _6975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5926_ _6013_/B _5926_/B vssd1 vssd1 vccd1 vccd1 _5953_/B sky130_fd_sc_hd__nand2_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4808_ _4808_/A vssd1 vssd1 vccd1 vccd1 _4808_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4739_ _6468_/Q _6469_/Q vssd1 vssd1 vccd1 vccd1 _4750_/A sky130_fd_sc_hd__or2b_1
XFILLER_119_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6409_ _6409_/A vssd1 vssd1 vccd1 vccd1 _7088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2854_ clkbuf_0__2854_/X vssd1 vssd1 vccd1 vccd1 _5784_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6345__31 _6347__33/A vssd1 vssd1 vccd1 vccd1 _7051_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5181__239 _5181__239/A vssd1 vssd1 vccd1 vccd1 _6521_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6760_ _6760_/CLK _6760_/D vssd1 vssd1 vccd1 vccd1 _6760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3972_ _3971_/X _3974_/A _3978_/B _3936_/A vssd1 vssd1 vccd1 vccd1 _3972_/X sky130_fd_sc_hd__a31o_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6691_ _6691_/CLK _6691_/D vssd1 vssd1 vccd1 vccd1 _6691_/Q sky130_fd_sc_hd__dfxtp_1
X_5642_ _5642_/A _5642_/B _5642_/C _5642_/D vssd1 vssd1 vccd1 vccd1 _5642_/X sky130_fd_sc_hd__or4_1
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5573_ _5573_/A vssd1 vssd1 vccd1 vccd1 _5573_/X sky130_fd_sc_hd__buf_1
X_4524_ _4481_/X _6532_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4455_ _4455_/A vssd1 vssd1 vccd1 vccd1 _6559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3406_ _3333_/X _7044_/Q _3410_/S vssd1 vssd1 vccd1 vccd1 _3407_/A sky130_fd_sc_hd__mux2_1
X_4386_ _4404_/A _4386_/B vssd1 vssd1 vccd1 vccd1 _4402_/S sky130_fd_sc_hd__or2_2
X_3337_ _4020_/A vssd1 vssd1 vccd1 vccd1 _3337_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_98_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3268_/A vssd1 vssd1 vccd1 vccd1 _7072_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5007_ _5007_/A vssd1 vssd1 vccd1 vccd1 _5007_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5574__395 _5577__398/A vssd1 vssd1 vccd1 vccd1 _6685_/CLK sky130_fd_sc_hd__inv_2
X_6958_ _6958_/CLK _6958_/D vssd1 vssd1 vccd1 vccd1 _6958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6889_ _6889_/CLK _6889_/D vssd1 vssd1 vccd1 vccd1 _6889_/Q sky130_fd_sc_hd__dfxtp_1
X_5909_ _5917_/B _5917_/C _6876_/Q vssd1 vssd1 vccd1 vccd1 _5912_/C sky130_fd_sc_hd__a21oi_1
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2837_ clkbuf_0__2837_/X vssd1 vssd1 vccd1 vccd1 _5709__439/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4240_ _4240_/A vssd1 vssd1 vccd1 vccd1 _6662_/D sky130_fd_sc_hd__clkbuf_1
X_4171_ _4171_/A vssd1 vssd1 vccd1 vccd1 _6693_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6812_ _6812_/CLK _6812_/D vssd1 vssd1 vccd1 vccd1 _6812_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__2871_ _5840_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2871_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6743_ _7093_/CLK _6743_/D vssd1 vssd1 vccd1 vccd1 _6743_/Q sky130_fd_sc_hd__dfxtp_2
X_3955_ _4804_/A vssd1 vssd1 vccd1 vccd1 _3968_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6674_ _6674_/CLK _6674_/D vssd1 vssd1 vccd1 vccd1 _6674_/Q sky130_fd_sc_hd__dfxtp_1
X_3886_ _6744_/Q vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__buf_2
X_5625_ _6168_/A _5917_/B _5890_/B vssd1 vssd1 vccd1 vccd1 _5895_/B sky130_fd_sc_hd__a21oi_4
XFILLER_117_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4507_ _4507_/A vssd1 vssd1 vccd1 vccd1 _6540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4438_ _3269_/X _6566_/Q _4438_/S vssd1 vssd1 vccd1 vccd1 _4439_/A sky130_fd_sc_hd__mux2_1
X_7157_ _7157_/A vssd1 vssd1 vccd1 vccd1 _7157_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4369_ _4384_/S vssd1 vssd1 vccd1 vccd1 _4378_/S sky130_fd_sc_hd__buf_2
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7088_ _7089_/CLK _7088_/D vssd1 vssd1 vccd1 vccd1 _7088_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5810__500 _5813__503/A vssd1 vssd1 vccd1 vccd1 _6806_/CLK sky130_fd_sc_hd__inv_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3740_ _3699_/X _6854_/Q _3744_/S vssd1 vssd1 vccd1 vccd1 _3741_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3671_ _3671_/A vssd1 vssd1 vccd1 vccd1 _6902_/D sky130_fd_sc_hd__clkbuf_1
X_6390_ _6390_/A vssd1 vssd1 vccd1 vccd1 _7082_/D sky130_fd_sc_hd__clkbuf_1
X_5410_ _5408_/X _5409_/X _5410_/S vssd1 vssd1 vccd1 vccd1 _5410_/X sky130_fd_sc_hd__mux2_1
Xoutput115 _7113_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[16] sky130_fd_sc_hd__buf_2
X_5341_ _5341_/A vssd1 vssd1 vccd1 vccd1 _5341_/X sky130_fd_sc_hd__buf_2
Xoutput126 _7123_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput159 _7127_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[2] sky130_fd_sc_hd__buf_2
Xoutput148 _7126_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput137 _7125_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[0] sky130_fd_sc_hd__buf_2
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7011_ _7011_/CLK _7011_/D vssd1 vssd1 vccd1 vccd1 _7011_/Q sky130_fd_sc_hd__dfxtp_1
X_5272_ _5334_/A vssd1 vssd1 vccd1 vccd1 _5394_/S sky130_fd_sc_hd__clkbuf_4
X_5525__356 _5527__358/A vssd1 vssd1 vccd1 vccd1 _6646_/CLK sky130_fd_sc_hd__inv_2
X_4223_ _4296_/A _4259_/B vssd1 vssd1 vccd1 vccd1 _4239_/S sky130_fd_sc_hd__or2_2
X_4154_ _4154_/A vssd1 vssd1 vccd1 vccd1 _6701_/D sky130_fd_sc_hd__clkbuf_1
X_4085_ _4070_/B _4085_/B _6318_/B vssd1 vssd1 vccd1 vccd1 _4086_/A sky130_fd_sc_hd__and3b_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2854_ _5756_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2854_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6726_ _6726_/CLK _6726_/D vssd1 vssd1 vccd1 vccd1 _6726_/Q sky130_fd_sc_hd__dfxtp_1
X_4987_ _4987_/A _6696_/Q _4987_/C vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__and3_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3938_ _4168_/A _4590_/B vssd1 vssd1 vccd1 vccd1 _4570_/S sky130_fd_sc_hd__nor2_2
X_3869_ _6804_/Q _3868_/X _3869_/S vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__mux2_1
X_6657_ _6657_/CLK _6657_/D vssd1 vssd1 vccd1 vccd1 _6657_/Q sky130_fd_sc_hd__dfxtp_1
X_5608_ _6170_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _5609_/B sky130_fd_sc_hd__nor2_1
X_6588_ _6588_/CLK _6588_/D vssd1 vssd1 vccd1 vccd1 _6588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 caravel_wb_data_i[22] vssd1 vssd1 vccd1 vccd1 _4999_/B sky130_fd_sc_hd__buf_4
Xinput28 caravel_wb_data_i[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0__3019_ clkbuf_0__3019_/X vssd1 vssd1 vccd1 vccd1 _6143__177/A sky130_fd_sc_hd__clkbuf_4
Xinput39 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 _7109_/A sky130_fd_sc_hd__buf_4
XFILLER_108_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5817__506 _5820__509/A vssd1 vssd1 vccd1 vccd1 _6812_/CLK sky130_fd_sc_hd__inv_2
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0__2740_ clkbuf_0__2740_/X vssd1 vssd1 vccd1 vccd1 _5527__358/A sky130_fd_sc_hd__clkbuf_4
X_4910_ _6764_/Q _6756_/Q _6719_/Q _6711_/Q _4956_/S _3959_/A vssd1 vssd1 vccd1 vccd1
+ _4910_/X sky130_fd_sc_hd__mux4_2
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5890_ _5890_/A _5890_/B vssd1 vssd1 vccd1 vccd1 _5891_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4841_ _4806_/X _4838_/X _4840_/X vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__a21o_1
X_4772_ _7040_/Q _6971_/Q _4772_/S vssd1 vssd1 vccd1 vccd1 _4772_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5531__360 _5534__363/A vssd1 vssd1 vccd1 vccd1 _6650_/CLK sky130_fd_sc_hd__inv_2
X_3723_ _3702_/X _6861_/Q _3725_/S vssd1 vssd1 vccd1 vccd1 _3724_/A sky130_fd_sc_hd__mux2_1
X_6511_ _6511_/CLK _6511_/D vssd1 vssd1 vccd1 vccd1 _6511_/Q sky130_fd_sc_hd__dfxtp_1
X_6442_ _6442_/CLK _6442_/D vssd1 vssd1 vccd1 vccd1 _6442_/Q sky130_fd_sc_hd__dfxtp_1
X_3654_ _3654_/A vssd1 vssd1 vccd1 vccd1 _6909_/D sky130_fd_sc_hd__clkbuf_1
X_3585_ _6935_/Q _3447_/X _3589_/S vssd1 vssd1 vccd1 vccd1 _3586_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5324_ _5324_/A vssd1 vssd1 vccd1 vccd1 _5324_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5255_ _7071_/Q _6697_/Q _6566_/Q _6844_/Q _5251_/X _5254_/X vssd1 vssd1 vccd1 vccd1
+ _5255_/X sky130_fd_sc_hd__mux4_2
XFILLER_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4206_ _4221_/S vssd1 vssd1 vccd1 vccd1 _4215_/S sky130_fd_sc_hd__buf_2
XFILLER_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4137_ _6707_/Q _3892_/X _4139_/S vssd1 vssd1 vccd1 vccd1 _4138_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4068_ _4068_/A _4068_/B _4068_/C _4068_/D vssd1 vssd1 vccd1 vccd1 _5739_/C sky130_fd_sc_hd__or4_4
X_5202__256 _5202__256/A vssd1 vssd1 vccd1 vccd1 _6538_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2869_ clkbuf_0__2869_/X vssd1 vssd1 vccd1 vccd1 _5831__517/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2837_ _5704_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2837_/X sky130_fd_sc_hd__clkbuf_16
X_6709_ _6709_/CLK _6709_/D vssd1 vssd1 vccd1 vccd1 _6709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2519_ clkbuf_0__2519_/X vssd1 vssd1 vccd1 vccd1 _5172__232/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5823__510 _5825__512/A vssd1 vssd1 vccd1 vccd1 _6816_/CLK sky130_fd_sc_hd__inv_2
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3370_ _3370_/A vssd1 vssd1 vccd1 vccd1 _7053_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6991_ _6991_/CLK _6991_/D vssd1 vssd1 vccd1 vccd1 _6991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5942_ _5945_/C _6013_/B _5926_/B _5951_/C vssd1 vssd1 vccd1 vccd1 _5942_/X sky130_fd_sc_hd__a31o_1
X_4824_ _4716_/A _4823_/X _4711_/X vssd1 vssd1 vccd1 vccd1 _4824_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4755_ _4798_/A _6377_/B vssd1 vssd1 vccd1 vccd1 _4969_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ _3705_/X _6889_/Q _3706_/S vssd1 vssd1 vccd1 vccd1 _3707_/A sky130_fd_sc_hd__mux2_1
X_4686_ _5050_/C _4686_/B vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__and2_2
X_6425_ _6425_/A _6425_/B vssd1 vssd1 vccd1 vccd1 _6426_/A sky130_fd_sc_hd__and2_1
X_3637_ _3388_/X _6915_/Q _3639_/S vssd1 vssd1 vccd1 vccd1 _3638_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__2870_ clkbuf_0__2870_/X vssd1 vssd1 vccd1 vccd1 _5836__521/A sky130_fd_sc_hd__clkbuf_4
X_3568_ _3568_/A vssd1 vssd1 vccd1 vccd1 _6943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5307_ _5306_/X _5355_/B vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__and2b_1
X_6287_ _7016_/Q _6292_/B vssd1 vssd1 vccd1 vccd1 _6287_/X sky130_fd_sc_hd__or2_1
XFILLER_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3499_ _3345_/X _6972_/Q _3503_/S vssd1 vssd1 vccd1 vccd1 _3500_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5238_ _5560_/A vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__buf_1
X_5169_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__buf_1
XFILLER_68_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5538__366 _5538__366/A vssd1 vssd1 vccd1 vccd1 _6656_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6372__54 _6372__54/A vssd1 vssd1 vccd1 vccd1 _7074_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2999_ clkbuf_0__2999_/X vssd1 vssd1 vccd1 vccd1 _6038__92/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5747__452 _5747__452/A vssd1 vssd1 vccd1 vccd1 _6756_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4540_ _4476_/X _6525_/Q _4548_/S vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4471_ _4471_/A vssd1 vssd1 vccd1 vccd1 _6552_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6210_ _6213_/B _6210_/B _6229_/C vssd1 vssd1 vccd1 vccd1 _6211_/A sky130_fd_sc_hd__and3b_1
X_3422_ _3422_/A vssd1 vssd1 vccd1 vccd1 _7038_/D sky130_fd_sc_hd__clkbuf_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _4032_/A vssd1 vssd1 vccd1 vccd1 _3353_/X sky130_fd_sc_hd__clkbuf_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3284_ _3284_/A vssd1 vssd1 vccd1 vccd1 _7067_/D sky130_fd_sc_hd__clkbuf_1
X_6072_ _6072_/A vssd1 vssd1 vccd1 vccd1 _6072_/X sky130_fd_sc_hd__buf_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_19 _7090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _7122_/A _7121_/A _7124_/A _7123_/A vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__and4_1
XFILLER_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6974_ _6974_/CLK _6974_/D vssd1 vssd1 vccd1 vccd1 _6974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5925_ _6869_/Q _6868_/Q vssd1 vssd1 vccd1 vccd1 _6013_/B sky130_fd_sc_hd__or2_2
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4807_ _7041_/Q _6972_/Q _4807_/S vssd1 vssd1 vccd1 vccd1 _4807_/X sky130_fd_sc_hd__mux2_2
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4738_ _4726_/X _4733_/X _4737_/X _4904_/A vssd1 vssd1 vccd1 vccd1 _4738_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4669_ _4669_/A vssd1 vssd1 vccd1 vccd1 _6441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6408_ _6408_/A _6408_/B vssd1 vssd1 vccd1 vccd1 _6409_/A sky130_fd_sc_hd__and2_1
XFILLER_115_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2853_ clkbuf_0__2853_/X vssd1 vssd1 vccd1 vccd1 _5752__456/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6074__121 _6075__122/A vssd1 vssd1 vccd1 vccd1 _6929_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5865__64 _5865__64/A vssd1 vssd1 vccd1 vccd1 _6850_/CLK sky130_fd_sc_hd__inv_2
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3019_ _6140_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3019_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5215__266 _5216__267/A vssd1 vssd1 vccd1 vccd1 _6548_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3971_ _4724_/A vssd1 vssd1 vccd1 vccd1 _3971_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5710_ _5716_/A vssd1 vssd1 vccd1 vccd1 _5710_/X sky130_fd_sc_hd__buf_1
X_6690_ _6690_/CLK _6690_/D vssd1 vssd1 vccd1 vccd1 _6690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5641_ _6999_/Q _5908_/B _5637_/X _5638_/Y _5640_/Y vssd1 vssd1 vccd1 vccd1 _5642_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4523_ _4523_/A vssd1 vssd1 vccd1 vccd1 _6533_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4454_ _4029_/X _6559_/Q _4456_/S vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__mux2_1
X_3405_ _3405_/A vssd1 vssd1 vccd1 vccd1 _7045_/D sky130_fd_sc_hd__clkbuf_1
X_4385_ _4385_/A vssd1 vssd1 vccd1 vccd1 _6598_/D sky130_fd_sc_hd__clkbuf_1
X_6138__173 _6139__174/A vssd1 vssd1 vccd1 vccd1 _6981_/CLK sky130_fd_sc_hd__inv_2
X_3336_ _6745_/Q vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5006_ _5014_/A _5006_/B vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__and2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _7072_/Q _3266_/X _3270_/S vssd1 vssd1 vccd1 vccd1 _3268_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6957_ _6957_/CLK _6957_/D vssd1 vssd1 vccd1 vccd1 _6957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5908_ _6873_/Q _5908_/B vssd1 vssd1 vccd1 vccd1 _5912_/B sky130_fd_sc_hd__xnor2_1
X_6888_ _6888_/CLK _6888_/D vssd1 vssd1 vccd1 vccd1 _6888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2519_ _5169_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2519_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_1_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5035__184 _5035__184/A vssd1 vssd1 vccd1 vccd1 _6440_/CLK sky130_fd_sc_hd__inv_2
XFILLER_114_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4170_ _4009_/X _6693_/Q _4178_/S vssd1 vssd1 vccd1 vccd1 _4171_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6811_ _6811_/CLK _6811_/D vssd1 vssd1 vccd1 vccd1 _6811_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2870_ _5834_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2870_/X sky130_fd_sc_hd__clkbuf_16
X_6742_ _7022_/CLK _6742_/D vssd1 vssd1 vccd1 vccd1 _6742_/Q sky130_fd_sc_hd__dfxtp_2
X_3954_ _6769_/Q vssd1 vssd1 vccd1 vccd1 _4804_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3885_ _3885_/A vssd1 vssd1 vccd1 vccd1 _6800_/D sky130_fd_sc_hd__clkbuf_1
X_6673_ _6673_/CLK _6673_/D vssd1 vssd1 vccd1 vccd1 _6673_/Q sky130_fd_sc_hd__dfxtp_1
X_5624_ _6167_/A _5664_/A _5913_/B vssd1 vssd1 vccd1 vccd1 _5917_/B sky130_fd_sc_hd__or3_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4506_ _4481_/X _6540_/Q _4512_/S vssd1 vssd1 vccd1 vccd1 _4507_/A sky130_fd_sc_hd__mux2_1
X_5486_ _5486_/A vssd1 vssd1 vccd1 vccd1 _5486_/X sky130_fd_sc_hd__buf_1
XFILLER_104_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4437_ _4437_/A vssd1 vssd1 vccd1 vccd1 _6567_/D sky130_fd_sc_hd__clkbuf_1
X_7156_ _7156_/A vssd1 vssd1 vccd1 vccd1 _7156_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _4368_/A _4404_/B vssd1 vssd1 vccd1 vccd1 _4384_/S sky130_fd_sc_hd__nor2_2
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3319_ _6778_/Q _4765_/A vssd1 vssd1 vccd1 vccd1 _3484_/A sky130_fd_sc_hd__and2_1
X_7087_ _7095_/CLK _7087_/D vssd1 vssd1 vccd1 vccd1 _7087_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4299_/A vssd1 vssd1 vccd1 vccd1 _6637_/D sky130_fd_sc_hd__clkbuf_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__2999_ _6035_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2999_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6087__131 _6088__132/A vssd1 vssd1 vccd1 vccd1 _6939_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6897_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3670_ _3337_/X _6902_/Q _3672_/S vssd1 vssd1 vccd1 vccd1 _3671_/A sky130_fd_sc_hd__mux2_1
Xoutput116 _7114_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[17] sky130_fd_sc_hd__buf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5340_ _5351_/B _5340_/B vssd1 vssd1 vccd1 vccd1 _5340_/Y sky130_fd_sc_hd__nor2_1
Xoutput127 _7124_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[27] sky130_fd_sc_hd__buf_2
Xoutput138 _7135_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput149 _7145_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5271_ _5265_/X _5269_/X _5429_/S vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__mux2_1
X_7010_ _7011_/CLK _7010_/D vssd1 vssd1 vccd1 vccd1 _7010_/Q sky130_fd_sc_hd__dfxtp_1
X_4222_ _4222_/A vssd1 vssd1 vccd1 vccd1 _6670_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4153_ _6701_/Q _4152_/X _4156_/S vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4084_ _6750_/Q _5739_/C _4083_/X vssd1 vssd1 vccd1 vccd1 _4085_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2853_ _5750_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2853_/X sky130_fd_sc_hd__clkbuf_16
X_4986_ _4992_/A input9/X _4970_/A _6161_/A vssd1 vssd1 vccd1 vccd1 _4986_/X sky130_fd_sc_hd__a22o_2
X_6725_ _6725_/CLK _6725_/D vssd1 vssd1 vccd1 vccd1 _6725_/Q sky130_fd_sc_hd__dfxtp_1
X_3937_ _3317_/A _3948_/B _5776_/A vssd1 vssd1 vccd1 vccd1 _3937_/Y sky130_fd_sc_hd__a21oi_1
X_5686__420 _5688__422/A vssd1 vssd1 vccd1 vccd1 _6714_/CLK sky130_fd_sc_hd__inv_2
X_3868_ _6741_/Q vssd1 vssd1 vccd1 vccd1 _3868_/X sky130_fd_sc_hd__buf_4
X_6656_ _6656_/CLK _6656_/D vssd1 vssd1 vccd1 vccd1 _6656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3799_ _3693_/X _6832_/Q _3801_/S vssd1 vssd1 vccd1 vccd1 _3800_/A sky130_fd_sc_hd__mux2_1
X_5607_ _5664_/A _5620_/A _5664_/C _5607_/D vssd1 vssd1 vccd1 vccd1 _5659_/B sky130_fd_sc_hd__or4_4
X_6587_ _6587_/CLK _6587_/D vssd1 vssd1 vccd1 vccd1 _6587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7139_ _7139_/A vssd1 vssd1 vccd1 vccd1 _7139_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2535_ clkbuf_0__2535_/X vssd1 vssd1 vccd1 vccd1 _5447__293/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 caravel_wb_data_i[23] vssd1 vssd1 vccd1 vccd1 _5001_/B sky130_fd_sc_hd__buf_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3018_ clkbuf_0__3018_/X vssd1 vssd1 vccd1 vccd1 _6139__174/A sky130_fd_sc_hd__clkbuf_4
Xinput29 caravel_wb_data_i[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5741__447 _5743__449/A vssd1 vssd1 vccd1 vccd1 _6751_/CLK sky130_fd_sc_hd__inv_2
XFILLER_97_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4840_ _4808_/X _4839_/X _4718_/A vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6510_ _6510_/CLK _6510_/D vssd1 vssd1 vccd1 vccd1 _6510_/Q sky130_fd_sc_hd__dfxtp_1
X_4771_ _4936_/S vssd1 vssd1 vccd1 vccd1 _4772_/S sky130_fd_sc_hd__buf_4
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3722_ _3722_/A vssd1 vssd1 vccd1 vccd1 _6862_/D sky130_fd_sc_hd__clkbuf_1
X_6441_ _6441_/CLK _6441_/D vssd1 vssd1 vccd1 vccd1 _6441_/Q sky130_fd_sc_hd__dfxtp_1
X_3653_ _3341_/X _6909_/Q _3653_/S vssd1 vssd1 vccd1 vccd1 _3654_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1_0__3153_ clkbuf_0__3153_/X vssd1 vssd1 vccd1 vccd1 _6338__26/A sky130_fd_sc_hd__clkbuf_4
X_3584_ _3584_/A vssd1 vssd1 vccd1 vccd1 _6936_/D sky130_fd_sc_hd__clkbuf_1
X_5323_ _6575_/Q _5250_/X _5322_/Y _5298_/X vssd1 vssd1 vccd1 vccd1 _6575_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5254_ _5338_/A vssd1 vssd1 vccd1 vccd1 _5254_/X sky130_fd_sc_hd__buf_2
X_4205_ _4205_/A _4259_/B vssd1 vssd1 vccd1 vccd1 _4221_/S sky130_fd_sc_hd__nor2_2
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _4136_/A vssd1 vssd1 vccd1 vccd1 _6708_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4067_ _3273_/B _6730_/Q _3222_/Y _3223_/X vssd1 vssd1 vccd1 vccd1 _4068_/D sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_1_1_0__2868_ clkbuf_0__2868_/X vssd1 vssd1 vccd1 vccd1 _5827__514/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__2836_ _5703_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2836_/X sky130_fd_sc_hd__clkbuf_16
X_4969_ _4969_/A _4969_/B vssd1 vssd1 vccd1 vccd1 _4970_/A sky130_fd_sc_hd__and2_1
X_6708_ _6708_/CLK _6708_/D vssd1 vssd1 vccd1 vccd1 _6708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6639_ _6639_/CLK _6639_/D vssd1 vssd1 vccd1 vccd1 _6639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6132__168 _6132__168/A vssd1 vssd1 vccd1 vccd1 _6976_/CLK sky130_fd_sc_hd__inv_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6990_ _6990_/CLK _6990_/D vssd1 vssd1 vccd1 vccd1 _6990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5941_ _5951_/C vssd1 vssd1 vccd1 vccd1 _5941_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5872_ _5878_/A vssd1 vssd1 vccd1 vccd1 _5872_/X sky130_fd_sc_hd__buf_1
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4823_ _6761_/Q _6753_/Q _6716_/Q _6708_/Q _4701_/A _4806_/A vssd1 vssd1 vccd1 vccd1
+ _4823_/X sky130_fd_sc_hd__mux4_1
XFILLER_21_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4754_ _4762_/C _4754_/B vssd1 vssd1 vccd1 vccd1 _6377_/B sky130_fd_sc_hd__or2_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3705_ _4032_/A vssd1 vssd1 vccd1 vccd1 _3705_/X sky130_fd_sc_hd__clkbuf_2
X_4685_ _4685_/A vssd1 vssd1 vccd1 vccd1 _4685_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_107_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6424_ _7128_/A _6173_/A _6424_/S vssd1 vssd1 vccd1 vccd1 _6425_/B sky130_fd_sc_hd__mux2_1
X_3636_ _3636_/A vssd1 vssd1 vccd1 vccd1 _6916_/D sky130_fd_sc_hd__clkbuf_1
X_6355_ _6355_/A vssd1 vssd1 vccd1 vccd1 _6355_/X sky130_fd_sc_hd__buf_1
X_3567_ _3372_/X _6943_/Q _3571_/S vssd1 vssd1 vccd1 vccd1 _3568_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6286_ _7016_/Q _6284_/X _6285_/X _6192_/X vssd1 vssd1 vccd1 vccd1 _7015_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5306_ _6923_/Q _6915_/Q _7032_/Q _7048_/Q _5281_/X _5282_/X vssd1 vssd1 vccd1 vccd1
+ _5306_/X sky130_fd_sc_hd__mux4_2
X_3498_ _3498_/A vssd1 vssd1 vccd1 vccd1 _6973_/D sky130_fd_sc_hd__clkbuf_1
X_5237_ _5597_/A vssd1 vssd1 vccd1 vccd1 _5237_/X sky130_fd_sc_hd__buf_1
XFILLER_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4119_ _6715_/Q _3892_/X _4121_/S vssd1 vssd1 vccd1 vccd1 _4120_/A sky130_fd_sc_hd__mux2_1
X_5099_ _5099_/A vssd1 vssd1 vccd1 vccd1 _6465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6373__1 _6376__4/A vssd1 vssd1 vccd1 vccd1 _7075_/CLK sky130_fd_sc_hd__inv_2
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6357__41 _6358__42/A vssd1 vssd1 vccd1 vccd1 _7061_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2998_ clkbuf_0__2998_/X vssd1 vssd1 vccd1 vccd1 _6032__88/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4470_ _4026_/X _6552_/Q _4474_/S vssd1 vssd1 vccd1 vccd1 _4471_/A sky130_fd_sc_hd__mux2_1
X_3421_ _3357_/X _7038_/Q _3429_/S vssd1 vssd1 vccd1 vccd1 _3422_/A sky130_fd_sc_hd__mux2_1
X_3352_ _6741_/Q vssd1 vssd1 vccd1 vccd1 _4032_/A sky130_fd_sc_hd__buf_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6140_ _6140_/A vssd1 vssd1 vccd1 vccd1 _6140_/X sky130_fd_sc_hd__buf_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3283_ _7067_/Q _3257_/X _3285_/S vssd1 vssd1 vccd1 vccd1 _3284_/A sky130_fd_sc_hd__mux2_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5022_ _6391_/A vssd1 vssd1 vccd1 vccd1 _6425_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6973_ _6973_/CLK _6973_/D vssd1 vssd1 vccd1 vccd1 _6973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5924_ _6888_/Q _6887_/Q _6886_/Q _5924_/D vssd1 vssd1 vccd1 vccd1 _6015_/B sky130_fd_sc_hd__and4_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _4806_/A vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7022_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_4737_ _4826_/A _4734_/X _4736_/X _4711_/X vssd1 vssd1 vccd1 vccd1 _4737_/X sky130_fd_sc_hd__o211a_1
X_4668_ _3853_/X _6441_/Q _4672_/S vssd1 vssd1 vccd1 vccd1 _4669_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__2535_ _5245_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2535_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2852_ clkbuf_0__2852_/X vssd1 vssd1 vccd1 vccd1 _5747__452/A sky130_fd_sc_hd__clkbuf_4
X_6407_ _7133_/A _6168_/A _6407_/S vssd1 vssd1 vccd1 vccd1 _6408_/B sky130_fd_sc_hd__mux2_1
X_3619_ _3619_/A vssd1 vssd1 vccd1 vccd1 _6923_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4599_ _4599_/A vssd1 vssd1 vccd1 vccd1 _6498_/D sky130_fd_sc_hd__clkbuf_1
X_5544__371 _5544__371/A vssd1 vssd1 vccd1 vccd1 _6661_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6269_ _6269_/A _6269_/B vssd1 vssd1 vccd1 vccd1 _6270_/B sky130_fd_sc_hd__xnor2_1
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3018_ _6134_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3018_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6027__84 _6027__84/A vssd1 vssd1 vccd1 vccd1 _6891_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _6771_/Q vssd1 vssd1 vccd1 vccd1 _4724_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5640_ _5913_/A _6178_/B vssd1 vssd1 vccd1 vccd1 _5640_/Y sky130_fd_sc_hd__xnor2_1
X_5487__325 _5488__326/A vssd1 vssd1 vccd1 vccd1 _6615_/CLK sky130_fd_sc_hd__inv_2
X_4522_ _4476_/X _6533_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4523_/A sky130_fd_sc_hd__mux2_1
X_5680__415 _5682__417/A vssd1 vssd1 vccd1 vccd1 _6709_/CLK sky130_fd_sc_hd__inv_2
X_4453_ _4453_/A vssd1 vssd1 vccd1 vccd1 _6560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3404_ _3329_/X _7045_/Q _3410_/S vssd1 vssd1 vccd1 vccd1 _3405_/A sky130_fd_sc_hd__mux2_1
X_6351__36 _6352__37/A vssd1 vssd1 vccd1 vccd1 _7056_/CLK sky130_fd_sc_hd__inv_2
X_4384_ _6598_/Q _3788_/A _4384_/S vssd1 vssd1 vccd1 vccd1 _4385_/A sky130_fd_sc_hd__mux2_1
X_3335_ _3335_/A vssd1 vssd1 vccd1 vccd1 _7060_/D sky130_fd_sc_hd__clkbuf_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5836__521 _5836__521/A vssd1 vssd1 vccd1 vccd1 _6827_/CLK sky130_fd_sc_hd__inv_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6072_/A vssd1 vssd1 vccd1 vccd1 _6054_/X sky130_fd_sc_hd__buf_1
X_3266_ _7024_/Q vssd1 vssd1 vccd1 vccd1 _3266_/X sky130_fd_sc_hd__buf_2
XFILLER_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5005_ _5005_/A vssd1 vssd1 vccd1 vccd1 _5014_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6956_ _6956_/CLK _6956_/D vssd1 vssd1 vccd1 vccd1 _6956_/Q sky130_fd_sc_hd__dfxtp_1
X_5907_ _4760_/X _6870_/Q _5905_/X _5906_/Y vssd1 vssd1 vccd1 vccd1 _5912_/A sky130_fd_sc_hd__a22o_1
XFILLER_53_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6887_ _6888_/CLK _6887_/D vssd1 vssd1 vccd1 vccd1 _6887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5769_ _5784_/A vssd1 vssd1 vccd1 vccd1 _5769_/X sky130_fd_sc_hd__buf_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2518_ _5163_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2518_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2835_ clkbuf_0__2835_/X vssd1 vssd1 vccd1 vccd1 _5701__433/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5221__271 _5224__274/A vssd1 vssd1 vccd1 vccd1 _6553_/CLK sky130_fd_sc_hd__inv_2
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6810_ _6810_/CLK _6810_/D vssd1 vssd1 vccd1 vccd1 _6810_/Q sky130_fd_sc_hd__dfxtp_1
X_5122__191 _5123__192/A vssd1 vssd1 vccd1 vccd1 _6473_/CLK sky130_fd_sc_hd__inv_2
X_6741_ _7022_/CLK _6741_/D vssd1 vssd1 vccd1 vccd1 _6741_/Q sky130_fd_sc_hd__dfxtp_2
X_3953_ _3953_/A vssd1 vssd1 vccd1 vccd1 _3974_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3884_ _6800_/Q _3883_/X _3887_/S vssd1 vssd1 vccd1 vccd1 _3885_/A sky130_fd_sc_hd__mux2_1
X_6672_ _6672_/CLK _6672_/D vssd1 vssd1 vccd1 vccd1 _6672_/Q sky130_fd_sc_hd__dfxtp_1
X_5623_ _5892_/B _5623_/B vssd1 vssd1 vccd1 vccd1 _5623_/X sky130_fd_sc_hd__and2_1
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5554_ _5554_/A vssd1 vssd1 vccd1 vccd1 _5554_/X sky130_fd_sc_hd__buf_1
XFILLER_117_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4505_ _4505_/A vssd1 vssd1 vccd1 vccd1 _6541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4436_ _3266_/X _6567_/Q _4438_/S vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__mux2_1
X_7155_ _7155_/A vssd1 vssd1 vccd1 vccd1 _7155_/X sky130_fd_sc_hd__clkbuf_1
X_4367_ _4367_/A vssd1 vssd1 vccd1 vccd1 _6606_/D sky130_fd_sc_hd__clkbuf_1
X_5164__225 _5166__227/A vssd1 vssd1 vccd1 vccd1 _6507_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3318_ _3318_/A _3318_/B _3318_/C _3318_/D vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__or4_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _7095_/CLK _7086_/D vssd1 vssd1 vccd1 vccd1 _7086_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _3764_/X _6637_/Q _4306_/S vssd1 vssd1 vccd1 vccd1 _4299_/A sky130_fd_sc_hd__mux2_1
X_3249_ _7078_/Q _3200_/X _3261_/S vssd1 vssd1 vccd1 vccd1 _3250_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2998_ _6028_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2998_/X sky130_fd_sc_hd__clkbuf_16
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _6939_/CLK _6939_/D vssd1 vssd1 vccd1 vccd1 _6939_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2749_ clkbuf_0__2749_/X vssd1 vssd1 vccd1 vccd1 _5572__394/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput117 _7115_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput128 _7099_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[2] sky130_fd_sc_hd__buf_2
Xoutput139 _7136_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_data_o[11] sky130_fd_sc_hd__buf_2
X_5270_ _5286_/A vssd1 vssd1 vccd1 vccd1 _5429_/S sky130_fd_sc_hd__buf_2
XFILLER_114_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4221_ _6670_/Q _4164_/X _4221_/S vssd1 vssd1 vccd1 vccd1 _4222_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5228__277 _5229__278/A vssd1 vssd1 vccd1 vccd1 _6559_/CLK sky130_fd_sc_hd__inv_2
XFILLER_95_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4152_ _7027_/Q vssd1 vssd1 vccd1 vccd1 _4152_/X sky130_fd_sc_hd__buf_4
XFILLER_95_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4083_ _4083_/A vssd1 vssd1 vccd1 vccd1 _4083_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2852_ _5744_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2852_/X sky130_fd_sc_hd__clkbuf_16
X_4985_ _7081_/Q vssd1 vssd1 vccd1 vccd1 _6161_/A sky130_fd_sc_hd__clkbuf_4
X_6724_ _6724_/CLK _6724_/D vssd1 vssd1 vccd1 vccd1 _6724_/Q sky130_fd_sc_hd__dfxtp_1
X_3936_ _3936_/A vssd1 vssd1 vccd1 vccd1 _5776_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3867_ _3867_/A vssd1 vssd1 vccd1 vccd1 _6805_/D sky130_fd_sc_hd__clkbuf_1
X_6655_ _6655_/CLK _6655_/D vssd1 vssd1 vccd1 vccd1 _6655_/Q sky130_fd_sc_hd__dfxtp_1
X_3798_ _3798_/A vssd1 vssd1 vccd1 vccd1 _6833_/D sky130_fd_sc_hd__clkbuf_1
X_5606_ _7087_/Q _7086_/Q _7085_/Q _7084_/Q vssd1 vssd1 vccd1 vccd1 _5607_/D sky130_fd_sc_hd__or4_1
XFILLER_11_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6586_ _6586_/CLK _6586_/D vssd1 vssd1 vccd1 vccd1 _6586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5468_ _5492_/A vssd1 vssd1 vccd1 vccd1 _5468_/X sky130_fd_sc_hd__buf_1
X_5399_ _6927_/Q _6919_/Q _7036_/Q _7052_/Q _4066_/A _5341_/X vssd1 vssd1 vccd1 vccd1
+ _5399_/X sky130_fd_sc_hd__mux4_2
X_4419_ _4419_/A vssd1 vssd1 vccd1 vccd1 _6583_/D sky130_fd_sc_hd__clkbuf_1
X_7138_ _7138_/A vssd1 vssd1 vccd1 vccd1 _7138_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5129__197 _5130__198/A vssd1 vssd1 vccd1 vccd1 _6479_/CLK sky130_fd_sc_hd__inv_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7069_ _7069_/CLK _7069_/D vssd1 vssd1 vccd1 vccd1 _7069_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__2534_ clkbuf_0__2534_/X vssd1 vssd1 vccd1 vccd1 _5242__287/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3017_ clkbuf_0__3017_/X vssd1 vssd1 vccd1 vccd1 _6132__168/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput19 caravel_wb_data_i[24] vssd1 vssd1 vccd1 vccd1 _5003_/B sky130_fd_sc_hd__buf_4
XFILLER_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4770_ _4933_/S _4770_/B vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__or2_1
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3721_ _3699_/X _6862_/Q _3725_/S vssd1 vssd1 vccd1 vccd1 _3722_/A sky130_fd_sc_hd__mux2_1
X_6440_ _6440_/CLK _6440_/D vssd1 vssd1 vccd1 vccd1 _6440_/Q sky130_fd_sc_hd__dfxtp_1
X_3652_ _3652_/A vssd1 vssd1 vccd1 vccd1 _6910_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1_0__3152_ clkbuf_0__3152_/X vssd1 vssd1 vccd1 vccd1 _6335__24/A sky130_fd_sc_hd__clkbuf_4
X_3583_ _6936_/Q _3444_/X _3589_/S vssd1 vssd1 vccd1 vccd1 _3584_/A sky130_fd_sc_hd__mux2_1
X_5322_ _4055_/X _5310_/X _5320_/Y _5321_/X vssd1 vssd1 vccd1 vccd1 _5322_/Y sky130_fd_sc_hd__o211ai_1
X_5253_ _5329_/A vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__buf_2
X_4204_ _4204_/A _4277_/C _6739_/Q vssd1 vssd1 vccd1 vccd1 _4259_/B sky130_fd_sc_hd__or3b_4
XFILLER_68_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4135_ _6708_/Q _3889_/X _4139_/S vssd1 vssd1 vccd1 vccd1 _4136_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4066_ _4066_/A vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__buf_2
XFILLER_52_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__2835_ _5697_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2835_/X sky130_fd_sc_hd__clkbuf_16
X_4968_ _4888_/X input33/X _4969_/B _4967_/X vssd1 vssd1 vccd1 vccd1 _4968_/X sky130_fd_sc_hd__a22o_2
XFILLER_51_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4899_ _3986_/X _6515_/Q _4898_/X _4806_/X vssd1 vssd1 vccd1 vccd1 _4899_/X sky130_fd_sc_hd__o211a_1
X_3919_ _3919_/A vssd1 vssd1 vccd1 vccd1 _6787_/D sky130_fd_sc_hd__clkbuf_1
X_6707_ _6707_/CLK _6707_/D vssd1 vssd1 vccd1 vccd1 _6707_/Q sky130_fd_sc_hd__dfxtp_1
X_6638_ _6638_/CLK _6638_/D vssd1 vssd1 vccd1 vccd1 _6638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6569_ _6569_/CLK _6569_/D vssd1 vssd1 vccd1 vccd1 _6569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5508__342 _5508__342/A vssd1 vssd1 vccd1 vccd1 _6632_/CLK sky130_fd_sc_hd__inv_2
XFILLER_105_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2517_ clkbuf_0__2517_/X vssd1 vssd1 vccd1 vccd1 _5160__222/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2532_ clkbuf_0__2532_/X vssd1 vssd1 vccd1 vccd1 _5529_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5177__235 _5179__237/A vssd1 vssd1 vccd1 vccd1 _6517_/CLK sky130_fd_sc_hd__inv_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5940_ _6871_/Q vssd1 vssd1 vccd1 vccd1 _5951_/C sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0__f__2875_ clkbuf_0__2875_/X vssd1 vssd1 vccd1 vccd1 _5857__57/A sky130_fd_sc_hd__clkbuf_16
X_5830__516 _5831__517/A vssd1 vssd1 vccd1 vccd1 _6822_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4822_ _4826_/A _4822_/B vssd1 vssd1 vccd1 vccd1 _4822_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4753_ _4725_/X _4738_/Y _4856_/B _4883_/B vssd1 vssd1 vccd1 vccd1 _4753_/X sky130_fd_sc_hd__o31a_1
X_3704_ _3704_/A vssd1 vssd1 vccd1 vccd1 _6890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6423_ _6423_/A vssd1 vssd1 vccd1 vccd1 _7092_/D sky130_fd_sc_hd__clkbuf_1
X_4684_ _5050_/B _4686_/B vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__and2_2
X_3635_ _3384_/X _6916_/Q _3639_/S vssd1 vssd1 vccd1 vccd1 _3636_/A sky130_fd_sc_hd__mux2_1
X_3566_ _3566_/A vssd1 vssd1 vccd1 vccd1 _6944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6285_ _7015_/Q _6292_/B vssd1 vssd1 vccd1 vccd1 _6285_/X sky130_fd_sc_hd__or2_1
XFILLER_88_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3497_ _3341_/X _6973_/Q _3497_/S vssd1 vssd1 vccd1 vccd1 _3498_/A sky130_fd_sc_hd__mux2_1
X_5305_ _5355_/B _5305_/B vssd1 vssd1 vccd1 vccd1 _5305_/Y sky130_fd_sc_hd__nor2_1
X_5877__74 _5877__74/A vssd1 vssd1 vccd1 vccd1 _6860_/CLK sky130_fd_sc_hd__inv_2
X_4118_ _4118_/A vssd1 vssd1 vccd1 vccd1 _6716_/D sky130_fd_sc_hd__clkbuf_1
X_5098_ _6465_/Q _7119_/A _5586_/S vssd1 vssd1 vccd1 vccd1 _5099_/A sky130_fd_sc_hd__mux2_1
X_6039__93 _6040__94/A vssd1 vssd1 vccd1 vccd1 _6901_/CLK sky130_fd_sc_hd__inv_2
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4049_ _6303_/B _4049_/B _4049_/C vssd1 vssd1 vccd1 vccd1 _4050_/A sky130_fd_sc_hd__and3_1
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2749_ _5567_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2749_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5699__431 _5701__433/A vssd1 vssd1 vccd1 vccd1 _6725_/CLK sky130_fd_sc_hd__inv_2
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5786__481 _5786__481/A vssd1 vssd1 vccd1 vccd1 _6787_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5708__438 _5709__439/A vssd1 vssd1 vccd1 vccd1 _6732_/CLK sky130_fd_sc_hd__inv_2
X_3420_ _3435_/S vssd1 vssd1 vccd1 vccd1 _3429_/S sky130_fd_sc_hd__clkbuf_2
X_3351_ _3351_/A vssd1 vssd1 vccd1 vccd1 _7056_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3282_ _3282_/A vssd1 vssd1 vccd1 vccd1 _7068_/D sky130_fd_sc_hd__clkbuf_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5021_ _5047_/A vssd1 vssd1 vccd1 vccd1 _6391_/A sky130_fd_sc_hd__clkinv_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5754__458 _5755__459/A vssd1 vssd1 vccd1 vccd1 _6762_/CLK sky130_fd_sc_hd__inv_2
XFILLER_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6972_ _6972_/CLK _6972_/D vssd1 vssd1 vccd1 vccd1 _6972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5923_ _6017_/A vssd1 vssd1 vccd1 vccd1 _5926_/B sky130_fd_sc_hd__clkbuf_2
X_5854_ _5866_/A vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__buf_1
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4805_ _4906_/A vssd1 vssd1 vccd1 vccd1 _4806_/A sky130_fd_sc_hd__buf_4
XFILLER_21_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4736_ _4875_/S _4736_/B vssd1 vssd1 vccd1 vccd1 _4736_/X sky130_fd_sc_hd__or2_1
XFILLER_119_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4667_ _4667_/A vssd1 vssd1 vccd1 vccd1 _6442_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2534_ _5239_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2534_/X sky130_fd_sc_hd__clkbuf_16
X_6406_ _6406_/A vssd1 vssd1 vccd1 vccd1 _7087_/D sky130_fd_sc_hd__clkbuf_1
X_3618_ _6923_/Q _3617_/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3619_/A sky130_fd_sc_hd__mux2_1
X_4598_ _6498_/Q _4020_/A _4600_/S vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3549_ _6951_/Q _3447_/X _3553_/S vssd1 vssd1 vccd1 vccd1 _3550_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6268_ _6268_/A vssd1 vssd1 vccd1 vccd1 _7010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5219_ _5231_/A vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__buf_1
X_6199_ _6271_/A _6271_/B vssd1 vssd1 vccd1 vccd1 _6282_/A sky130_fd_sc_hd__and2b_1
X_5247__291 _5448__294/A vssd1 vssd1 vccd1 vccd1 _6573_/CLK sky130_fd_sc_hd__inv_2
XFILLER_28_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__3017_ _6128_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3017_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6081__127 _6082__128/A vssd1 vssd1 vccd1 vccd1 _6935_/CLK sky130_fd_sc_hd__inv_2
XFILLER_100_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5871__69 _5871__69/A vssd1 vssd1 vccd1 vccd1 _6855_/CLK sky130_fd_sc_hd__inv_2
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4521_ _4536_/S vssd1 vssd1 vccd1 vccd1 _4530_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_117_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4452_ _4026_/X _6560_/Q _4456_/S vssd1 vssd1 vccd1 vccd1 _4453_/A sky130_fd_sc_hd__mux2_1
X_5760__462 _5760__462/A vssd1 vssd1 vccd1 vccd1 _6766_/CLK sky130_fd_sc_hd__inv_2
X_3403_ _3403_/A vssd1 vssd1 vccd1 vccd1 _7046_/D sky130_fd_sc_hd__clkbuf_1
X_4383_ _4383_/A vssd1 vssd1 vccd1 vccd1 _6599_/D sky130_fd_sc_hd__clkbuf_1
X_3334_ _3333_/X _7060_/Q _3342_/S vssd1 vssd1 vccd1 vccd1 _3335_/A sky130_fd_sc_hd__mux2_1
X_6122_ _6128_/A vssd1 vssd1 vccd1 vccd1 _6122_/X sky130_fd_sc_hd__buf_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6053_ _6084_/A vssd1 vssd1 vccd1 vccd1 _6053_/X sky130_fd_sc_hd__buf_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3265_/A vssd1 vssd1 vccd1 vccd1 _7073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5004_ _5004_/A vssd1 vssd1 vccd1 vccd1 _5004_/X sky130_fd_sc_hd__clkbuf_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6955_ _6955_/CLK _6955_/D vssd1 vssd1 vccd1 vccd1 _6955_/Q sky130_fd_sc_hd__dfxtp_1
X_5906_ _6872_/Q _5906_/B _5906_/C vssd1 vssd1 vccd1 vccd1 _5906_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6886_ _6888_/CLK _6886_/D vssd1 vssd1 vccd1 vccd1 _6886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6145__179 _6145__179/A vssd1 vssd1 vccd1 vccd1 _6987_/CLK sky130_fd_sc_hd__inv_2
X_4719_ _4719_/A vssd1 vssd1 vccd1 vccd1 _4719_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__2517_ _5157_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2517_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2834_ clkbuf_0__2834_/X vssd1 vssd1 vccd1 vccd1 _5696__429/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5493__330 _5494__331/A vssd1 vssd1 vccd1 vccd1 _6620_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6740_ _6740_/CLK _6740_/D vssd1 vssd1 vccd1 vccd1 _6740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3952_ _6770_/Q vssd1 vssd1 vccd1 vccd1 _3953_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3883_ _6745_/Q vssd1 vssd1 vccd1 vccd1 _3883_/X sky130_fd_sc_hd__clkbuf_4
X_6671_ _6671_/CLK _6671_/D vssd1 vssd1 vccd1 vccd1 _6671_/Q sky130_fd_sc_hd__dfxtp_1
X_5622_ _5890_/A _5890_/B _4974_/X vssd1 vssd1 vccd1 vccd1 _5623_/B sky130_fd_sc_hd__a21bo_1
X_4504_ _4476_/X _6541_/Q _4512_/S vssd1 vssd1 vccd1 vccd1 _4505_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4435_ _4435_/A vssd1 vssd1 vccd1 vccd1 _6568_/D sky130_fd_sc_hd__clkbuf_1
X_7154_ _7154_/A vssd1 vssd1 vccd1 vccd1 _7154_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4366_ _6606_/Q _3788_/A _4366_/S vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5799__491 _5799__491/A vssd1 vssd1 vccd1 vccd1 _6797_/CLK sky130_fd_sc_hd__inv_2
X_3317_ _3317_/A _3961_/B vssd1 vssd1 vccd1 vccd1 _3318_/D sky130_fd_sc_hd__xnor2_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5502__337 _5502__337/A vssd1 vssd1 vccd1 vccd1 _6627_/CLK sky130_fd_sc_hd__inv_2
X_7085_ _7089_/CLK _7085_/D vssd1 vssd1 vccd1 vccd1 _7085_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4312_/S vssd1 vssd1 vccd1 vccd1 _4306_/S sky130_fd_sc_hd__buf_2
XFILLER_100_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3248_ _3270_/S vssd1 vssd1 vccd1 vccd1 _3261_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6938_ _6938_/CLK _6938_/D vssd1 vssd1 vccd1 vccd1 _6938_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6869_ _6883_/CLK _6869_/D vssd1 vssd1 vccd1 vccd1 _6869_/Q sky130_fd_sc_hd__dfxtp_1
X_5767__468 _5768__469/A vssd1 vssd1 vccd1 vccd1 _6772_/CLK sky130_fd_sc_hd__inv_2
XFILLER_108_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2748_ clkbuf_0__2748_/X vssd1 vssd1 vccd1 vccd1 _5566__389/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5557__382 _5557__382/A vssd1 vssd1 vccd1 vccd1 _6672_/CLK sky130_fd_sc_hd__inv_2
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput107 _6467_/Q vssd1 vssd1 vccd1 vccd1 caravel_uart_tx sky130_fd_sc_hd__buf_2
Xoutput118 _7116_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[19] sky130_fd_sc_hd__buf_2
Xoutput129 _7100_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[3] sky130_fd_sc_hd__buf_2
X_6094__137 _6094__137/A vssd1 vssd1 vccd1 vccd1 _6945_/CLK sky130_fd_sc_hd__inv_2
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4220_ _4220_/A vssd1 vssd1 vccd1 vccd1 _6671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4151_ _4151_/A vssd1 vssd1 vccd1 vccd1 _6702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4082_ _5281_/A vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__buf_4
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4984_ _5005_/A vssd1 vssd1 vccd1 vccd1 _4992_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6723_ _6723_/CLK _6723_/D vssd1 vssd1 vccd1 vccd1 _6723_/Q sky130_fd_sc_hd__dfxtp_1
X_3935_ _6777_/Q _6778_/Q _3485_/B _5723_/B vssd1 vssd1 vccd1 vccd1 _6777_/D sky130_fd_sc_hd__o211a_1
X_6654_ _6654_/CLK _6654_/D vssd1 vssd1 vccd1 vccd1 _6654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5170__230 _5172__232/A vssd1 vssd1 vccd1 vccd1 _6512_/CLK sky130_fd_sc_hd__inv_2
X_3866_ _6805_/Q _3865_/X _3869_/S vssd1 vssd1 vccd1 vccd1 _3867_/A sky130_fd_sc_hd__mux2_1
X_5605_ _7089_/Q _7088_/Q vssd1 vssd1 vccd1 vccd1 _5664_/C sky130_fd_sc_hd__or2_2
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3797_ _3690_/X _6833_/Q _3801_/S vssd1 vssd1 vccd1 vccd1 _3798_/A sky130_fd_sc_hd__mux2_1
X_6585_ _6585_/CLK _6585_/D vssd1 vssd1 vccd1 vccd1 _6585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5536_ _5554_/A vssd1 vssd1 vccd1 vccd1 _5536_/X sky130_fd_sc_hd__buf_1
X_5467_ _5529_/A vssd1 vssd1 vccd1 vccd1 _5467_/X sky130_fd_sc_hd__buf_1
X_4418_ _3266_/X _6583_/Q _4420_/S vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__mux2_1
X_5398_ _5437_/A _5398_/B vssd1 vssd1 vccd1 vccd1 _5398_/Y sky130_fd_sc_hd__nor2_1
X_7137_ _7137_/A vssd1 vssd1 vccd1 vccd1 _7137_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4349_ _4349_/A vssd1 vssd1 vccd1 vccd1 _6614_/D sky130_fd_sc_hd__clkbuf_1
X_5693__426 _5694__427/A vssd1 vssd1 vccd1 vccd1 _6720_/CLK sky130_fd_sc_hd__inv_2
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7068_ _7068_/CLK _7068_/D vssd1 vssd1 vccd1 vccd1 _7068_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__2533_ clkbuf_0__2533_/X vssd1 vssd1 vccd1 vccd1 _5461_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6019_ _6021_/B _6019_/B _6019_/C vssd1 vssd1 vccd1 vccd1 _6020_/A sky130_fd_sc_hd__and3b_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5849__532 _5849__532/A vssd1 vssd1 vccd1 vccd1 _6838_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__3016_ clkbuf_0__3016_/X vssd1 vssd1 vccd1 vccd1 _6124__161/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6154__10 _6154__10/A vssd1 vssd1 vccd1 vccd1 _6993_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5780__476 _5780__476/A vssd1 vssd1 vccd1 vccd1 _6782_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3720_ _3720_/A vssd1 vssd1 vccd1 vccd1 _6863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5234__282 _5235__283/A vssd1 vssd1 vccd1 vccd1 _6564_/CLK sky130_fd_sc_hd__inv_2
X_3651_ _3337_/X _6910_/Q _3653_/S vssd1 vssd1 vccd1 vccd1 _3652_/A sky130_fd_sc_hd__mux2_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3582_ _3582_/A vssd1 vssd1 vccd1 vccd1 _6937_/D sky130_fd_sc_hd__clkbuf_1
X_6102__144 _6102__144/A vssd1 vssd1 vccd1 vccd1 _6952_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0__3151_ clkbuf_0__3151_/X vssd1 vssd1 vccd1 vccd1 _6329__19/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5321_ _5321_/A vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5252_ _5258_/A vssd1 vssd1 vccd1 vccd1 _5329_/A sky130_fd_sc_hd__buf_2
X_4203_ _4203_/A vssd1 vssd1 vccd1 vccd1 _6678_/D sky130_fd_sc_hd__clkbuf_1
X_4134_ _4134_/A vssd1 vssd1 vccd1 vccd1 _6709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4065_ _5281_/A vssd1 vssd1 vccd1 vccd1 _4066_/A sky130_fd_sc_hd__clkbuf_4
X_5241__286 _5244__289/A vssd1 vssd1 vccd1 vccd1 _6568_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_0__2834_ _5691_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2834_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _6168_/A _4987_/C _4856_/Y vssd1 vssd1 vccd1 vccd1 _4967_/X sky130_fd_sc_hd__a21o_1
X_6369__51 _6372__54/A vssd1 vssd1 vccd1 vccd1 _7071_/CLK sky130_fd_sc_hd__inv_2
X_4898_ _4898_/A _6499_/Q vssd1 vssd1 vccd1 vccd1 _4898_/X sky130_fd_sc_hd__or2_1
X_3918_ _6787_/Q _3871_/X _3926_/S vssd1 vssd1 vccd1 vccd1 _3919_/A sky130_fd_sc_hd__mux2_1
X_6706_ _6706_/CLK _6706_/D vssd1 vssd1 vccd1 vccd1 _6706_/Q sky130_fd_sc_hd__dfxtp_1
X_3849_ _3849_/A vssd1 vssd1 vccd1 vccd1 _6811_/D sky130_fd_sc_hd__clkbuf_1
X_6637_ _6637_/CLK _6637_/D vssd1 vssd1 vccd1 vccd1 _6637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6568_ _6568_/CLK _6568_/D vssd1 vssd1 vccd1 vccd1 _6568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6499_ _6499_/CLK _6499_/D vssd1 vssd1 vccd1 vccd1 _6499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5701__433 _5701__433/A vssd1 vssd1 vccd1 vccd1 _6727_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2516_ clkbuf_0__2516_/X vssd1 vssd1 vccd1 vccd1 _5156__219/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4821_ _6472_/Q _6624_/Q _7057_/Q _6782_/Q _3958_/A _4956_/S vssd1 vssd1 vccd1 vccd1
+ _4822_/B sky130_fd_sc_hd__mux4_1
X_4752_ _4762_/C _4752_/B _4766_/C vssd1 vssd1 vccd1 vccd1 _4883_/B sky130_fd_sc_hd__or3_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3703_ _3702_/X _6890_/Q _3706_/S vssd1 vssd1 vccd1 vccd1 _3704_/A sky130_fd_sc_hd__mux2_1
X_4683_ _5005_/A _4683_/B _4683_/C _4683_/D vssd1 vssd1 vccd1 vccd1 _4686_/B sky130_fd_sc_hd__and4_4
X_6422_ _6425_/A _6422_/B vssd1 vssd1 vccd1 vccd1 _6423_/A sky130_fd_sc_hd__and2_1
X_3634_ _3634_/A vssd1 vssd1 vccd1 vccd1 _6917_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3565_ _3368_/X _6944_/Q _3571_/S vssd1 vssd1 vccd1 vccd1 _3566_/A sky130_fd_sc_hd__mux2_1
X_6284_ _6284_/A vssd1 vssd1 vccd1 vccd1 _6284_/X sky130_fd_sc_hd__clkbuf_2
X_3496_ _3496_/A vssd1 vssd1 vccd1 vccd1 _6974_/D sky130_fd_sc_hd__clkbuf_1
X_5304_ _6947_/Q _6679_/Q _6591_/Q _6813_/Q _4083_/X _4070_/A vssd1 vssd1 vccd1 vccd1
+ _5305_/B sky130_fd_sc_hd__mux4_1
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4117_ _6716_/Q _3889_/X _4121_/S vssd1 vssd1 vccd1 vccd1 _4118_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5097_ _5097_/A vssd1 vssd1 vccd1 vccd1 _6464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4048_ _4048_/A _4052_/B vssd1 vssd1 vccd1 vccd1 _4049_/C sky130_fd_sc_hd__nand2_1
XFILLER_71_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5999_ _5999_/A vssd1 vssd1 vccd1 vccd1 _6881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__2748_ _5561_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2748_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5183__240 _5187__244/A vssd1 vssd1 vccd1 vccd1 _6522_/CLK sky130_fd_sc_hd__inv_2
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6363__46 _6363__46/A vssd1 vssd1 vccd1 vccd1 _7066_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3350_ _3349_/X _7056_/Q _3354_/S vssd1 vssd1 vccd1 vccd1 _3351_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _6444_/Q vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__inv_2
X_3281_ _7068_/Q _3254_/X _3285_/S vssd1 vssd1 vccd1 vccd1 _3282_/A sky130_fd_sc_hd__mux2_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5793__486 _5796__489/A vssd1 vssd1 vccd1 vccd1 _6792_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5457__301 _5458__302/A vssd1 vssd1 vccd1 vccd1 _6591_/CLK sky130_fd_sc_hd__inv_2
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6971_ _6971_/CLK _6971_/D vssd1 vssd1 vccd1 vccd1 _6971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5922_ _5922_/A _5922_/B _5922_/C _5922_/D vssd1 vssd1 vccd1 vccd1 _6017_/A sky130_fd_sc_hd__or4_4
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5853_ _6115_/A vssd1 vssd1 vccd1 vccd1 _5853_/X sky130_fd_sc_hd__buf_1
X_4804_ _4804_/A _4804_/B vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__or2_1
X_5784_ _5784_/A vssd1 vssd1 vccd1 vccd1 _5784_/X sky130_fd_sc_hd__buf_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4735_ _6542_/Q _6722_/Q _6860_/Q _6526_/Q _4845_/A _4701_/A vssd1 vssd1 vccd1 vccd1
+ _4736_/B sky130_fd_sc_hd__mux4_1
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4666_ _3850_/X _6442_/Q _4672_/S vssd1 vssd1 vccd1 vccd1 _4667_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_0__2533_ _5238_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2533_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4597_ _4597_/A vssd1 vssd1 vccd1 vccd1 _6499_/D sky130_fd_sc_hd__clkbuf_1
X_6405_ _6408_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6406_/A sky130_fd_sc_hd__and2_1
X_3617_ _7024_/Q vssd1 vssd1 vccd1 vccd1 _3617_/X sky130_fd_sc_hd__clkbuf_4
X_6336_ _6336_/A vssd1 vssd1 vccd1 vccd1 _6336_/X sky130_fd_sc_hd__buf_1
X_3548_ _3548_/A vssd1 vssd1 vccd1 vccd1 _6952_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6267_ _6267_/A _6267_/B _6269_/B vssd1 vssd1 vccd1 vccd1 _6268_/A sky130_fd_sc_hd__and3_1
X_3479_ _3479_/A vssd1 vssd1 vccd1 vccd1 _6980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6198_ _6995_/Q _6179_/X _6290_/A vssd1 vssd1 vccd1 vccd1 _6270_/A sky130_fd_sc_hd__o21ai_2
Xclkbuf_0__3016_ _6122_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3016_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_56_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5551__377 _5553__379/A vssd1 vssd1 vccd1 vccd1 _6667_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5856__56 _5857__57/A vssd1 vssd1 vccd1 vccd1 _6842_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5714__443 _5715__444/A vssd1 vssd1 vccd1 vccd1 _6737_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6033__89 _6033__89/A vssd1 vssd1 vccd1 vccd1 _6896_/CLK sky130_fd_sc_hd__inv_2
X_5452__297 _5453__298/A vssd1 vssd1 vccd1 vccd1 _6587_/CLK sky130_fd_sc_hd__inv_2
X_4520_ _4608_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4536_/S sky130_fd_sc_hd__or2_2
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4451_ _4451_/A vssd1 vssd1 vccd1 vccd1 _6561_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6058__108 _6059__109/A vssd1 vssd1 vccd1 vccd1 _6916_/CLK sky130_fd_sc_hd__inv_2
X_3402_ _3294_/X _7046_/Q _3410_/S vssd1 vssd1 vccd1 vccd1 _3403_/A sky130_fd_sc_hd__mux2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ _6599_/Q _3785_/A _4384_/S vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__mux2_1
X_3333_ _4017_/A vssd1 vssd1 vccd1 vccd1 _3333_/X sky130_fd_sc_hd__buf_2
XFILLER_98_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5801__493 _5802__494/A vssd1 vssd1 vccd1 vccd1 _6799_/CLK sky130_fd_sc_hd__inv_2
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _7073_/Q _3263_/X _3270_/S vssd1 vssd1 vccd1 vccd1 _3265_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5003_ _5003_/A _5003_/B vssd1 vssd1 vccd1 vccd1 _5004_/A sky130_fd_sc_hd__and2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6954_ _6954_/CLK _6954_/D vssd1 vssd1 vccd1 vccd1 _6954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5905_ _5906_/B _5906_/C _5951_/B vssd1 vssd1 vccd1 vccd1 _5905_/X sky130_fd_sc_hd__a21bo_1
X_6885_ _7008_/CLK _6885_/D vssd1 vssd1 vccd1 vccd1 _6885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5134__201 _5137__204/A vssd1 vssd1 vccd1 vccd1 _6483_/CLK sky130_fd_sc_hd__inv_2
XFILLER_22_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4718_ _4718_/A vssd1 vssd1 vccd1 vccd1 _4826_/A sky130_fd_sc_hd__clkbuf_2
X_5843__527 _5843__527/A vssd1 vssd1 vccd1 vccd1 _6833_/CLK sky130_fd_sc_hd__inv_2
XFILLER_30_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2516_ _5151_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2516_/X sky130_fd_sc_hd__clkbuf_16
X_4649_ _4649_/A vssd1 vssd1 vccd1 vccd1 _6476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2833_ clkbuf_0__2833_/X vssd1 vssd1 vccd1 vccd1 _5688__422/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6319_ _6319_/A vssd1 vssd1 vccd1 vccd1 _7030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3951_ _6771_/Q vssd1 vssd1 vccd1 vccd1 _3951_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_63_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3882_ _3882_/A vssd1 vssd1 vccd1 vccd1 _6801_/D sky130_fd_sc_hd__clkbuf_1
X_6670_ _6670_/CLK _6670_/D vssd1 vssd1 vccd1 vccd1 _6670_/Q sky130_fd_sc_hd__dfxtp_1
X_5621_ _5913_/A _5913_/B _5664_/C vssd1 vssd1 vccd1 vccd1 _5890_/B sky130_fd_sc_hd__nor3_4
XFILLER_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4503_ _4518_/S vssd1 vssd1 vccd1 vccd1 _4512_/S sky130_fd_sc_hd__buf_2
X_4434_ _3263_/X _6568_/Q _4438_/S vssd1 vssd1 vccd1 vccd1 _4435_/A sky130_fd_sc_hd__mux2_1
X_7153_ _7153_/A vssd1 vssd1 vccd1 vccd1 _7153_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4365_ _4365_/A vssd1 vssd1 vccd1 vccd1 _6607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3316_ _6776_/Q _6771_/Q vssd1 vssd1 vccd1 vccd1 _3961_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7084_ _7095_/CLK _7084_/D vssd1 vssd1 vccd1 vccd1 _7084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6035_ _6047_/A vssd1 vssd1 vccd1 vccd1 _6035_/X sky130_fd_sc_hd__buf_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _4296_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4312_/S sky130_fd_sc_hd__or2_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _4422_/A _4205_/A vssd1 vssd1 vccd1 vccd1 _3270_/S sky130_fd_sc_hd__nor2_2
XFILLER_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6937_ _6937_/CLK _6937_/D vssd1 vssd1 vccd1 vccd1 _6937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6868_ _6888_/CLK _6868_/D vssd1 vssd1 vccd1 vccd1 _6868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6799_ _6799_/CLK _6799_/D vssd1 vssd1 vccd1 vccd1 _6799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5808__499 _5808__499/A vssd1 vssd1 vccd1 vccd1 _6805_/CLK sky130_fd_sc_hd__inv_2
XFILLER_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2747_ clkbuf_0__2747_/X vssd1 vssd1 vccd1 vccd1 _5573_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput119 _7098_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[1] sky130_fd_sc_hd__buf_2
Xoutput108 _7097_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[0] sky130_fd_sc_hd__buf_2
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5564__387 _5564__387/A vssd1 vssd1 vccd1 vccd1 _6677_/CLK sky130_fd_sc_hd__inv_2
XFILLER_68_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4150_ _6702_/Q _4149_/X _4156_/S vssd1 vssd1 vccd1 vccd1 _4151_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4081_ _4081_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _6731_/D sky130_fd_sc_hd__nor2_1
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4983_ _4973_/X input8/X _4970_/A _6155_/A vssd1 vssd1 vccd1 vccd1 _4983_/X sky130_fd_sc_hd__a22o_2
XFILLER_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6722_ _6722_/CLK _6722_/D vssd1 vssd1 vccd1 vccd1 _6722_/Q sky130_fd_sc_hd__dfxtp_1
X_3934_ _3947_/A vssd1 vssd1 vccd1 vccd1 _5723_/B sky130_fd_sc_hd__buf_4
XFILLER_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3865_ _6742_/Q vssd1 vssd1 vccd1 vccd1 _3865_/X sky130_fd_sc_hd__clkbuf_4
X_6653_ _6653_/CLK _6653_/D vssd1 vssd1 vccd1 vccd1 _6653_/Q sky130_fd_sc_hd__dfxtp_1
X_5604_ _7091_/Q _7090_/Q vssd1 vssd1 vccd1 vccd1 _5620_/A sky130_fd_sc_hd__or2_1
X_3796_ _3796_/A vssd1 vssd1 vccd1 vccd1 _6834_/D sky130_fd_sc_hd__clkbuf_1
X_6584_ _6584_/CLK _6584_/D vssd1 vssd1 vccd1 vccd1 _6584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4417_ _4417_/A vssd1 vssd1 vccd1 vccd1 _6584_/D sky130_fd_sc_hd__clkbuf_1
X_5397_ _6951_/Q _6683_/Q _6595_/Q _6817_/Q _5337_/X _5338_/X vssd1 vssd1 vccd1 vccd1
+ _5398_/B sky130_fd_sc_hd__mux4_2
XFILLER_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7136_ _7136_/A vssd1 vssd1 vccd1 vccd1 _7136_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4348_ _3788_/X _6614_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7067_ _7067_/CLK _7067_/D vssd1 vssd1 vccd1 vccd1 _7067_/Q sky130_fd_sc_hd__dfxtp_1
X_4279_ _4294_/S vssd1 vssd1 vccd1 vccd1 _4288_/S sky130_fd_sc_hd__buf_2
XFILLER_100_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6018_ _5924_/D _5929_/B _6017_/Y _6886_/Q vssd1 vssd1 vccd1 vccd1 _6019_/C sky130_fd_sc_hd__a31o_1
XFILLER_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5773__473 _5773__473/A vssd1 vssd1 vccd1 vccd1 _6777_/CLK sky130_fd_sc_hd__inv_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0__3015_ clkbuf_0__3015_/X vssd1 vssd1 vccd1 vccd1 _6121__159/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5147__211 _5147__211/A vssd1 vssd1 vccd1 vccd1 _6493_/CLK sky130_fd_sc_hd__inv_2
XFILLER_2_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3650_ _3650_/A vssd1 vssd1 vccd1 vccd1 _6911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3581_ _6937_/Q _3437_/X _3589_/S vssd1 vssd1 vccd1 vccd1 _3582_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5320_ _5366_/A _5320_/B vssd1 vssd1 vccd1 vccd1 _5320_/Y sky130_fd_sc_hd__nand2_1
X_5251_ _5281_/A vssd1 vssd1 vccd1 vccd1 _5251_/X sky130_fd_sc_hd__buf_4
XFILLER_114_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4202_ _6678_/Q _4164_/X _4202_/S vssd1 vssd1 vccd1 vccd1 _4203_/A sky130_fd_sc_hd__mux2_1
X_5182_ _5188_/A vssd1 vssd1 vccd1 vccd1 _5182_/X sky130_fd_sc_hd__buf_1
XFILLER_114_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4133_ _6709_/Q _3886_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4134_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4064_ _6730_/Q vssd1 vssd1 vccd1 vccd1 _5281_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1_0__2865_ clkbuf_0__2865_/X vssd1 vssd1 vccd1 vccd1 _5814__504/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__2833_ _5685_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2833_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6705_ _7093_/CLK _6705_/D vssd1 vssd1 vccd1 vccd1 _6705_/Q sky130_fd_sc_hd__dfxtp_2
X_4966_ _7088_/Q vssd1 vssd1 vccd1 vccd1 _6168_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4897_ _4893_/X _4895_/X _4896_/X _4933_/S _4722_/X vssd1 vssd1 vccd1 vccd1 _4904_/B
+ sky130_fd_sc_hd__o221a_1
X_3917_ _3932_/S vssd1 vssd1 vccd1 vccd1 _3926_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3848_ _6811_/Q _3845_/X _3860_/S vssd1 vssd1 vccd1 vccd1 _3849_/A sky130_fd_sc_hd__mux2_1
X_6636_ _6636_/CLK _6636_/D vssd1 vssd1 vccd1 vccd1 _6636_/Q sky130_fd_sc_hd__dfxtp_1
X_3779_ _3779_/A vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__clkbuf_2
X_6567_ _6567_/CLK _6567_/D vssd1 vssd1 vccd1 vccd1 _6567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7079_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_6498_ _6498_/CLK _6498_/D vssd1 vssd1 vccd1 vccd1 _6498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5449_ _5449_/A vssd1 vssd1 vccd1 vccd1 _5449_/X sky130_fd_sc_hd__buf_1
XFILLER_99_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7119_ _7119_/A vssd1 vssd1 vccd1 vccd1 _7119_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2515_ clkbuf_0__2515_/X vssd1 vssd1 vccd1 vccd1 _5147__211/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5515__348 _5516__349/A vssd1 vssd1 vccd1 vccd1 _6638_/CLK sky130_fd_sc_hd__inv_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5596__409 _5596__409/A vssd1 vssd1 vccd1 vccd1 _6702_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4820_ _4802_/X _4804_/X _4812_/X _4819_/X _4904_/A vssd1 vssd1 vccd1 vccd1 _4820_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4795_/A _4794_/C vssd1 vssd1 vccd1 vccd1 _4766_/C sky130_fd_sc_hd__nand2_1
XFILLER_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3702_ _4029_/A vssd1 vssd1 vccd1 vccd1 _3702_/X sky130_fd_sc_hd__buf_2
X_4682_ _4682_/A _4682_/B vssd1 vssd1 vccd1 vccd1 _4683_/D sky130_fd_sc_hd__nor2_2
X_6421_ _7129_/A _4885_/X _6424_/S vssd1 vssd1 vccd1 vccd1 _6422_/B sky130_fd_sc_hd__mux2_1
X_3633_ _3380_/X _6917_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _3634_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3564_ _3564_/A vssd1 vssd1 vccd1 vccd1 _6945_/D sky130_fd_sc_hd__clkbuf_1
X_6283_ _6300_/B vssd1 vssd1 vccd1 vccd1 _6284_/A sky130_fd_sc_hd__inv_2
X_3495_ _3337_/X _6974_/Q _3497_/S vssd1 vssd1 vccd1 vccd1 _3496_/A sky130_fd_sc_hd__mux2_1
X_5303_ _5439_/B vssd1 vssd1 vccd1 vccd1 _5355_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4116_ _4116_/A vssd1 vssd1 vccd1 vccd1 _6717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ _6464_/Q _7118_/A _5586_/S vssd1 vssd1 vccd1 vccd1 _5097_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4047_ _4051_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _4052_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _6002_/A _5998_/B vssd1 vssd1 vccd1 vccd1 _5999_/A sky130_fd_sc_hd__and2_1
X_4949_ _6766_/Q _6758_/Q _6721_/Q _6713_/Q _4923_/X _4892_/X vssd1 vssd1 vccd1 vccd1
+ _4949_/X sky130_fd_sc_hd__mux4_2
XFILLER_20_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2747_ _5560_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2747_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6619_ _6619_/CLK _6619_/D vssd1 vssd1 vccd1 vccd1 _6619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5883__79 _5883__79/A vssd1 vssd1 vccd1 vccd1 _6865_/CLK sky130_fd_sc_hd__inv_2
X_6051__103 _6052__104/A vssd1 vssd1 vccd1 vccd1 _6911_/CLK sky130_fd_sc_hd__inv_2
XFILLER_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6045__98 _6046__99/A vssd1 vssd1 vccd1 vccd1 _6906_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5038__185 _5040__187/A vssd1 vssd1 vccd1 vccd1 _6441_/CLK sky130_fd_sc_hd__inv_2
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3280_ _3280_/A vssd1 vssd1 vccd1 vccd1 _7069_/D sky130_fd_sc_hd__clkbuf_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6970_ _6970_/CLK _6970_/D vssd1 vssd1 vccd1 vccd1 _6970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5921_ _5921_/A _5921_/B _5921_/C _5921_/D vssd1 vssd1 vccd1 vccd1 _5922_/D sky130_fd_sc_hd__or4_1
XFILLER_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5852_ _5852_/A vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__buf_1
X_4803_ _6900_/Q _6560_/Q _6908_/Q _6488_/Q _4719_/A _4807_/S vssd1 vssd1 vccd1 vccd1
+ _4804_/B sky130_fd_sc_hd__mux4_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4734_ _6889_/Q _6518_/Q _6494_/Q _6510_/Q _4891_/B _4709_/X vssd1 vssd1 vccd1 vccd1
+ _4734_/X sky130_fd_sc_hd__mux4_1
X_4665_ _4665_/A vssd1 vssd1 vccd1 vccd1 _6443_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__2532_ _5237_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2532_/X sky130_fd_sc_hd__clkbuf_16
X_4596_ _6499_/Q _4017_/A _4600_/S vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__mux2_1
X_6404_ _7134_/A _5663_/A _6407_/S vssd1 vssd1 vccd1 vccd1 _6405_/B sky130_fd_sc_hd__mux2_1
X_3616_ _3616_/A vssd1 vssd1 vccd1 vccd1 _6924_/D sky130_fd_sc_hd__clkbuf_1
X_3547_ _6952_/Q _3444_/X _3553_/S vssd1 vssd1 vccd1 vccd1 _3548_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6266_ _6266_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6269_/B sky130_fd_sc_hd__nand2_1
X_3478_ _3384_/X _6980_/Q _3482_/S vssd1 vssd1 vccd1 vccd1 _3479_/A sky130_fd_sc_hd__mux2_1
X_6197_ _6216_/C _6187_/B _6196_/Y _6192_/X vssd1 vssd1 vccd1 vccd1 _6996_/D sky130_fd_sc_hd__o211a_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3015_ _6116_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3015_/X sky130_fd_sc_hd__clkbuf_16
X_5079_ _5079_/A vssd1 vssd1 vccd1 vccd1 _6456_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4450_ _4023_/X _6561_/Q _4450_/S vssd1 vssd1 vccd1 vccd1 _4451_/A sky130_fd_sc_hd__mux2_1
X_3401_ _3416_/S vssd1 vssd1 vccd1 vccd1 _3410_/S sky130_fd_sc_hd__clkbuf_2
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _6600_/D sky130_fd_sc_hd__clkbuf_1
X_3332_ _6746_/Q vssd1 vssd1 vccd1 vccd1 _4017_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3263_ _7025_/Q vssd1 vssd1 vccd1 vccd1 _3263_/X sky130_fd_sc_hd__clkbuf_4
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5002_ _5002_/A vssd1 vssd1 vccd1 vccd1 _5002_/X sky130_fd_sc_hd__clkbuf_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6953_ _6953_/CLK _6953_/D vssd1 vssd1 vccd1 vccd1 _6953_/Q sky130_fd_sc_hd__dfxtp_1
X_5904_ _6872_/Q vssd1 vssd1 vccd1 vccd1 _5951_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6884_ _7008_/CLK _6884_/D vssd1 vssd1 vccd1 vccd1 _6884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5697_ _5697_/A vssd1 vssd1 vccd1 vccd1 _5697_/X sky130_fd_sc_hd__buf_1
X_4717_ _4732_/A vssd1 vssd1 vccd1 vccd1 _4718_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_0__2515_ _5145_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2515_/X sky130_fd_sc_hd__clkbuf_16
X_4648_ _3850_/X _6476_/Q _4654_/S vssd1 vssd1 vccd1 vccd1 _4649_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0__2832_ clkbuf_0__2832_/X vssd1 vssd1 vccd1 vccd1 _5682__417/A sky130_fd_sc_hd__clkbuf_4
X_4579_ _4579_/A vssd1 vssd1 vccd1 vccd1 _6507_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6318_ _7132_/A _6318_/B _6318_/C vssd1 vssd1 vccd1 vccd1 _6319_/A sky130_fd_sc_hd__and3_1
X_6249_ _7006_/Q _6250_/A _6249_/C _6249_/D vssd1 vssd1 vccd1 vccd1 _6249_/X sky130_fd_sc_hd__and4_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5861__60 _5862__61/A vssd1 vssd1 vccd1 vccd1 _6846_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7093_/CLK
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5196__251 _5196__251/A vssd1 vssd1 vccd1 vccd1 _6533_/CLK sky130_fd_sc_hd__inv_2
XFILLER_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3950_ _3950_/A vssd1 vssd1 vccd1 vccd1 _6772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6064__113 _6064__113/A vssd1 vssd1 vccd1 vccd1 _6921_/CLK sky130_fd_sc_hd__inv_2
X_3881_ _6801_/Q _3880_/X _3887_/S vssd1 vssd1 vccd1 vccd1 _3882_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5620_ _5620_/A vssd1 vssd1 vccd1 vccd1 _5913_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_117_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4502_ _4502_/A _4662_/B vssd1 vssd1 vccd1 vccd1 _4518_/S sky130_fd_sc_hd__or2_2
XFILLER_104_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4433_ _4433_/A vssd1 vssd1 vccd1 vccd1 _6569_/D sky130_fd_sc_hd__clkbuf_1
X_7152_ _7152_/A vssd1 vssd1 vccd1 vccd1 _7152_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4364_ _6607_/Q _3785_/A _4366_/S vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3315_ _6775_/Q _6774_/Q _6773_/Q _3315_/D vssd1 vssd1 vccd1 vccd1 _3317_/A sky130_fd_sc_hd__and4_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7083_ _7095_/CLK _7083_/D vssd1 vssd1 vccd1 vccd1 _7083_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6109_/A vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__buf_1
X_4295_ _4295_/A vssd1 vssd1 vccd1 vccd1 _6638_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6034_ _6897_/Q _5976_/A _6013_/X vssd1 vssd1 vccd1 vccd1 _6897_/D sky130_fd_sc_hd__a21o_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _4368_/A vssd1 vssd1 vccd1 vccd1 _4205_/A sky130_fd_sc_hd__buf_4
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6936_ _6936_/CLK _6936_/D vssd1 vssd1 vccd1 vccd1 _6936_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6867_ _6867_/CLK _6867_/D vssd1 vssd1 vccd1 vccd1 _6867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6798_ _6798_/CLK _6798_/D vssd1 vssd1 vccd1 vccd1 _6798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2746_ clkbuf_0__2746_/X vssd1 vssd1 vccd1 vccd1 _5557__382/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput109 _7107_/X vssd1 vssd1 vccd1 vccd1 caravel_wb_adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4080_ _4070_/A _4070_/B _4037_/X vssd1 vssd1 vccd1 vccd1 _4081_/B sky130_fd_sc_hd__o21ai_1
Xclkbuf_1_1_0__2881_ clkbuf_0__2881_/X vssd1 vssd1 vccd1 vccd1 _5887__81/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4982_ _7082_/Q vssd1 vssd1 vccd1 vccd1 _6155_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6721_ _6721_/CLK _6721_/D vssd1 vssd1 vccd1 vccd1 _6721_/Q sky130_fd_sc_hd__dfxtp_1
X_3933_ _3933_/A vssd1 vssd1 vccd1 vccd1 _6780_/D sky130_fd_sc_hd__clkbuf_1
X_3864_ _3864_/A vssd1 vssd1 vccd1 vccd1 _6806_/D sky130_fd_sc_hd__clkbuf_1
X_6652_ _6652_/CLK _6652_/D vssd1 vssd1 vccd1 vccd1 _6652_/Q sky130_fd_sc_hd__dfxtp_1
X_5603_ _5619_/A vssd1 vssd1 vccd1 vccd1 _5664_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3795_ _3687_/X _6834_/Q _3801_/S vssd1 vssd1 vccd1 vccd1 _3796_/A sky130_fd_sc_hd__mux2_1
X_6583_ _6583_/CLK _6583_/D vssd1 vssd1 vccd1 vccd1 _6583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4416_ _3263_/X _6584_/Q _4420_/S vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__mux2_1
X_7135_ _7135_/A vssd1 vssd1 vccd1 vccd1 _7135_/X sky130_fd_sc_hd__clkbuf_1
X_5396_ _5395_/X _5435_/B vssd1 vssd1 vccd1 vccd1 _5396_/X sky130_fd_sc_hd__and2b_1
XFILLER_113_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4347_ _4347_/A vssd1 vssd1 vccd1 vccd1 _6615_/D sky130_fd_sc_hd__clkbuf_1
X_6376__4 _6376__4/A vssd1 vssd1 vccd1 vccd1 _7078_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0__2531_ clkbuf_0__2531_/X vssd1 vssd1 vccd1 vccd1 _5236__284/A sky130_fd_sc_hd__clkbuf_4
X_7066_ _7066_/CLK _7066_/D vssd1 vssd1 vccd1 vccd1 _7066_/Q sky130_fd_sc_hd__dfxtp_1
X_4278_ _4368_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4294_/S sky130_fd_sc_hd__nor2_2
XFILLER_74_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3229_ _6469_/Q _6468_/Q vssd1 vssd1 vccd1 vccd1 _5044_/A sky130_fd_sc_hd__and2b_1
X_6017_ _6017_/A vssd1 vssd1 vccd1 vccd1 _6017_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6919_ _6919_/CLK _6919_/D vssd1 vssd1 vccd1 vccd1 _6919_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3014_ clkbuf_0__3014_/X vssd1 vssd1 vccd1 vccd1 _6140_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2729_ clkbuf_0__2729_/X vssd1 vssd1 vccd1 vccd1 _5492_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5570__392 _5572__394/A vssd1 vssd1 vccd1 vccd1 _6682_/CLK sky130_fd_sc_hd__inv_2
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3580_ _3595_/S vssd1 vssd1 vccd1 vccd1 _3589_/S sky130_fd_sc_hd__buf_2
XFILLER_114_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5250_ _5250_/A vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4201_ _4201_/A vssd1 vssd1 vccd1 vccd1 _6679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4132_ _4132_/A vssd1 vssd1 vccd1 vccd1 _6710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4063_ _4063_/A vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_0__2864_ clkbuf_0__2864_/X vssd1 vssd1 vccd1 vccd1 _5806__497/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__2832_ _5679_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2832_/X sky130_fd_sc_hd__clkbuf_16
X_4965_ _6435_/Q _6695_/Q _5736_/B vssd1 vssd1 vccd1 vccd1 _4969_/B sky130_fd_sc_hd__and3_1
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3916_ _4644_/A _4168_/A vssd1 vssd1 vccd1 vccd1 _3932_/S sky130_fd_sc_hd__nor2_2
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6704_ _6704_/CLK _6704_/D vssd1 vssd1 vccd1 vccd1 _6704_/Q sky130_fd_sc_hd__dfxtp_1
X_4896_ _6903_/Q _6563_/Q _6911_/Q _6491_/Q _4806_/A _4701_/X vssd1 vssd1 vccd1 vccd1
+ _4896_/X sky130_fd_sc_hd__mux4_2
XFILLER_20_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3847_ _3869_/S vssd1 vssd1 vccd1 vccd1 _3860_/S sky130_fd_sc_hd__clkbuf_2
X_6635_ _6635_/CLK _6635_/D vssd1 vssd1 vccd1 vccd1 _6635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3778_ _3778_/A vssd1 vssd1 vccd1 vccd1 _6840_/D sky130_fd_sc_hd__clkbuf_1
X_6566_ _6566_/CLK _6566_/D vssd1 vssd1 vccd1 vccd1 _6566_/Q sky130_fd_sc_hd__dfxtp_1
X_5517_ _5523_/A vssd1 vssd1 vccd1 vccd1 _5517_/X sky130_fd_sc_hd__buf_1
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6497_ _6497_/CLK _6497_/D vssd1 vssd1 vccd1 vccd1 _6497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5031__180 _5033__182/A vssd1 vssd1 vccd1 vccd1 _6436_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5379_ _5437_/A _5379_/B vssd1 vssd1 vccd1 vccd1 _5379_/Y sky130_fd_sc_hd__nor2_1
X_7118_ _7118_/A vssd1 vssd1 vccd1 vccd1 _7118_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2514_ clkbuf_0__2514_/X vssd1 vssd1 vccd1 vccd1 _5169_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7049_ _7049_/CLK _7049_/D vssd1 vssd1 vccd1 vccd1 _7049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5676__412 _5678__414/A vssd1 vssd1 vccd1 vccd1 _6706_/CLK sky130_fd_sc_hd__inv_2
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4750_/A _4762_/D vssd1 vssd1 vccd1 vccd1 _4794_/C sky130_fd_sc_hd__nor2_1
X_3701_ _3701_/A vssd1 vssd1 vccd1 vccd1 _6891_/D sky130_fd_sc_hd__clkbuf_1
X_4681_ _4987_/A vssd1 vssd1 vccd1 vccd1 _5005_/A sky130_fd_sc_hd__clkinv_4
X_6420_ _6420_/A vssd1 vssd1 vccd1 vccd1 _7091_/D sky130_fd_sc_hd__clkbuf_1
X_3632_ _3632_/A vssd1 vssd1 vccd1 vccd1 _6918_/D sky130_fd_sc_hd__clkbuf_1
X_3563_ _3357_/X _6945_/Q _3571_/S vssd1 vssd1 vccd1 vccd1 _3564_/A sky130_fd_sc_hd__mux2_1
X_5302_ _5302_/A vssd1 vssd1 vccd1 vccd1 _5439_/B sky130_fd_sc_hd__buf_2
X_6282_ _6282_/A vssd1 vssd1 vccd1 vccd1 _6300_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3494_ _3494_/A vssd1 vssd1 vccd1 vccd1 _6975_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4115_ _6717_/Q _3886_/X _4115_/S vssd1 vssd1 vccd1 vccd1 _4116_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5095_ _5588_/S vssd1 vssd1 vccd1 vccd1 _5586_/S sky130_fd_sc_hd__buf_4
X_5577__398 _5577__398/A vssd1 vssd1 vccd1 vccd1 _6688_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4046_ _6305_/A vssd1 vssd1 vccd1 vccd1 _6303_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5997_ _6881_/Q _5966_/X _5996_/Y _5970_/X vssd1 vssd1 vccd1 vccd1 _5998_/B sky130_fd_sc_hd__a22o_1
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4948_ _4954_/S _4948_/B vssd1 vssd1 vccd1 vccd1 _4948_/X sky130_fd_sc_hd__or2_1
X_4879_ _4808_/X _4878_/X _4718_/A vssd1 vssd1 vccd1 vccd1 _4879_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_0__2746_ _5554_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2746_/X sky130_fd_sc_hd__clkbuf_16
X_6618_ _6618_/CLK _6618_/D vssd1 vssd1 vccd1 vccd1 _6618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6549_ _6549_/CLK _6549_/D vssd1 vssd1 vccd1 vccd1 _6549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5868__66 _5871__69/A vssd1 vssd1 vccd1 vccd1 _6852_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5521__353 _5522__354/A vssd1 vssd1 vccd1 vccd1 _6643_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6152__9 _6152__9/A vssd1 vssd1 vccd1 vccd1 _6992_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5190__246 _5190__246/A vssd1 vssd1 vccd1 vccd1 _6528_/CLK sky130_fd_sc_hd__inv_2
X_6348__34 _6348__34/A vssd1 vssd1 vccd1 vccd1 _7054_/CLK sky130_fd_sc_hd__inv_2
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5920_ _5915_/X _5916_/Y _5917_/X _5919_/Y vssd1 vssd1 vccd1 vccd1 _5921_/D sky130_fd_sc_hd__a211o_1
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4802_ _4802_/A vssd1 vssd1 vccd1 vccd1 _4802_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4733_ _4729_/X _4731_/X _4905_/A vssd1 vssd1 vccd1 vccd1 _4733_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2531_ _5231_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2531_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4664_ _3845_/X _6443_/Q _4672_/S vssd1 vssd1 vccd1 vccd1 _4665_/A sky130_fd_sc_hd__mux2_1
X_6403_ _6403_/A vssd1 vssd1 vccd1 vccd1 _7086_/D sky130_fd_sc_hd__clkbuf_1
X_4595_ _4595_/A vssd1 vssd1 vccd1 vccd1 _6500_/D sky130_fd_sc_hd__clkbuf_1
X_5464__307 _5464__307/A vssd1 vssd1 vccd1 vccd1 _6597_/CLK sky130_fd_sc_hd__inv_2
X_3615_ _6924_/Q _3614_/X _3621_/S vssd1 vssd1 vccd1 vccd1 _3616_/A sky130_fd_sc_hd__mux2_1
X_3546_ _3546_/A vssd1 vssd1 vccd1 vccd1 _6953_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6265_ _6266_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6267_/B sky130_fd_sc_hd__or2_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3477_ _3477_/A vssd1 vssd1 vccd1 vccd1 _6981_/D sky130_fd_sc_hd__clkbuf_1
X_6196_ _6207_/C vssd1 vssd1 vccd1 vccd1 _6196_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3014_ _6115_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3014_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5078_ _6456_/Q _7110_/A _5082_/S vssd1 vssd1 vccd1 vccd1 _5079_/A sky130_fd_sc_hd__mux2_1
X_4029_ _4029_/A vssd1 vssd1 vccd1 vccd1 _4029_/X sky130_fd_sc_hd__clkbuf_4
X_5813__503 _5813__503/A vssd1 vssd1 vccd1 vccd1 _6809_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2729_ _5467_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2729_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_119_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3400_ _4590_/A _4626_/A vssd1 vssd1 vccd1 vccd1 _3416_/S sky130_fd_sc_hd__or2_2
X_4380_ _6600_/Q _3782_/A _4384_/S vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__mux2_1
X_5528__359 _5528__359/A vssd1 vssd1 vccd1 vccd1 _6649_/CLK sky130_fd_sc_hd__inv_2
X_3331_ _3331_/A vssd1 vssd1 vccd1 vccd1 _7061_/D sky130_fd_sc_hd__clkbuf_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3262_/A vssd1 vssd1 vccd1 vccd1 _7074_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5001_ _5003_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _5002_/A sky130_fd_sc_hd__and2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6952_ _6952_/CLK _6952_/D vssd1 vssd1 vccd1 vccd1 _6952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5903_ _5892_/B _5623_/B _6879_/Q vssd1 vssd1 vccd1 vccd1 _5921_/B sky130_fd_sc_hd__a21oi_1
X_6883_ _6883_/CLK _6883_/D vssd1 vssd1 vccd1 vccd1 _6883_/Q sky130_fd_sc_hd__dfxtp_1
X_5834_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5834_/X sky130_fd_sc_hd__buf_1
X_5470__311 _5470__311/A vssd1 vssd1 vccd1 vccd1 _6601_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4716_ _4716_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4716_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_0__2514_ _5144_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2514_/X sky130_fd_sc_hd__clkbuf_16
X_4647_ _4647_/A vssd1 vssd1 vccd1 vccd1 _6477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4578_ _4484_/X _6507_/Q _4582_/S vssd1 vssd1 vccd1 vccd1 _4579_/A sky130_fd_sc_hd__mux2_1
X_6317_ _6317_/A vssd1 vssd1 vccd1 vccd1 _7029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3529_ _3529_/A vssd1 vssd1 vccd1 vccd1 _6960_/D sky130_fd_sc_hd__clkbuf_1
X_6248_ _6248_/A vssd1 vssd1 vccd1 vccd1 _7005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6179_ _6172_/X _6175_/X _6178_/X _6994_/Q vssd1 vssd1 vccd1 vccd1 _6179_/X sky130_fd_sc_hd__o31a_1
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5141__207 _5143__209/A vssd1 vssd1 vccd1 vccd1 _6489_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5534__363 _5534__363/A vssd1 vssd1 vccd1 vccd1 _6653_/CLK sky130_fd_sc_hd__inv_2
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3880_ _6746_/Q vssd1 vssd1 vccd1 vccd1 _3880_/X sky130_fd_sc_hd__buf_2
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4501_ _4501_/A vssd1 vssd1 vccd1 vccd1 _6542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4432_ _3260_/X _6569_/Q _4432_/S vssd1 vssd1 vccd1 vccd1 _4433_/A sky130_fd_sc_hd__mux2_1
X_7151_ _7151_/A vssd1 vssd1 vccd1 vccd1 _7151_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4363_ _4363_/A vssd1 vssd1 vccd1 vccd1 _6608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3314_ _3485_/A _3962_/A vssd1 vssd1 vccd1 vccd1 _3318_/C sky130_fd_sc_hd__xnor2_1
X_7082_ _7095_/CLK _7082_/D vssd1 vssd1 vccd1 vccd1 _7082_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _6638_/Q _4164_/X _4294_/S vssd1 vssd1 vccd1 vccd1 _4295_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3361_/A _4051_/A _3418_/C vssd1 vssd1 vccd1 vccd1 _4368_/A sky130_fd_sc_hd__or3_4
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5205__259 _5205__259/A vssd1 vssd1 vccd1 vccd1 _6541_/CLK sky130_fd_sc_hd__inv_2
XFILLER_66_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6935_ _6935_/CLK _6935_/D vssd1 vssd1 vccd1 vccd1 _6935_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6866_ _6866_/CLK _6866_/D vssd1 vssd1 vccd1 vccd1 _6866_/Q sky130_fd_sc_hd__dfxtp_1
X_6797_ _6797_/CLK _6797_/D vssd1 vssd1 vccd1 vccd1 _6797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2529_ clkbuf_0__2529_/X vssd1 vssd1 vccd1 vccd1 _5223__273/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5679_ _5697_/A vssd1 vssd1 vccd1 vccd1 _5679_/X sky130_fd_sc_hd__buf_1
XFILLER_116_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__2745_ clkbuf_0__2745_/X vssd1 vssd1 vccd1 vccd1 _5550__376/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5477__317 _5478__318/A vssd1 vssd1 vccd1 vccd1 _6607_/CLK sky130_fd_sc_hd__inv_2
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__3159_ clkbuf_0__3159_/X vssd1 vssd1 vccd1 vccd1 _6370__52/A sky130_fd_sc_hd__clkbuf_4
X_5826__513 _5827__514/A vssd1 vssd1 vccd1 vccd1 _6819_/CLK sky130_fd_sc_hd__inv_2
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2880_ clkbuf_0__2880_/X vssd1 vssd1 vccd1 vccd1 _6028_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _4973_/X input7/X _4970_/X _6170_/A vssd1 vssd1 vccd1 vccd1 _4981_/X sky130_fd_sc_hd__a22o_2
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6720_ _6720_/CLK _6720_/D vssd1 vssd1 vccd1 vccd1 _6720_/Q sky130_fd_sc_hd__dfxtp_1
X_3932_ _6780_/Q _3895_/X _3932_/S vssd1 vssd1 vccd1 vccd1 _3933_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3863_ _6806_/Q _3862_/X _3869_/S vssd1 vssd1 vccd1 vccd1 _3864_/A sky130_fd_sc_hd__mux2_1
X_6651_ _6651_/CLK _6651_/D vssd1 vssd1 vccd1 vccd1 _6651_/Q sky130_fd_sc_hd__dfxtp_1
X_5602_ _7095_/Q _7094_/Q _7093_/Q _7092_/Q vssd1 vssd1 vccd1 vccd1 _5619_/A sky130_fd_sc_hd__or4_1
X_6582_ _6582_/CLK _6582_/D vssd1 vssd1 vccd1 vccd1 _6582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3794_ _3794_/A vssd1 vssd1 vccd1 vccd1 _6835_/D sky130_fd_sc_hd__clkbuf_1
X_5211__263 _5212__264/A vssd1 vssd1 vccd1 vccd1 _6545_/CLK sky130_fd_sc_hd__inv_2
X_4415_ _4415_/A vssd1 vssd1 vccd1 vccd1 _6585_/D sky130_fd_sc_hd__clkbuf_1
X_5395_ _6793_/Q _6983_/Q _6991_/Q _6967_/Q _5341_/A _5276_/X vssd1 vssd1 vccd1 vccd1
+ _5395_/X sky130_fd_sc_hd__mux4_2
X_7134_ _7134_/A vssd1 vssd1 vccd1 vccd1 _7134_/X sky130_fd_sc_hd__clkbuf_1
X_4346_ _3785_/X _6615_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__mux2_1
XFILLER_100_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2530_ clkbuf_0__2530_/X vssd1 vssd1 vccd1 vccd1 _5229__278/A sky130_fd_sc_hd__clkbuf_4
X_7065_ _7065_/CLK _7065_/D vssd1 vssd1 vccd1 vccd1 _7065_/Q sky130_fd_sc_hd__dfxtp_1
X_4277_ _4277_/A _4277_/B _4277_/C vssd1 vssd1 vccd1 vccd1 _4350_/B sky130_fd_sc_hd__nand3_4
XFILLER_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3228_ _6749_/Q _5043_/B vssd1 vssd1 vccd1 vccd1 _4051_/B sky130_fd_sc_hd__and2_1
X_6016_ _5924_/D _5926_/B _6015_/X vssd1 vssd1 vccd1 vccd1 _6021_/B sky130_fd_sc_hd__a21oi_1
XFILLER_54_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6918_ _6918_/CLK _6918_/D vssd1 vssd1 vccd1 vccd1 _6918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6849_ _6849_/CLK _6849_/D vssd1 vssd1 vccd1 vccd1 _6849_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3013_ clkbuf_0__3013_/X vssd1 vssd1 vccd1 vccd1 _6113__153/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2728_ clkbuf_0__2728_/X vssd1 vssd1 vccd1 vccd1 _5464__307/A sky130_fd_sc_hd__clkbuf_4
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5154__217 _5155__218/A vssd1 vssd1 vccd1 vccd1 _6499_/CLK sky130_fd_sc_hd__inv_2
XFILLER_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4200_ _6679_/Q _4161_/X _4202_/S vssd1 vssd1 vccd1 vccd1 _4201_/A sky130_fd_sc_hd__mux2_1
XFILLER_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4131_ _6710_/Q _3883_/X _4133_/S vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4062_ _5341_/A vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__clkbuf_8
Xclkbuf_1_1_0__2863_ clkbuf_0__2863_/X vssd1 vssd1 vccd1 vccd1 _5802__494/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4964_ _4888_/X input32/X _4695_/X _4963_/X vssd1 vssd1 vccd1 vccd1 _4964_/X sky130_fd_sc_hd__a22o_2
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6703_ _6703_/CLK _6703_/D vssd1 vssd1 vccd1 vccd1 _6703_/Q sky130_fd_sc_hd__dfxtp_1
X_3915_ _3915_/A vssd1 vssd1 vccd1 vccd1 _6788_/D sky130_fd_sc_hd__clkbuf_1
X_4895_ _4774_/X _4894_/X _4865_/A vssd1 vssd1 vccd1 vccd1 _4895_/X sky130_fd_sc_hd__a21o_1
X_3846_ _4590_/A _3873_/B vssd1 vssd1 vccd1 vccd1 _3869_/S sky130_fd_sc_hd__nor2_2
X_6634_ _6634_/CLK _6634_/D vssd1 vssd1 vccd1 vccd1 _6634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6565_ _6565_/CLK _6565_/D vssd1 vssd1 vccd1 vccd1 _6565_/Q sky130_fd_sc_hd__dfxtp_1
X_3777_ _3776_/X _6840_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__mux2_1
X_6496_ _6496_/CLK _6496_/D vssd1 vssd1 vccd1 vccd1 _6496_/Q sky130_fd_sc_hd__dfxtp_1
X_6077__124 _6077__124/A vssd1 vssd1 vccd1 vccd1 _6932_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5378_ _6950_/Q _6682_/Q _6594_/Q _6816_/Q _5337_/X _5338_/X vssd1 vssd1 vccd1 vccd1
+ _5379_/B sky130_fd_sc_hd__mux4_2
X_7117_ _7117_/A vssd1 vssd1 vccd1 vccd1 _7117_/X sky130_fd_sc_hd__clkbuf_1
X_4329_ _4329_/A vssd1 vssd1 vccd1 vccd1 _6623_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2513_ clkbuf_0__2513_/X vssd1 vssd1 vccd1 vccd1 _5140__206/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7048_ _7048_/CLK _7048_/D vssd1 vssd1 vccd1 vccd1 _7048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5218__269 _5218__269/A vssd1 vssd1 vccd1 vccd1 _6551_/CLK sky130_fd_sc_hd__inv_2
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3699_/X _6891_/Q _3706_/S vssd1 vssd1 vccd1 vccd1 _3701_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ _6435_/Q vssd1 vssd1 vccd1 vccd1 _4987_/A sky130_fd_sc_hd__buf_6
X_5119__189 _5119__189/A vssd1 vssd1 vccd1 vccd1 _6471_/CLK sky130_fd_sc_hd__inv_2
X_3631_ _3376_/X _6918_/Q _3633_/S vssd1 vssd1 vccd1 vccd1 _3632_/A sky130_fd_sc_hd__mux2_1
X_3562_ _3577_/S vssd1 vssd1 vccd1 vccd1 _3571_/S sky130_fd_sc_hd__buf_2
X_5301_ _5300_/X _5351_/B vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__and2b_1
X_6281_ _6995_/Q _6272_/A _6280_/X _7014_/Q _6247_/A vssd1 vssd1 vccd1 vccd1 _7014_/D
+ sky130_fd_sc_hd__o221a_1
X_3493_ _3333_/X _6975_/Q _3497_/S vssd1 vssd1 vccd1 vccd1 _3494_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5163_ _5163_/A vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__buf_1
X_4114_ _4114_/A vssd1 vssd1 vccd1 vccd1 _6718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5094_ _5094_/A vssd1 vssd1 vccd1 vccd1 _6463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4045_ _4277_/C _4049_/B _4044_/X _4037_/X vssd1 vssd1 vccd1 vccd1 _6737_/D sky130_fd_sc_hd__o211a_1
XFILLER_71_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _6004_/C _5996_/B vssd1 vssd1 vccd1 vccd1 _5996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4947_ _6477_/Q _6629_/Q _7062_/Q _6787_/Q _4719_/X _4772_/S vssd1 vssd1 vccd1 vccd1
+ _4948_/B sky130_fd_sc_hd__mux4_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4878_ _6893_/Q _6522_/Q _4878_/S vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_0__2745_ _5548_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2745_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_20_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3829_ _6819_/Q _3597_/X _3837_/S vssd1 vssd1 vccd1 vccd1 _3830_/A sky130_fd_sc_hd__mux2_1
X_6617_ _6617_/CLK _6617_/D vssd1 vssd1 vccd1 vccd1 _6617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6548_ _6548_/CLK _6548_/D vssd1 vssd1 vccd1 vccd1 _6548_/Q sky130_fd_sc_hd__dfxtp_1
X_6479_ _6479_/CLK _6479_/D vssd1 vssd1 vccd1 vccd1 _6479_/Q sky130_fd_sc_hd__dfxtp_1
XINSDIODE2_0 _3614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__3159_ _6367_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3159_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4801_ _7094_/Q vssd1 vssd1 vccd1 vccd1 _5910_/A sky130_fd_sc_hd__clkbuf_4
X_4732_ _4732_/A vssd1 vssd1 vccd1 vccd1 _4905_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__2530_ _5225_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2530_/X sky130_fd_sc_hd__clkbuf_16
X_4663_ _4678_/S vssd1 vssd1 vccd1 vccd1 _4672_/S sky130_fd_sc_hd__buf_2
XFILLER_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6402_ _6408_/A _6402_/B vssd1 vssd1 vccd1 vccd1 _6403_/A sky130_fd_sc_hd__and2_1
X_3614_ _7025_/Q vssd1 vssd1 vccd1 vccd1 _3614_/X sky130_fd_sc_hd__buf_4
X_4594_ _6500_/Q _4014_/A _4600_/S vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__mux2_1
X_3545_ _6953_/Q _3437_/X _3553_/S vssd1 vssd1 vccd1 vccd1 _3546_/A sky130_fd_sc_hd__mux2_1
X_6264_ _6264_/A vssd1 vssd1 vccd1 vccd1 _7009_/D sky130_fd_sc_hd__clkbuf_1
X_3476_ _3380_/X _6981_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3477_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6195_ _6216_/C _6254_/C vssd1 vssd1 vccd1 vccd1 _6207_/C sky130_fd_sc_hd__and2_1
Xclkbuf_0__3013_ _6109_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3013_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5873__70 _5876__73/A vssd1 vssd1 vccd1 vccd1 _6856_/CLK sky130_fd_sc_hd__inv_2
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5077_ _5077_/A vssd1 vssd1 vccd1 vccd1 _6455_/D sky130_fd_sc_hd__clkbuf_1
X_4028_ _4028_/A vssd1 vssd1 vccd1 vccd1 _6753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5979_ _6877_/Q _5978_/C _6878_/Q vssd1 vssd1 vccd1 vccd1 _5980_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_0__2728_ _5461_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2728_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3330_ _3329_/X _7061_/Q _3342_/S vssd1 vssd1 vccd1 vccd1 _3331_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5000_ _5000_/A vssd1 vssd1 vccd1 vccd1 _5000_/X sky130_fd_sc_hd__clkbuf_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _7074_/Q _3260_/X _3261_/S vssd1 vssd1 vccd1 vccd1 _3262_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6951_ _6951_/CLK _6951_/D vssd1 vssd1 vccd1 vccd1 _6951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5902_ _6881_/Q _5902_/B vssd1 vssd1 vccd1 vccd1 _5921_/A sky130_fd_sc_hd__xnor2_1
X_6882_ _6883_/CLK _6882_/D vssd1 vssd1 vccd1 vccd1 _6882_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5689__423 _5690__424/A vssd1 vssd1 vccd1 vccd1 _6717_/CLK sky130_fd_sc_hd__inv_2
XFILLER_62_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4715_ _6502_/Q _6436_/Q _6534_/Q _6686_/Q _4936_/S _3959_/A vssd1 vssd1 vccd1 vccd1
+ _4716_/B sky130_fd_sc_hd__mux4_2
XFILLER_108_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2513_ _5138_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2513_/X sky130_fd_sc_hd__clkbuf_16
X_4646_ _3845_/X _6477_/Q _4654_/S vssd1 vssd1 vccd1 vccd1 _4647_/A sky130_fd_sc_hd__mux2_1
X_4577_ _4577_/A vssd1 vssd1 vccd1 vccd1 _6508_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6316_ _7131_/A _6318_/B _6318_/C vssd1 vssd1 vccd1 vccd1 _6317_/A sky130_fd_sc_hd__and3_1
XFILLER_115_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3528_ _6960_/Q _3444_/X _3534_/S vssd1 vssd1 vccd1 vccd1 _3529_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6247_ _6247_/A _6247_/B vssd1 vssd1 vccd1 vccd1 _6248_/A sky130_fd_sc_hd__and2_1
X_3459_ _3785_/A vssd1 vssd1 vccd1 vccd1 _3459_/X sky130_fd_sc_hd__clkbuf_2
X_6178_ _6178_/A _6178_/B _6177_/X vssd1 vssd1 vccd1 vccd1 _6178_/X sky130_fd_sc_hd__or3b_1
XFILLER_29_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4500_ _4499_/X _6542_/Q _4500_/S vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__mux2_1
X_5480_ _5486_/A vssd1 vssd1 vccd1 vccd1 _5480_/X sky130_fd_sc_hd__buf_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4431_ _4431_/A vssd1 vssd1 vccd1 vccd1 _6570_/D sky130_fd_sc_hd__clkbuf_1
X_7150_ _7150_/A vssd1 vssd1 vccd1 vccd1 _7150_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4362_ _6608_/Q _3782_/A _4366_/S vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3313_ _6774_/Q _6769_/Q vssd1 vssd1 vccd1 vccd1 _3962_/A sky130_fd_sc_hd__xor2_1
X_7081_ _7095_/CLK _7081_/D vssd1 vssd1 vccd1 vccd1 _7081_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071__119 _6071__119/A vssd1 vssd1 vccd1 vccd1 _6927_/CLK sky130_fd_sc_hd__inv_2
X_4293_ _4293_/A vssd1 vssd1 vccd1 vccd1 _6639_/D sky130_fd_sc_hd__clkbuf_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _4051_/B _4036_/A vssd1 vssd1 vccd1 vccd1 _3418_/C sky130_fd_sc_hd__nand2_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6934_ _6934_/CLK _6934_/D vssd1 vssd1 vccd1 vccd1 _6934_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6865_ _6865_/CLK _6865_/D vssd1 vssd1 vccd1 vccd1 _6865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6796_ _6796_/CLK _6796_/D vssd1 vssd1 vccd1 vccd1 _6796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2528_ clkbuf_0__2528_/X vssd1 vssd1 vccd1 vccd1 _5216__267/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4629_ _4629_/A vssd1 vssd1 vccd1 vccd1 _6485_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0_0__2744_ clkbuf_0__2744_/X vssd1 vssd1 vccd1 vccd1 _5547__374/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5600__410 _5601__411/A vssd1 vssd1 vccd1 vccd1 _6703_/CLK sky130_fd_sc_hd__inv_2
XFILLER_103_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__3158_ clkbuf_0__3158_/X vssd1 vssd1 vccd1 vccd1 _6366__49/A sky130_fd_sc_hd__clkbuf_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _7083_/Q vssd1 vssd1 vccd1 vccd1 _6170_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3931_ _3931_/A vssd1 vssd1 vccd1 vccd1 _6781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3862_ _6743_/Q vssd1 vssd1 vccd1 vccd1 _3862_/X sky130_fd_sc_hd__buf_4
X_6650_ _6650_/CLK _6650_/D vssd1 vssd1 vccd1 vccd1 _6650_/Q sky130_fd_sc_hd__dfxtp_1
X_6581_ _6888_/CLK _6581_/D vssd1 vssd1 vccd1 vccd1 _6581_/Q sky130_fd_sc_hd__dfxtp_1
X_3793_ _3680_/X _6835_/Q _3801_/S vssd1 vssd1 vccd1 vccd1 _3794_/A sky130_fd_sc_hd__mux2_1
X_5582__402 _5583__403/A vssd1 vssd1 vccd1 vccd1 _6692_/CLK sky130_fd_sc_hd__inv_2
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4414_ _3260_/X _6585_/Q _4414_/S vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__mux2_1
X_5394_ _5390_/X _5393_/X _5394_/S vssd1 vssd1 vccd1 vccd1 _5394_/X sky130_fd_sc_hd__mux2_1
X_7133_ _7133_/A vssd1 vssd1 vccd1 vccd1 _7133_/X sky130_fd_sc_hd__clkbuf_1
X_4345_ _4345_/A vssd1 vssd1 vccd1 vccd1 _6616_/D sky130_fd_sc_hd__clkbuf_1
X_6320__11 _6323__14/A vssd1 vssd1 vccd1 vccd1 _7031_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7064_ _7064_/CLK _7064_/D vssd1 vssd1 vccd1 vccd1 _7064_/Q sky130_fd_sc_hd__dfxtp_1
X_4276_ _4276_/A vssd1 vssd1 vccd1 vccd1 _6646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6015_ _6868_/Q _6015_/B _6886_/Q vssd1 vssd1 vccd1 vccd1 _6015_/X sky130_fd_sc_hd__or3b_1
X_3227_ _3227_/A _3227_/B _3227_/C _3226_/X vssd1 vssd1 vccd1 vccd1 _5043_/B sky130_fd_sc_hd__or4b_2
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6917_ _6917_/CLK _6917_/D vssd1 vssd1 vccd1 vccd1 _6917_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3012_ clkbuf_0__3012_/X vssd1 vssd1 vccd1 vccd1 _6108__149/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6848_ _6848_/CLK _6848_/D vssd1 vssd1 vccd1 vccd1 _6848_/Q sky130_fd_sc_hd__dfxtp_1
X_6779_ _7096_/CLK _6779_/D vssd1 vssd1 vccd1 vccd1 _6779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5483__322 _5483__322/A vssd1 vssd1 vccd1 vccd1 _6612_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2727_ clkbuf_0__2727_/X vssd1 vssd1 vccd1 vccd1 _5460__304/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6141__175 _6143__177/A vssd1 vssd1 vccd1 vccd1 _6983_/CLK sky130_fd_sc_hd__inv_2
X_4130_ _4130_/A vssd1 vssd1 vccd1 vccd1 _6711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4061_ _5258_/A vssd1 vssd1 vccd1 vccd1 _5341_/A sky130_fd_sc_hd__buf_2
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2862_ clkbuf_0__2862_/X vssd1 vssd1 vccd1 vccd1 _5795__488/A sky130_fd_sc_hd__clkbuf_4
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4963_ _4856_/Y _4951_/X _4961_/X _4987_/C _6167_/A vssd1 vssd1 vccd1 vccd1 _4963_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6702_ _6702_/CLK _6702_/D vssd1 vssd1 vccd1 vccd1 _6702_/Q sky130_fd_sc_hd__dfxtp_1
X_3914_ _6788_/Q _3620_/X _3914_/S vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__mux2_1
X_4894_ _6483_/Q _6555_/Q _4900_/S vssd1 vssd1 vccd1 vccd1 _4894_/X sky130_fd_sc_hd__mux2_1
X_6633_ _6633_/CLK _6633_/D vssd1 vssd1 vccd1 vccd1 _6633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3845_ _6748_/Q vssd1 vssd1 vccd1 vccd1 _3845_/X sky130_fd_sc_hd__buf_6
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6564_ _6564_/CLK _6564_/D vssd1 vssd1 vccd1 vccd1 _6564_/Q sky130_fd_sc_hd__dfxtp_1
X_3776_ _3776_/A vssd1 vssd1 vccd1 vccd1 _3776_/X sky130_fd_sc_hd__clkbuf_2
X_6495_ _6495_/CLK _6495_/D vssd1 vssd1 vccd1 vccd1 _6495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5547__374 _5547__374/A vssd1 vssd1 vccd1 vccd1 _6664_/CLK sky130_fd_sc_hd__inv_2
XFILLER_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5377_ _5376_/X _5435_/B vssd1 vssd1 vccd1 vccd1 _5377_/X sky130_fd_sc_hd__and2b_1
X_7116_ _7116_/A vssd1 vssd1 vccd1 vccd1 _7116_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4328_ _6623_/Q _3892_/X _4330_/S vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_0__2512_ clkbuf_0__2512_/X vssd1 vssd1 vccd1 vccd1 _5136__203/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4259_ _4350_/A _4259_/B vssd1 vssd1 vccd1 vccd1 _4275_/S sky130_fd_sc_hd__nor2_2
X_7047_ _7047_/CLK _7047_/D vssd1 vssd1 vccd1 vccd1 _7047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5448__294 _5448__294/A vssd1 vssd1 vccd1 vccd1 _6584_/CLK sky130_fd_sc_hd__inv_2
XFILLER_111_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5160__222 _5160__222/A vssd1 vssd1 vccd1 vccd1 _6504_/CLK sky130_fd_sc_hd__inv_2
XFILLER_93_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5683__418 _5684__419/A vssd1 vssd1 vccd1 vccd1 _6712_/CLK sky130_fd_sc_hd__inv_2
X_3630_ _3630_/A vssd1 vssd1 vccd1 vccd1 _6919_/D sky130_fd_sc_hd__clkbuf_1
X_3561_ _3579_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _3577_/S sky130_fd_sc_hd__or2_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5300_ _6789_/Q _6979_/Q _6987_/Q _6963_/Q _5290_/X _4069_/A vssd1 vssd1 vccd1 vccd1
+ _5300_/X sky130_fd_sc_hd__mux4_1
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6280_ _6271_/X _6280_/B _7013_/Q _7012_/Q vssd1 vssd1 vccd1 vccd1 _6280_/X sky130_fd_sc_hd__and4b_1
X_3492_ _3492_/A vssd1 vssd1 vccd1 vccd1 _6976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5231_ _5231_/A vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__buf_1
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5839__524 _5839__524/A vssd1 vssd1 vccd1 vccd1 _6830_/CLK sky130_fd_sc_hd__inv_2
X_4113_ _6718_/Q _3883_/X _4115_/S vssd1 vssd1 vccd1 vccd1 _4114_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5093_ _6463_/Q _7117_/A _5093_/S vssd1 vssd1 vccd1 vccd1 _5094_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4044_ _4044_/A _4044_/B vssd1 vssd1 vccd1 vccd1 _4044_/X sky130_fd_sc_hd__or2_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5995_ _5994_/B _5994_/C _6881_/Q vssd1 vssd1 vccd1 vccd1 _5996_/B sky130_fd_sc_hd__a21oi_1
X_4946_ _4927_/A _4945_/X _4802_/X vssd1 vssd1 vccd1 vccd1 _4946_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _3986_/A _6514_/Q _4876_/X _4728_/X vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__o211a_1
Xclkbuf_0__2744_ _5542_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2744_/X sky130_fd_sc_hd__clkbuf_16
X_3828_ _3843_/S vssd1 vssd1 vccd1 vccd1 _3837_/S sky130_fd_sc_hd__clkbuf_2
X_6616_ _6616_/CLK _6616_/D vssd1 vssd1 vccd1 vccd1 _6616_/Q sky130_fd_sc_hd__dfxtp_1
X_6547_ _6547_/CLK _6547_/D vssd1 vssd1 vccd1 vccd1 _6547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3759_ _3759_/A vssd1 vssd1 vccd1 vccd1 _6846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6478_ _6478_/CLK _6478_/D vssd1 vssd1 vccd1 vccd1 _6478_/Q sky130_fd_sc_hd__dfxtp_1
X_5429_ _5427_/X _5428_/X _5429_/S vssd1 vssd1 vccd1 vccd1 _5429_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_1 _3845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__3158_ _6361_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3158_/X sky130_fd_sc_hd__clkbuf_16
X_5224__274 _5224__274/A vssd1 vssd1 vccd1 vccd1 _6556_/CLK sky130_fd_sc_hd__inv_2
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5125__194 _5125__194/A vssd1 vssd1 vccd1 vccd1 _6476_/CLK sky130_fd_sc_hd__inv_2
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_wb_clk_i clkbuf_4_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _7030_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_4800_ _4691_/X input14/X _4764_/X _4799_/X vssd1 vssd1 vccd1 vccd1 _4800_/X sky130_fd_sc_hd__a22o_2
XFILLER_22_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _6898_/Q _6558_/Q _6906_/Q _6486_/Q _3958_/A _4956_/S vssd1 vssd1 vccd1 vccd1
+ _4731_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4662_ _4662_/A _4662_/B vssd1 vssd1 vccd1 vccd1 _4678_/S sky130_fd_sc_hd__or2_2
XFILLER_9_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6354__39 _6354__39/A vssd1 vssd1 vccd1 vccd1 _7059_/CLK sky130_fd_sc_hd__inv_2
X_6401_ _7135_/A _4974_/X _6401_/S vssd1 vssd1 vccd1 vccd1 _6402_/B sky130_fd_sc_hd__mux2_1
X_3613_ _3613_/A vssd1 vssd1 vccd1 vccd1 _6925_/D sky130_fd_sc_hd__clkbuf_1
X_4593_ _4593_/A vssd1 vssd1 vccd1 vccd1 _6501_/D sky130_fd_sc_hd__clkbuf_1
X_3544_ _3559_/S vssd1 vssd1 vccd1 vccd1 _3553_/S sky130_fd_sc_hd__clkbuf_2
X_5167__228 _5168__229/A vssd1 vssd1 vccd1 vccd1 _6510_/CLK sky130_fd_sc_hd__inv_2
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6263_ _6266_/B _6267_/A _6263_/C vssd1 vssd1 vccd1 vccd1 _6264_/A sky130_fd_sc_hd__and3b_1
X_3475_ _3475_/A vssd1 vssd1 vccd1 vccd1 _6982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6194_ _6995_/Q _6994_/Q vssd1 vssd1 vccd1 vccd1 _6254_/C sky130_fd_sc_hd__nand2_1
Xclkbuf_0__3012_ _6103_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3012_/X sky130_fd_sc_hd__clkbuf_16
X_5145_ _5169_/A vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__buf_1
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _6455_/Q _7109_/A _5082_/S vssd1 vssd1 vccd1 vccd1 _5077_/A sky130_fd_sc_hd__mux2_1
X_4027_ _4026_/X _6753_/Q _4033_/S vssd1 vssd1 vccd1 vccd1 _4028_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5978_ _6878_/Q _6877_/Q _5978_/C vssd1 vssd1 vccd1 vccd1 _5985_/B sky130_fd_sc_hd__and3_1
X_4929_ _3968_/A _4928_/X _4782_/X vssd1 vssd1 vccd1 vccd1 _4929_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2727_ _5455_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2727_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_118_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5820__509 _5820__509/A vssd1 vssd1 vccd1 vccd1 _6815_/CLK sky130_fd_sc_hd__inv_2
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3260_ _7026_/Q vssd1 vssd1 vccd1 vccd1 _3260_/X sky130_fd_sc_hd__buf_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6950_ _6950_/CLK _6950_/D vssd1 vssd1 vccd1 vccd1 _6950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2836_ clkbuf_0__2836_/X vssd1 vssd1 vccd1 vccd1 _5716_/A sky130_fd_sc_hd__clkbuf_16
X_5901_ _6879_/Q _5623_/X _5897_/Y _5898_/X _5900_/Y vssd1 vssd1 vccd1 vccd1 _5922_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6881_ _7008_/CLK _6881_/D vssd1 vssd1 vccd1 vccd1 _6881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5763_ _5784_/A vssd1 vssd1 vccd1 vccd1 _5763_/X sky130_fd_sc_hd__buf_1
X_4714_ _4876_/A vssd1 vssd1 vccd1 vccd1 _4936_/S sky130_fd_sc_hd__clkbuf_4
X_6327__17 _6328__18/A vssd1 vssd1 vccd1 vccd1 _7037_/CLK sky130_fd_sc_hd__inv_2
XFILLER_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2512_ _5132_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2512_/X sky130_fd_sc_hd__clkbuf_16
X_4645_ _4660_/S vssd1 vssd1 vccd1 vccd1 _4654_/S sky130_fd_sc_hd__buf_2
X_4576_ _4481_/X _6508_/Q _4582_/S vssd1 vssd1 vccd1 vccd1 _4577_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3527_ _3527_/A vssd1 vssd1 vccd1 vccd1 _6961_/D sky130_fd_sc_hd__clkbuf_1
X_6315_ _6315_/A vssd1 vssd1 vccd1 vccd1 _7028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6246_ _6187_/B _6243_/X _6244_/Y _6245_/Y _6250_/A vssd1 vssd1 vccd1 vccd1 _6247_/B
+ sky130_fd_sc_hd__a32o_1
X_3458_ _3458_/A vssd1 vssd1 vccd1 vccd1 _6988_/D sky130_fd_sc_hd__clkbuf_1
X_6177_ _6167_/Y _6241_/C _5648_/X _5649_/X _6269_/A vssd1 vssd1 vccd1 vccd1 _6177_/X
+ sky130_fd_sc_hd__o2111a_1
X_3389_ _3388_/X _7048_/Q _3393_/S vssd1 vssd1 vccd1 vccd1 _3390_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5059_ _6448_/Q _7102_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5060_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6105__146 _6108__149/A vssd1 vssd1 vccd1 vccd1 _6954_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4430_ _3257_/X _6570_/Q _4432_/S vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4361_/A vssd1 vssd1 vccd1 vccd1 _6609_/D sky130_fd_sc_hd__clkbuf_1
X_3312_ _3661_/A _3315_/D vssd1 vssd1 vccd1 vccd1 _3485_/A sky130_fd_sc_hd__nand2_1
X_7080_ _7089_/CLK _7080_/D vssd1 vssd1 vccd1 vccd1 _7080_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _6639_/Q _4161_/X _4294_/S vssd1 vssd1 vccd1 vccd1 _4293_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3243_ _7128_/A _3242_/X _5047_/A vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__a21oi_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5541__369 _5541__369/A vssd1 vssd1 vccd1 vccd1 _6659_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6933_ _6933_/CLK _6933_/D vssd1 vssd1 vccd1 vccd1 _6933_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6864_ _6864_/CLK _6864_/D vssd1 vssd1 vccd1 vccd1 _6864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5815_ _5815_/A vssd1 vssd1 vccd1 vccd1 _5815_/X sky130_fd_sc_hd__buf_1
XFILLER_50_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6795_ _6795_/CLK _6795_/D vssd1 vssd1 vccd1 vccd1 _6795_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1_0__2527_ clkbuf_0__2527_/X vssd1 vssd1 vccd1 vccd1 _5210__262/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2458_ clkbuf_0__2458_/X vssd1 vssd1 vccd1 vccd1 _5040__187/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4628_ _3845_/X _6485_/Q _4636_/S vssd1 vssd1 vccd1 vccd1 _4629_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4559_ _4559_/A vssd1 vssd1 vccd1 vccd1 _6516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2743_ clkbuf_0__2743_/X vssd1 vssd1 vccd1 vccd1 _5538__366/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6229_ _6237_/C _6229_/B _6229_/C vssd1 vssd1 vccd1 vccd1 _6230_/A sky130_fd_sc_hd__and3b_1
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3157_ clkbuf_0__3157_/X vssd1 vssd1 vccd1 vccd1 _6360__44/A sky130_fd_sc_hd__clkbuf_4
XFILLER_41_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5833__519 _5833__519/A vssd1 vssd1 vccd1 vccd1 _6825_/CLK sky130_fd_sc_hd__inv_2
XFILLER_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3930_ _6781_/Q _3892_/X _3932_/S vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _3861_/A vssd1 vssd1 vccd1 vccd1 _6807_/D sky130_fd_sc_hd__clkbuf_1
X_3792_ _3807_/S vssd1 vssd1 vccd1 vccd1 _3801_/S sky130_fd_sc_hd__buf_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6580_ _6888_/CLK _6580_/D vssd1 vssd1 vccd1 vccd1 _6580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5393_ _5391_/X _5392_/X _5429_/S vssd1 vssd1 vccd1 vccd1 _5393_/X sky130_fd_sc_hd__mux2_1
X_4413_ _4413_/A vssd1 vssd1 vccd1 vccd1 _6586_/D sky130_fd_sc_hd__clkbuf_1
X_7132_ _7132_/A vssd1 vssd1 vccd1 vccd1 _7132_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_113_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4344_ _3782_/X _6616_/Q _4348_/S vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7063_ _7063_/CLK _7063_/D vssd1 vssd1 vccd1 vccd1 _7063_/Q sky130_fd_sc_hd__dfxtp_1
X_6014_ _6885_/Q _6011_/X _6012_/Y _6013_/X vssd1 vssd1 vccd1 vccd1 _6885_/D sky130_fd_sc_hd__o211a_1
X_4275_ _6646_/Q _4164_/X _4275_/S vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3226_ _3226_/A _3623_/B _4068_/C vssd1 vssd1 vccd1 vccd1 _3226_/X sky130_fd_sc_hd__or3_1
XFILLER_100_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6916_ _6916_/CLK _6916_/D vssd1 vssd1 vccd1 vccd1 _6916_/Q sky130_fd_sc_hd__dfxtp_1
X_6847_ _6847_/CLK _6847_/D vssd1 vssd1 vccd1 vccd1 _6847_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3011_ clkbuf_0__3011_/X vssd1 vssd1 vccd1 vccd1 _6102__144/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _7019_/CLK
+ sky130_fd_sc_hd__clkbuf_4
X_6778_ _7011_/CLK _6778_/D vssd1 vssd1 vccd1 vccd1 _6778_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5729_ _5729_/A vssd1 vssd1 vccd1 vccd1 _6745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0__2726_ clkbuf_0__2726_/X vssd1 vssd1 vccd1 vccd1 _5453__298/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5789__484 _5789__484/A vssd1 vssd1 vccd1 vccd1 _6790_/CLK sky130_fd_sc_hd__inv_2
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4060_ _5437_/A vssd1 vssd1 vccd1 vccd1 _4071_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_1_1_0__2861_ clkbuf_0__2861_/X vssd1 vssd1 vccd1 vccd1 _5809_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962_ _7089_/Q vssd1 vssd1 vccd1 vccd1 _6167_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4893_ _6975_/Q _3986_/X _4891_/X _4892_/X vssd1 vssd1 vccd1 vccd1 _4893_/X sky130_fd_sc_hd__o211a_1
X_6701_ _6701_/CLK _6701_/D vssd1 vssd1 vccd1 vccd1 _6701_/Q sky130_fd_sc_hd__dfxtp_1
X_3913_ _3913_/A vssd1 vssd1 vccd1 vccd1 _6789_/D sky130_fd_sc_hd__clkbuf_1
X_6632_ _6632_/CLK _6632_/D vssd1 vssd1 vccd1 vccd1 _6632_/Q sky130_fd_sc_hd__dfxtp_1
X_3844_ _3844_/A vssd1 vssd1 vccd1 vccd1 _6812_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__2518_ clkbuf_0__2518_/X vssd1 vssd1 vccd1 vccd1 _5168__229/A sky130_fd_sc_hd__clkbuf_16
X_6563_ _6563_/CLK _6563_/D vssd1 vssd1 vccd1 vccd1 _6563_/Q sky130_fd_sc_hd__dfxtp_1
X_3775_ _3775_/A vssd1 vssd1 vccd1 vccd1 _6841_/D sky130_fd_sc_hd__clkbuf_1
X_6494_ _6494_/CLK _6494_/D vssd1 vssd1 vccd1 vccd1 _6494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5445_ _6581_/Q _5321_/X _5444_/X _5406_/X vssd1 vssd1 vccd1 vccd1 _6581_/D sky130_fd_sc_hd__o211a_1
XFILLER_105_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7115_ _7115_/A vssd1 vssd1 vccd1 vccd1 _7115_/X sky130_fd_sc_hd__clkbuf_1
X_5376_ _6792_/Q _6982_/Q _6990_/Q _6966_/Q _5264_/A _5276_/X vssd1 vssd1 vccd1 vccd1
+ _5376_/X sky130_fd_sc_hd__mux4_1
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4327_ _4327_/A vssd1 vssd1 vccd1 vccd1 _6624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6118__156 _6119__157/A vssd1 vssd1 vccd1 vccd1 _6964_/CLK sky130_fd_sc_hd__inv_2
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__2511_ clkbuf_0__2511_/X vssd1 vssd1 vccd1 vccd1 _5131__199/A sky130_fd_sc_hd__clkbuf_4
X_7046_ _7046_/CLK _7046_/D vssd1 vssd1 vccd1 vccd1 _7046_/Q sky130_fd_sc_hd__dfxtp_1
X_4258_ _4258_/A vssd1 vssd1 vccd1 vccd1 _6654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3209_ _3273_/B _6730_/Q vssd1 vssd1 vccd1 vccd1 _4068_/A sky130_fd_sc_hd__and2_1
XFILLER_103_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4189_ _4189_/A vssd1 vssd1 vccd1 vccd1 _6685_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5717__445 _5718__446/A vssd1 vssd1 vccd1 vccd1 _6739_/CLK sky130_fd_sc_hd__inv_2
XFILLER_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3560_ _3560_/A vssd1 vssd1 vccd1 vccd1 _6946_/D sky130_fd_sc_hd__clkbuf_1
X_3491_ _3329_/X _6976_/Q _3497_/S vssd1 vssd1 vccd1 vccd1 _3492_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5804__495 _5808__499/A vssd1 vssd1 vccd1 vccd1 _6801_/CLK sky130_fd_sc_hd__inv_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4112_ _4112_/A vssd1 vssd1 vccd1 vccd1 _6719_/D sky130_fd_sc_hd__clkbuf_1
X_5092_ _5092_/A vssd1 vssd1 vccd1 vccd1 _6462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4043_ _4040_/A _4049_/B _4042_/X _4037_/X vssd1 vssd1 vccd1 vccd1 _6738_/D sky130_fd_sc_hd__o211a_1
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5994_ _6881_/Q _5994_/B _5994_/C vssd1 vssd1 vccd1 vccd1 _6004_/C sky130_fd_sc_hd__and3_1
X_4945_ _6859_/Q _6835_/Q _6811_/Q _6803_/Q _4923_/X _4892_/X vssd1 vssd1 vccd1 vccd1
+ _4945_/X sky130_fd_sc_hd__mux4_2
XFILLER_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _4876_/A _6498_/Q vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__or2_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__2743_ _5536_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2743_/X sky130_fd_sc_hd__clkbuf_16
X_6615_ _6615_/CLK _6615_/D vssd1 vssd1 vccd1 vccd1 _6615_/Q sky130_fd_sc_hd__dfxtp_1
X_3827_ _3827_/A _4386_/B vssd1 vssd1 vccd1 vccd1 _3843_/S sky130_fd_sc_hd__nor2_2
XFILLER_118_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6546_ _6546_/CLK _6546_/D vssd1 vssd1 vccd1 vccd1 _6546_/Q sky130_fd_sc_hd__dfxtp_1
X_3758_ _6846_/Q _3614_/X _3762_/S vssd1 vssd1 vccd1 vccd1 _3759_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3689_ _3689_/A vssd1 vssd1 vccd1 vccd1 _6895_/D sky130_fd_sc_hd__clkbuf_1
X_6477_ _6477_/CLK _6477_/D vssd1 vssd1 vccd1 vccd1 _6477_/Q sky130_fd_sc_hd__dfxtp_1
X_5428_ _6677_/Q _6669_/Q _6661_/Q _6653_/Q _5263_/X _5264_/X vssd1 vssd1 vccd1 vccd1
+ _5428_/X sky130_fd_sc_hd__mux4_2
XFILLER_102_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5359_ _7074_/Q _6700_/Q _6569_/Q _6847_/Q _5311_/X _5312_/X vssd1 vssd1 vccd1 vccd1
+ _5359_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XINSDIODE2_2 _3856_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0__3157_ _6355_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3157_/X sky130_fd_sc_hd__clkbuf_16
X_6090__134 _6090__134/A vssd1 vssd1 vccd1 vccd1 _6942_/CLK sky130_fd_sc_hd__inv_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7029_ _7030_/CLK _7029_/D vssd1 vssd1 vccd1 vccd1 _7029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5496__333 _5497__334/A vssd1 vssd1 vccd1 vccd1 _6623_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4923_/A vssd1 vssd1 vccd1 vccd1 _4956_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_119_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4661_ _4661_/A vssd1 vssd1 vccd1 vccd1 _6470_/D sky130_fd_sc_hd__clkbuf_1
X_6400_ _6400_/A vssd1 vssd1 vccd1 vccd1 _7085_/D sky130_fd_sc_hd__clkbuf_1
X_3612_ _6925_/Q _3611_/X _3612_/S vssd1 vssd1 vccd1 vccd1 _3613_/A sky130_fd_sc_hd__mux2_1
X_4592_ _6501_/Q _4009_/A _4600_/S vssd1 vssd1 vccd1 vccd1 _4593_/A sky130_fd_sc_hd__mux2_1
X_3543_ _4205_/A _4386_/B vssd1 vssd1 vccd1 vccd1 _3559_/S sky130_fd_sc_hd__nor2_2
XFILLER_88_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6262_ _6262_/A _6262_/B vssd1 vssd1 vccd1 vccd1 _6263_/C sky130_fd_sc_hd__nand2_1
X_3474_ _3376_/X _6982_/Q _3476_/S vssd1 vssd1 vccd1 vccd1 _3475_/A sky130_fd_sc_hd__mux2_1
X_5213_ _5213_/A vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__buf_1
X_6193_ _6245_/A _6188_/C _6190_/Y _6192_/X vssd1 vssd1 vccd1 vccd1 _6995_/D sky130_fd_sc_hd__o211a_1
X_5144_ _5175_/A vssd1 vssd1 vccd1 vccd1 _5144_/X sky130_fd_sc_hd__buf_1
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__3011_ _6097_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3011_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _5075_/A vssd1 vssd1 vccd1 vccd1 _6454_/D sky130_fd_sc_hd__clkbuf_1
X_4026_ _4026_/A vssd1 vssd1 vccd1 vccd1 _4026_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2758_ clkbuf_0__2758_/X vssd1 vssd1 vccd1 vccd1 _5678__414/A sky130_fd_sc_hd__clkbuf_4
X_5977_ _6013_/A vssd1 vssd1 vccd1 vccd1 _6002_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4928_ _6765_/Q _6757_/Q _6720_/Q _6712_/Q _4923_/X _4892_/X vssd1 vssd1 vccd1 vccd1
+ _4928_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_0__2726_ _5449_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2726_/X sky130_fd_sc_hd__clkbuf_16
X_4859_ _7093_/Q vssd1 vssd1 vccd1 vccd1 _6173_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6529_ _6529_/CLK _6529_/D vssd1 vssd1 vccd1 vccd1 _6529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5900_ _5888_/C _5610_/X _6012_/D vssd1 vssd1 vccd1 vccd1 _5900_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6880_ _7008_/CLK _6880_/D vssd1 vssd1 vccd1 vccd1 _6880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5173__233 _5174__234/A vssd1 vssd1 vccd1 vccd1 _6515_/CLK sky130_fd_sc_hd__inv_2
X_4713_ _4868_/S vssd1 vssd1 vccd1 vccd1 _4876_/A sky130_fd_sc_hd__buf_2
Xclkbuf_0__2511_ _5126_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2511_/X sky130_fd_sc_hd__clkbuf_16
X_4644_ _4644_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4660_/S sky130_fd_sc_hd__or2_2
X_4575_ _4575_/A vssd1 vssd1 vccd1 vccd1 _6509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6314_ _7130_/A _6314_/B _6318_/C vssd1 vssd1 vccd1 vccd1 _6315_/A sky130_fd_sc_hd__and3_1
X_3526_ _6961_/Q _3437_/X _3534_/S vssd1 vssd1 vccd1 vccd1 _3527_/A sky130_fd_sc_hd__mux2_1
X_6245_ _6245_/A _6245_/B vssd1 vssd1 vccd1 vccd1 _6245_/Y sky130_fd_sc_hd__nor2_1
X_5696__429 _5696__429/A vssd1 vssd1 vccd1 vccd1 _6723_/CLK sky130_fd_sc_hd__inv_2
X_3457_ _6988_/Q _3456_/X _3463_/S vssd1 vssd1 vccd1 vccd1 _3458_/A sky130_fd_sc_hd__mux2_1
X_6176_ _7002_/Q vssd1 vssd1 vccd1 vccd1 _6241_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3388_ _3785_/A vssd1 vssd1 vccd1 vccd1 _3388_/X sky130_fd_sc_hd__buf_2
X_5058_ _5058_/A vssd1 vssd1 vccd1 vccd1 _6447_/D sky130_fd_sc_hd__clkbuf_1
X_5592__405 _5594__407/A vssd1 vssd1 vccd1 vccd1 _6698_/CLK sky130_fd_sc_hd__inv_2
X_4009_ _4009_/A vssd1 vssd1 vccd1 vccd1 _4009_/X sky130_fd_sc_hd__buf_4
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5783__479 _5783__479/A vssd1 vssd1 vccd1 vccd1 _6785_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4360_ _6609_/Q _3779_/A _4360_/S vssd1 vssd1 vccd1 vccd1 _4361_/A sky130_fd_sc_hd__mux2_1
X_3311_ _3308_/X _3309_/X _3960_/A vssd1 vssd1 vccd1 vccd1 _3318_/B sky130_fd_sc_hd__mux2_1
X_6332__21 _6335__24/A vssd1 vssd1 vccd1 vccd1 _7041_/CLK sky130_fd_sc_hd__inv_2
XFILLER_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _4291_/A vssd1 vssd1 vccd1 vccd1 _6640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3242_ _3242_/A vssd1 vssd1 vccd1 vccd1 _3242_/X sky130_fd_sc_hd__buf_4
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5244__289 _5244__289/A vssd1 vssd1 vccd1 vccd1 _6571_/CLK sky130_fd_sc_hd__inv_2
XFILLER_82_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6932_ _6932_/CLK _6932_/D vssd1 vssd1 vccd1 vccd1 _6932_/Q sky130_fd_sc_hd__dfxtp_1
X_6863_ _6863_/CLK _6863_/D vssd1 vssd1 vccd1 vccd1 _6863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0__2526_ clkbuf_0__2526_/X vssd1 vssd1 vccd1 vccd1 _5213_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6794_ _6794_/CLK _6794_/D vssd1 vssd1 vccd1 vccd1 _6794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2457_ clkbuf_0__2457_/X vssd1 vssd1 vccd1 vccd1 _5037_/A sky130_fd_sc_hd__clkbuf_4
X_4627_ _4642_/S vssd1 vssd1 vccd1 vccd1 _4636_/S sky130_fd_sc_hd__buf_2
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4558_ _6516_/Q _4014_/A _4562_/S vssd1 vssd1 vccd1 vccd1 _4559_/A sky130_fd_sc_hd__mux2_1
X_4489_ _4489_/A vssd1 vssd1 vccd1 vccd1 _6546_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3509_ _3509_/A vssd1 vssd1 vccd1 vccd1 _6969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__2742_ clkbuf_0__2742_/X vssd1 vssd1 vccd1 vccd1 _5535__364/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6228_ _6241_/C _6228_/B vssd1 vssd1 vccd1 vccd1 _6229_/B sky130_fd_sc_hd__or2_1
Xclkbuf_1_1_0__3009_ clkbuf_0__3009_/X vssd1 vssd1 vccd1 vccd1 _6088__132/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6159_ _6155_/A _6262_/A _6168_/B _6168_/A vssd1 vssd1 vccd1 vccd1 _6159_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_0__3156_ clkbuf_0__3156_/X vssd1 vssd1 vccd1 vccd1 _6352__37/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6111__151 _6113__153/A vssd1 vssd1 vccd1 vccd1 _6959_/CLK sky130_fd_sc_hd__inv_2
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _6807_/Q _3859_/X _3860_/S vssd1 vssd1 vccd1 vccd1 _3861_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3791_ _4458_/A _3873_/B vssd1 vssd1 vccd1 vccd1 _3807_/S sky130_fd_sc_hd__or2_2
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5530_ _5554_/A vssd1 vssd1 vccd1 vccd1 _5530_/X sky130_fd_sc_hd__buf_1
XFILLER_118_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5461_ _5461_/A vssd1 vssd1 vccd1 vccd1 _5461_/X sky130_fd_sc_hd__buf_1
X_4412_ _3257_/X _6586_/Q _4414_/S vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__mux2_1
X_5392_ _6603_/Q _6587_/Q _6841_/Q _6825_/Q _5329_/X _5330_/X vssd1 vssd1 vccd1 vccd1
+ _5392_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_7131_ _7131_/A vssd1 vssd1 vccd1 vccd1 _7131_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4343_ _4343_/A vssd1 vssd1 vccd1 vccd1 _6617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7062_ _7062_/CLK _7062_/D vssd1 vssd1 vccd1 vccd1 _7062_/Q sky130_fd_sc_hd__dfxtp_1
X_4274_ _4274_/A vssd1 vssd1 vccd1 vccd1 _6647_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6013_ _6013_/A _6013_/B vssd1 vssd1 vccd1 vccd1 _6013_/X sky130_fd_sc_hd__and2_2
X_3225_ _4277_/C _3221_/A _3226_/A _4068_/B _3224_/X vssd1 vssd1 vccd1 vccd1 _3227_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_94_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6915_ _6915_/CLK _6915_/D vssd1 vssd1 vccd1 vccd1 _6915_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__3010_ clkbuf_0__3010_/X vssd1 vssd1 vccd1 vccd1 _6094__137/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6846_ _6846_/CLK _6846_/D vssd1 vssd1 vccd1 vccd1 _6846_/Q sky130_fd_sc_hd__dfxtp_1
X_6777_ _6777_/CLK _6777_/D vssd1 vssd1 vccd1 vccd1 _6777_/Q sky130_fd_sc_hd__dfxtp_1
X_5728_ _7019_/Q _5734_/B vssd1 vssd1 vccd1 vccd1 _5729_/A sky130_fd_sc_hd__and2_1
X_3989_ _3989_/A vssd1 vssd1 vccd1 vccd1 _6767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5659_ _7083_/Q _5659_/B vssd1 vssd1 vccd1 vccd1 _5897_/B sky130_fd_sc_hd__xor2_2
X_5186__243 _5186__243/A vssd1 vssd1 vccd1 vccd1 _6525_/CLK sky130_fd_sc_hd__inv_2
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5490__328 _5491__329/A vssd1 vssd1 vccd1 vccd1 _6618_/CLK sky130_fd_sc_hd__inv_2
XFILLER_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__3154_ clkbuf_0__3154_/X vssd1 vssd1 vccd1 vccd1 _6355_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5796__489 _5796__489/A vssd1 vssd1 vccd1 vccd1 _6795_/CLK sky130_fd_sc_hd__inv_2
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0__2860_ clkbuf_0__2860_/X vssd1 vssd1 vccd1 vccd1 _5786__481/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4961_ _4726_/X _4954_/X _4960_/X _3971_/X vssd1 vssd1 vccd1 vccd1 _4961_/X sky130_fd_sc_hd__a211o_1
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4892_ _4914_/A vssd1 vssd1 vccd1 vccd1 _4892_/X sky130_fd_sc_hd__clkbuf_4
X_6700_ _6700_/CLK _6700_/D vssd1 vssd1 vccd1 vccd1 _6700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3912_ _6789_/Q _3617_/X _3914_/S vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__mux2_1
X_3843_ _6812_/Q _3620_/X _3843_/S vssd1 vssd1 vccd1 vccd1 _3844_/A sky130_fd_sc_hd__mux2_1
X_6631_ _6631_/CLK _6631_/D vssd1 vssd1 vccd1 vccd1 _6631_/Q sky130_fd_sc_hd__dfxtp_1
X_6562_ _6562_/CLK _6562_/D vssd1 vssd1 vccd1 vccd1 _6562_/Q sky130_fd_sc_hd__dfxtp_1
X_3774_ _3773_/X _6841_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3775_/A sky130_fd_sc_hd__mux2_1
X_6493_ _6493_/CLK _6493_/D vssd1 vssd1 vccd1 vccd1 _6493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5444_ _5324_/X _5433_/X _5443_/Y vssd1 vssd1 vccd1 vccd1 _5444_/X sky130_fd_sc_hd__a21o_1
X_7114_ _7114_/A vssd1 vssd1 vccd1 vccd1 _7114_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_99_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5375_ _5371_/X _5374_/X _5394_/S vssd1 vssd1 vccd1 vccd1 _5375_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4326_ _6624_/Q _3889_/X _4330_/S vssd1 vssd1 vccd1 vccd1 _4327_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0__2510_ clkbuf_0__2510_/X vssd1 vssd1 vccd1 vccd1 _5123__192/A sky130_fd_sc_hd__clkbuf_4
X_7045_ _7045_/CLK _7045_/D vssd1 vssd1 vccd1 vccd1 _7045_/Q sky130_fd_sc_hd__dfxtp_1
X_4257_ _3788_/X _6654_/Q _4257_/S vssd1 vssd1 vccd1 vccd1 _4258_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4188_ _6685_/Q _4141_/X _4196_/S vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3208_ _6735_/Q vssd1 vssd1 vccd1 vccd1 _3273_/B sky130_fd_sc_hd__inv_2
XFILLER_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6829_ _6829_/CLK _6829_/D vssd1 vssd1 vccd1 vccd1 _6829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6366__49 _6366__49/A vssd1 vssd1 vccd1 vccd1 _7069_/CLK sky130_fd_sc_hd__inv_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3490_ _3490_/A vssd1 vssd1 vccd1 vccd1 _6977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4111_ _6719_/Q _3880_/X _4115_/S vssd1 vssd1 vccd1 vccd1 _4112_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5091_ _6462_/Q _7116_/A _5093_/S vssd1 vssd1 vccd1 vccd1 _5092_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4042_ _4044_/A _4044_/B _4277_/B vssd1 vssd1 vccd1 vccd1 _4042_/X sky130_fd_sc_hd__a21o_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _5993_/A vssd1 vssd1 vccd1 vccd1 _6880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4944_ _4944_/A _4944_/B vssd1 vssd1 vccd1 vccd1 _4944_/X sky130_fd_sc_hd__or2_1
X_5137__204 _5137__204/A vssd1 vssd1 vccd1 vccd1 _6486_/CLK sky130_fd_sc_hd__inv_2
X_4875_ _4873_/X _4874_/X _4875_/S vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2742_ _5530_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2742_/X sky130_fd_sc_hd__clkbuf_16
X_6124__161 _6124__161/A vssd1 vssd1 vccd1 vccd1 _6969_/CLK sky130_fd_sc_hd__inv_2
X_6614_ _6614_/CLK _6614_/D vssd1 vssd1 vccd1 vccd1 _6614_/Q sky130_fd_sc_hd__dfxtp_1
X_3826_ _3826_/A vssd1 vssd1 vccd1 vccd1 _6820_/D sky130_fd_sc_hd__clkbuf_1
X_6545_ _6545_/CLK _6545_/D vssd1 vssd1 vccd1 vccd1 _6545_/Q sky130_fd_sc_hd__dfxtp_1
X_3757_ _3757_/A vssd1 vssd1 vccd1 vccd1 _6847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3688_ _3687_/X _6895_/Q _3697_/S vssd1 vssd1 vccd1 vccd1 _3689_/A sky130_fd_sc_hd__mux2_1
X_6476_ _6476_/CLK _6476_/D vssd1 vssd1 vccd1 vccd1 _6476_/Q sky130_fd_sc_hd__dfxtp_1
X_5427_ _7078_/Q _6704_/Q _6573_/Q _6851_/Q _5257_/X _5259_/X vssd1 vssd1 vccd1 vccd1
+ _5427_/X sky130_fd_sc_hd__mux4_1
X_5358_ _4071_/A _5351_/X _5353_/Y _5355_/X _5357_/Y vssd1 vssd1 vccd1 vccd1 _5358_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XINSDIODE2_3 _3877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__3156_ _6349_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3156_/X sky130_fd_sc_hd__clkbuf_16
X_4309_ _4309_/A vssd1 vssd1 vccd1 vccd1 _6632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7028_ _7030_/CLK _7028_/D vssd1 vssd1 vccd1 vccd1 _7028_/Q sky130_fd_sc_hd__dfxtp_1
X_5289_ _5435_/B vssd1 vssd1 vccd1 vccd1 _5289_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5859__59 _5859__59/A vssd1 vssd1 vccd1 vccd1 _6845_/CLK sky130_fd_sc_hd__inv_2
XFILLER_3_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6067__115 _6069__117/A vssd1 vssd1 vccd1 vccd1 _6923_/CLK sky130_fd_sc_hd__inv_2
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6339__27 _6341__29/A vssd1 vssd1 vccd1 vccd1 _7047_/CLK sky130_fd_sc_hd__inv_2
XFILLER_119_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _3868_/X _6470_/Q _4660_/S vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__mux2_1
X_3611_ _7026_/Q vssd1 vssd1 vccd1 vccd1 _3611_/X sky130_fd_sc_hd__buf_4
X_4591_ _4606_/S vssd1 vssd1 vccd1 vccd1 _4600_/S sky130_fd_sc_hd__clkbuf_2
X_6330_ _6330_/A vssd1 vssd1 vccd1 vccd1 _6330_/X sky130_fd_sc_hd__buf_1
X_3542_ _4277_/A _4277_/B _4044_/A vssd1 vssd1 vccd1 vccd1 _4386_/B sky130_fd_sc_hd__or3_4
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6261_ _6262_/A _6262_/B vssd1 vssd1 vccd1 vccd1 _6266_/B sky130_fd_sc_hd__nor2_1
X_3473_ _3473_/A vssd1 vssd1 vccd1 vccd1 _6983_/D sky130_fd_sc_hd__clkbuf_1
X_6192_ _6247_/A vssd1 vssd1 vccd1 vccd1 _6192_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_0__3010_ _6091_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__3010_/X sky130_fd_sc_hd__clkbuf_16
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5074_ _6454_/Q _7108_/A _5082_/S vssd1 vssd1 vccd1 vccd1 _5075_/A sky130_fd_sc_hd__mux2_1
X_4025_ _4025_/A vssd1 vssd1 vccd1 vccd1 _6754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5976_ _5976_/A _5976_/B vssd1 vssd1 vccd1 vccd1 _6877_/D sky130_fd_sc_hd__nor2_1
X_4927_ _4927_/A _4927_/B vssd1 vssd1 vccd1 vccd1 _4927_/X sky130_fd_sc_hd__or2_1
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4858_ _4844_/X _4855_/X _4856_/Y _4857_/Y _5739_/C vssd1 vssd1 vccd1 vccd1 _4858_/X
+ sky130_fd_sc_hd__a32o_1
X_3809_ _3827_/A _4404_/B vssd1 vssd1 vccd1 vccd1 _3825_/S sky130_fd_sc_hd__nor2_2
XFILLER_119_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4789_ _6471_/Q _6623_/Q _7056_/Q _6781_/Q _4709_/X _4772_/S vssd1 vssd1 vccd1 vccd1
+ _4790_/B sky130_fd_sc_hd__mux4_1
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6528_ _6528_/CLK _6528_/D vssd1 vssd1 vccd1 vccd1 _6528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6459_ _7089_/CLK _6459_/D vssd1 vssd1 vccd1 vccd1 _6459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6344__30 _6348__34/A vssd1 vssd1 vccd1 vccd1 _7050_/CLK sky130_fd_sc_hd__inv_2
XFILLER_112_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4712_ _4716_/A _4710_/X _4711_/X vssd1 vssd1 vccd1 vccd1 _4712_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_0__2510_ _5120_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__2510_/X sky130_fd_sc_hd__clkbuf_16
X_4643_ _4643_/A vssd1 vssd1 vccd1 vccd1 _6478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4574_ _4476_/X _6509_/Q _4582_/S vssd1 vssd1 vccd1 vccd1 _4575_/A sky130_fd_sc_hd__mux2_1
X_6313_ _6313_/A vssd1 vssd1 vccd1 vccd1 _7027_/D sky130_fd_sc_hd__clkbuf_1
X_3525_ _3540_/S vssd1 vssd1 vccd1 vccd1 _3534_/S sky130_fd_sc_hd__buf_2
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _6250_/A _6249_/D vssd1 vssd1 vccd1 vccd1 _6244_/Y sky130_fd_sc_hd__nand2_1
X_3456_ _3782_/A vssd1 vssd1 vccd1 vccd1 _3456_/X sky130_fd_sc_hd__buf_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6175_ _6175_/A _6175_/B _5652_/C vssd1 vssd1 vccd1 vccd1 _6175_/X sky130_fd_sc_hd__or3b_1
X_3387_ _7024_/Q vssd1 vssd1 vccd1 vccd1 _3785_/A sky130_fd_sc_hd__clkbuf_4
X_5180__238 _5181__239/A vssd1 vssd1 vccd1 vccd1 _6520_/CLK sky130_fd_sc_hd__inv_2
X_5126_ _5138_/A vssd1 vssd1 vccd1 vccd1 _5126_/X sky130_fd_sc_hd__buf_1
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5057_ _6447_/Q _7101_/A _5116_/B vssd1 vssd1 vccd1 vccd1 _5058_/A sky130_fd_sc_hd__mux2_1
X_4008_ _4008_/A vssd1 vssd1 vccd1 vccd1 _6759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5959_ _5976_/A _5959_/B vssd1 vssd1 vccd1 vccd1 _6874_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3310_ _6773_/Q _6768_/Q vssd1 vssd1 vccd1 vccd1 _3960_/A sky130_fd_sc_hd__xor2_1
XFILLER_6_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ _6640_/Q _4158_/X _4294_/S vssd1 vssd1 vccd1 vccd1 _4291_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3241_ _6694_/Q _5044_/A _3241_/C _5044_/B vssd1 vssd1 vccd1 vccd1 _3242_/A sky130_fd_sc_hd__and4_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6931_ _6931_/CLK _6931_/D vssd1 vssd1 vccd1 vccd1 _6931_/Q sky130_fd_sc_hd__dfxtp_1
X_6862_ _6862_/CLK _6862_/D vssd1 vssd1 vccd1 vccd1 _6862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0__2525_ clkbuf_0__2525_/X vssd1 vssd1 vccd1 vccd1 _5202__256/A sky130_fd_sc_hd__clkbuf_4
X_6793_ _6793_/CLK _6793_/D vssd1 vssd1 vccd1 vccd1 _6793_/Q sky130_fd_sc_hd__dfxtp_1
X_5744_ _5750_/A vssd1 vssd1 vccd1 vccd1 _5744_/X sky130_fd_sc_hd__buf_1
Xclkbuf_1_1_0__2456_ clkbuf_0__2456_/X vssd1 vssd1 vccd1 vccd1 _5035__184/A sky130_fd_sc_hd__clkbuf_4
X_5675_ _5675_/A vssd1 vssd1 vccd1 vccd1 _6705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4626_ _4626_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4642_/S sky130_fd_sc_hd__or2_2
XFILLER_116_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4557_ _4557_/A vssd1 vssd1 vccd1 vccd1 _6517_/D sky130_fd_sc_hd__clkbuf_1
X_4488_ _4487_/X _6546_/Q _4491_/S vssd1 vssd1 vccd1 vccd1 _4489_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3508_ _6969_/Q _3437_/X _3516_/S vssd1 vssd1 vccd1 vccd1 _3509_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0__2741_ clkbuf_0__2741_/X vssd1 vssd1 vccd1 vccd1 _5548_/A sky130_fd_sc_hd__clkbuf_4
X_6227_ _6241_/C _6228_/B vssd1 vssd1 vccd1 vccd1 _6237_/C sky130_fd_sc_hd__and2_1
Xclkbuf_1_1_0__3008_ clkbuf_0__3008_/X vssd1 vssd1 vccd1 vccd1 _6097_/A sky130_fd_sc_hd__clkbuf_4
X_3439_ _4277_/A _4277_/B _4277_/C vssd1 vssd1 vccd1 vccd1 _3898_/B sky130_fd_sc_hd__or3_4
XFILLER_106_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_6158_ _7003_/Q vssd1 vssd1 vccd1 vccd1 _6168_/B sky130_fd_sc_hd__inv_2
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _6578_/Q _6579_/Q _6580_/Q _6581_/Q _6886_/Q _6887_/Q vssd1 vssd1 vccd1 vccd1
+ _5109_/X sky130_fd_sc_hd__mux4_1
XFILLER_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0__3155_ clkbuf_0__3155_/X vssd1 vssd1 vccd1 vccd1 _6347__33/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _3790_/A vssd1 vssd1 vccd1 vccd1 _6836_/D sky130_fd_sc_hd__clkbuf_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4411_ _4411_/A vssd1 vssd1 vccd1 vccd1 _6587_/D sky130_fd_sc_hd__clkbuf_1
X_5391_ _6643_/Q _6635_/Q _6619_/Q _6611_/Q _4083_/A _4063_/A vssd1 vssd1 vccd1 vccd1
+ _5391_/X sky130_fd_sc_hd__mux4_1
X_7130_ _7130_/A vssd1 vssd1 vccd1 vccd1 _7130_/X sky130_fd_sc_hd__clkbuf_1
X_4342_ _3779_/X _6617_/Q _4342_/S vssd1 vssd1 vccd1 vccd1 _4343_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7061_ _7061_/CLK _7061_/D vssd1 vssd1 vccd1 vccd1 _7061_/Q sky130_fd_sc_hd__dfxtp_1
X_4273_ _6647_/Q _4161_/X _4275_/S vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6012_ _5954_/B _6012_/B _6885_/Q _6012_/D vssd1 vssd1 vccd1 vccd1 _6012_/Y sky130_fd_sc_hd__nand4b_1
X_3224_ _3273_/B _6730_/Q _3222_/Y _3223_/X vssd1 vssd1 vccd1 vccd1 _3224_/X sky130_fd_sc_hd__o211a_1
.ends

