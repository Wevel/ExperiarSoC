VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Art
  CLASS BLOCK ;
  FOREIGN Art ;
  ORIGIN 0.800 1.000 ;
  SIZE 504.920 BY 501.000 ;
  PIN dumyPin
    PORT
      LAYER met2 ;
        RECT 9.000 -1.000 11.000 1.000 ;
    END
  END dumyPin
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -0.80000 0.00000 0.80000 500.00000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 499.20000 0.00000 500.80000 500.00000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.000 30.000 105.000 70.000 ;
        RECT 5.000 5.000 25.000 25.000 ;
      LAYER met1 ;
        RECT 85.000 60.000 105.000 70.120 ;
        RECT 65.000 50.000 105.000 60.000 ;
        RECT 45.000 40.000 105.000 50.000 ;
        RECT 25.000 30.120 105.000 40.000 ;
        RECT 25.000 30.000 85.000 30.120 ;
        RECT 25.000 5.000 45.000 25.000 ;
      LAYER met2 ;
        RECT 45.000 60.000 65.000 70.000 ;
        RECT 25.000 50.000 45.000 60.000 ;
        RECT 85.000 50.000 105.000 60.000 ;
        RECT 5.000 40.000 25.000 50.000 ;
        RECT 65.000 40.000 105.000 50.000 ;
        RECT 45.000 30.000 105.000 40.000 ;
        RECT 45.000 5.000 65.000 25.000 ;
      LAYER met3 ;
        RECT 25.000 60.000 45.000 70.000 ;
        RECT 5.000 50.000 25.000 60.000 ;
        RECT 85.000 40.000 105.000 50.000 ;
        RECT 65.000 30.000 105.000 40.000 ;
        RECT 65.000 5.000 85.000 25.000 ;
      LAYER met4 ;
        RECT -0.800 0.000 0.800 500.000 ;
        RECT 45.770 486.600 51.770 488.600 ;
        RECT 45.770 484.600 47.770 486.600 ;
        RECT 43.770 482.600 47.770 484.600 ;
        RECT 49.770 484.600 51.770 486.600 ;
        RECT 49.770 482.600 53.770 484.600 ;
        RECT 43.770 478.600 45.770 482.600 ;
        RECT 41.770 476.600 45.770 478.600 ;
        RECT 51.770 478.600 53.770 482.600 ;
        RECT 51.770 476.600 55.770 478.600 ;
        RECT 41.770 472.600 43.770 476.600 ;
        RECT 39.770 470.600 43.770 472.600 ;
        RECT 45.770 470.600 49.770 474.600 ;
        RECT 53.770 472.600 55.770 476.600 ;
        RECT 53.770 470.600 57.770 472.600 ;
        RECT 39.770 466.600 41.770 470.600 ;
        RECT 37.770 464.600 41.770 466.600 ;
        RECT 43.770 468.600 49.770 470.600 ;
        RECT 55.770 468.600 57.770 470.600 ;
        RECT 43.770 466.600 51.770 468.600 ;
        RECT 55.770 466.600 59.770 468.600 ;
        RECT 43.770 464.600 53.770 466.600 ;
        RECT 37.770 462.600 39.770 464.600 ;
        RECT 35.770 460.600 39.770 462.600 ;
        RECT 41.770 460.600 49.770 464.600 ;
        RECT 35.770 456.600 37.770 460.600 ;
        RECT 33.770 454.600 37.770 456.600 ;
        RECT 39.770 456.600 49.770 460.600 ;
        RECT 51.770 460.600 55.770 464.600 ;
        RECT 57.770 462.600 59.770 466.600 ;
        RECT 57.770 460.600 61.770 462.600 ;
        RECT 51.770 456.600 57.770 460.600 ;
        RECT 39.770 454.600 51.770 456.600 ;
        RECT 33.770 452.600 35.770 454.600 ;
        RECT 27.770 450.600 35.770 452.600 ;
        RECT 37.770 450.600 51.770 454.600 ;
        RECT 53.770 454.600 57.770 456.600 ;
        RECT 59.770 456.600 61.770 460.600 ;
        RECT 59.770 454.600 63.770 456.600 ;
        RECT 53.770 452.600 59.770 454.600 ;
        RECT 53.770 450.600 55.770 452.600 ;
        RECT 61.770 450.600 63.770 454.600 ;
        RECT 17.770 448.600 29.770 450.600 ;
        RECT 37.770 448.600 53.770 450.600 ;
        RECT 55.770 448.600 59.770 450.600 ;
        RECT 61.770 448.600 71.770 450.600 ;
        RECT 11.770 446.600 19.770 448.600 ;
        RECT 29.770 446.600 33.770 448.600 ;
        RECT 11.770 442.600 13.770 446.600 ;
        RECT 19.770 444.600 33.770 446.600 ;
        RECT 35.770 444.600 61.770 448.600 ;
        RECT 69.770 446.600 79.770 448.600 ;
        RECT 63.770 444.600 65.770 446.600 ;
        RECT 77.770 444.600 87.770 446.600 ;
        RECT 19.770 442.600 35.770 444.600 ;
        RECT 45.770 442.600 57.770 444.600 ;
        RECT 61.770 442.600 69.770 444.600 ;
        RECT 85.770 442.600 91.770 444.600 ;
        RECT 11.770 440.600 19.770 442.600 ;
        RECT 29.770 440.600 45.770 442.600 ;
        RECT 57.770 440.600 75.770 442.600 ;
        RECT 89.770 440.600 91.770 442.600 ;
        RECT 17.770 438.600 29.770 440.600 ;
        RECT 39.770 438.600 79.770 440.600 ;
        RECT 87.770 438.600 91.770 440.600 ;
        RECT 27.770 436.600 39.770 438.600 ;
        RECT 49.770 436.600 77.770 438.600 ;
        RECT 85.770 436.600 89.770 438.600 ;
        RECT 29.770 434.600 31.770 436.600 ;
        RECT 27.770 432.600 31.770 434.600 ;
        RECT 33.770 434.600 49.770 436.600 ;
        RECT 59.770 434.600 69.770 436.600 ;
        RECT 77.770 434.600 87.770 436.600 ;
        RECT 33.770 432.600 59.770 434.600 ;
        RECT 69.770 432.600 79.770 434.600 ;
        RECT 27.770 426.600 29.770 432.600 ;
        RECT 31.770 430.600 49.770 432.600 ;
        RECT 59.770 430.600 71.770 432.600 ;
        RECT 31.770 428.600 47.770 430.600 ;
        RECT 33.770 426.600 47.770 428.600 ;
        RECT 49.770 428.600 53.770 430.600 ;
        RECT 57.770 428.600 59.770 430.600 ;
        RECT 63.770 428.600 65.770 430.600 ;
        RECT 69.770 428.600 71.770 430.600 ;
        RECT 79.770 428.600 85.770 430.600 ;
        RECT 49.770 426.600 51.770 428.600 ;
        RECT 63.770 426.600 71.770 428.600 ;
        RECT 77.770 426.600 81.770 428.600 ;
        RECT 83.770 426.600 85.770 428.600 ;
        RECT 25.770 424.600 31.770 426.600 ;
        RECT 23.770 422.600 27.770 424.600 ;
        RECT 29.770 422.600 35.770 424.600 ;
        RECT 37.770 422.600 47.770 426.600 ;
        RECT 51.770 424.600 53.770 426.600 ;
        RECT 63.770 424.600 67.770 426.600 ;
        RECT 73.770 424.600 79.770 426.600 ;
        RECT 81.770 424.600 85.770 426.600 ;
        RECT 61.770 422.600 67.770 424.600 ;
        RECT 69.770 422.600 75.770 424.600 ;
        RECT 21.770 420.600 25.770 422.600 ;
        RECT 27.770 420.600 37.770 422.600 ;
        RECT 41.770 420.600 49.770 422.600 ;
        RECT 55.770 420.600 71.770 422.600 ;
        RECT 75.770 420.600 79.770 422.600 ;
        RECT 21.770 414.600 23.770 420.600 ;
        RECT 19.770 412.600 23.770 414.600 ;
        RECT 25.770 418.600 39.770 420.600 ;
        RECT 43.770 418.600 49.770 420.600 ;
        RECT 59.770 418.600 67.770 420.600 ;
        RECT 71.770 418.600 81.770 420.600 ;
        RECT 83.770 418.600 85.770 424.600 ;
        RECT 25.770 416.600 43.770 418.600 ;
        RECT 45.770 416.600 49.770 418.600 ;
        RECT 57.770 416.600 63.770 418.600 ;
        RECT 67.770 416.600 77.770 418.600 ;
        RECT 81.770 416.600 85.770 418.600 ;
        RECT 25.770 414.600 45.770 416.600 ;
        RECT 53.770 414.600 59.770 416.600 ;
        RECT 63.770 414.600 75.770 416.600 ;
        RECT 25.770 412.600 65.770 414.600 ;
        RECT 73.770 412.600 75.770 414.600 ;
        RECT 77.770 414.600 83.770 416.600 ;
        RECT 77.770 412.600 79.770 414.600 ;
        RECT 19.770 392.600 21.770 412.600 ;
        RECT 23.770 410.600 39.770 412.600 ;
        RECT 41.770 410.600 43.770 412.600 ;
        RECT 47.770 410.600 59.770 412.600 ;
        RECT 23.770 408.600 37.770 410.600 ;
        RECT 39.770 408.600 41.770 410.600 ;
        RECT 43.770 408.600 47.770 410.600 ;
        RECT 53.770 408.600 57.770 410.600 ;
        RECT 59.770 408.600 61.770 410.600 ;
        RECT 75.770 408.600 79.770 412.600 ;
        RECT 23.770 406.600 39.770 408.600 ;
        RECT 41.770 406.600 43.770 408.600 ;
        RECT 23.770 404.600 37.770 406.600 ;
        RECT 39.770 404.600 43.770 406.600 ;
        RECT 47.770 406.600 57.770 408.600 ;
        RECT 61.770 406.600 79.770 408.600 ;
        RECT 47.770 404.600 49.770 406.600 ;
        RECT 55.770 404.600 59.770 406.600 ;
        RECT 63.770 404.600 65.770 406.600 ;
        RECT 77.770 404.600 81.770 406.600 ;
        RECT 23.770 402.600 39.770 404.600 ;
        RECT 41.770 402.600 43.770 404.600 ;
        RECT 49.770 402.600 53.770 404.600 ;
        RECT 23.770 400.600 41.770 402.600 ;
        RECT 43.770 400.600 45.770 402.600 ;
        RECT 51.770 400.600 53.770 402.600 ;
        RECT 55.770 402.600 57.770 404.600 ;
        RECT 55.770 400.600 59.770 402.600 ;
        RECT 61.770 400.600 63.770 404.600 ;
        RECT 79.770 402.600 83.770 404.600 ;
        RECT 75.770 400.600 79.770 402.600 ;
        RECT 23.770 398.600 39.770 400.600 ;
        RECT 45.770 398.600 47.770 400.600 ;
        RECT 53.770 398.600 61.770 400.600 ;
        RECT 63.770 398.600 67.770 400.600 ;
        RECT 71.770 398.600 77.770 400.600 ;
        RECT 81.770 398.600 83.770 402.600 ;
        RECT 23.770 396.600 41.770 398.600 ;
        RECT 47.770 396.600 49.770 398.600 ;
        RECT 57.770 396.600 63.770 398.600 ;
        RECT 67.770 396.600 71.770 398.600 ;
        RECT 77.770 396.600 83.770 398.600 ;
        RECT 23.770 394.600 39.770 396.600 ;
        RECT 49.770 394.600 51.770 396.600 ;
        RECT 59.770 394.600 67.770 396.600 ;
        RECT 71.770 394.600 79.770 396.600 ;
        RECT 23.770 392.600 37.770 394.600 ;
        RECT 39.770 392.600 41.770 394.600 ;
        RECT 51.770 392.600 55.770 394.600 ;
        RECT 65.770 392.600 73.770 394.600 ;
        RECT 19.770 390.600 23.770 392.600 ;
        RECT 21.770 374.600 23.770 390.600 ;
        RECT 25.770 388.600 35.770 392.600 ;
        RECT 37.770 390.600 39.770 392.600 ;
        RECT 41.770 390.600 43.770 392.600 ;
        RECT 55.770 390.600 69.770 392.600 ;
        RECT 39.770 388.600 41.770 390.600 ;
        RECT 55.770 388.600 65.770 390.600 ;
        RECT 25.770 386.600 39.770 388.600 ;
        RECT 41.770 386.600 43.770 388.600 ;
        RECT 57.770 386.600 65.770 388.600 ;
        RECT 25.770 384.600 37.770 386.600 ;
        RECT 39.770 384.600 41.770 386.600 ;
        RECT 25.770 382.600 39.770 384.600 ;
        RECT 41.770 382.600 43.770 384.600 ;
        RECT 57.770 382.600 67.770 386.600 ;
        RECT 25.770 380.600 41.770 382.600 ;
        RECT 25.770 378.600 39.770 380.600 ;
        RECT 41.770 378.600 43.770 380.600 ;
        RECT 59.770 378.600 67.770 382.600 ;
        RECT 25.770 376.600 41.770 378.600 ;
        RECT 25.770 374.600 39.770 376.600 ;
        RECT 41.770 374.600 43.770 376.600 ;
        RECT 61.770 374.600 67.770 378.600 ;
        RECT 21.770 372.600 25.770 374.600 ;
        RECT 27.770 372.600 41.770 374.600 ;
        RECT 59.770 372.600 61.770 374.600 ;
        RECT 65.770 372.600 67.770 374.600 ;
        RECT 23.770 370.600 25.770 372.600 ;
        RECT 31.770 370.600 39.770 372.600 ;
        RECT 41.770 370.600 43.770 372.600 ;
        RECT 45.770 370.600 47.770 372.600 ;
        RECT 49.770 370.600 51.770 372.600 ;
        RECT 53.770 370.600 55.770 372.600 ;
        RECT 57.770 370.600 59.770 372.600 ;
        RECT 61.770 370.600 67.770 372.600 ;
        RECT 23.770 368.600 31.770 370.600 ;
        RECT 39.770 368.600 41.770 370.600 ;
        RECT 43.770 368.600 45.770 370.600 ;
        RECT 47.770 368.600 49.770 370.600 ;
        RECT 51.770 368.600 53.770 370.600 ;
        RECT 55.770 368.600 65.770 370.600 ;
        RECT 29.770 366.600 47.770 368.600 ;
        RECT 49.770 366.600 63.770 368.600 ;
        RECT 45.770 364.600 51.770 366.600 ;
        RECT 5.000 60.000 25.000 70.000 ;
        RECT 85.000 30.000 105.000 40.000 ;
        RECT 85.000 5.000 105.000 25.000 ;
        RECT 499.200 0.000 500.800 500.000 ;
  END
END Art
END LIBRARY

