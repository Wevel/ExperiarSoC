VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ExperiarCore
  CLASS BLOCK ;
  FOREIGN ExperiarCore ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 800.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END addr0[8]
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END addr1[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END clk0
  PIN clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END clk1
  PIN coreIndex[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 796.000 6.350 800.000 ;
    END
  END coreIndex[0]
  PIN coreIndex[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 796.000 18.770 800.000 ;
    END
  END coreIndex[1]
  PIN coreIndex[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 796.000 31.650 800.000 ;
    END
  END coreIndex[2]
  PIN coreIndex[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 796.000 44.530 800.000 ;
    END
  END coreIndex[3]
  PIN coreIndex[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 796.000 57.410 800.000 ;
    END
  END coreIndex[4]
  PIN coreIndex[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 796.000 70.290 800.000 ;
    END
  END coreIndex[5]
  PIN coreIndex[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 796.000 83.170 800.000 ;
    END
  END coreIndex[6]
  PIN coreIndex[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 796.000 96.050 800.000 ;
    END
  END coreIndex[7]
  PIN core_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 8.880 500.000 9.480 ;
    END
  END core_wb_ack_i
  PIN core_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 32.680 500.000 33.280 ;
    END
  END core_wb_adr_o[0]
  PIN core_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 167.320 500.000 167.920 ;
    END
  END core_wb_adr_o[10]
  PIN core_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 178.880 500.000 179.480 ;
    END
  END core_wb_adr_o[11]
  PIN core_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 191.120 500.000 191.720 ;
    END
  END core_wb_adr_o[12]
  PIN core_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 202.680 500.000 203.280 ;
    END
  END core_wb_adr_o[13]
  PIN core_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 214.920 500.000 215.520 ;
    END
  END core_wb_adr_o[14]
  PIN core_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 226.480 500.000 227.080 ;
    END
  END core_wb_adr_o[15]
  PIN core_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 238.720 500.000 239.320 ;
    END
  END core_wb_adr_o[16]
  PIN core_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 250.280 500.000 250.880 ;
    END
  END core_wb_adr_o[17]
  PIN core_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 262.520 500.000 263.120 ;
    END
  END core_wb_adr_o[18]
  PIN core_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 274.080 500.000 274.680 ;
    END
  END core_wb_adr_o[19]
  PIN core_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 48.320 500.000 48.920 ;
    END
  END core_wb_adr_o[1]
  PIN core_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 286.320 500.000 286.920 ;
    END
  END core_wb_adr_o[20]
  PIN core_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 297.880 500.000 298.480 ;
    END
  END core_wb_adr_o[21]
  PIN core_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 310.120 500.000 310.720 ;
    END
  END core_wb_adr_o[22]
  PIN core_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 321.680 500.000 322.280 ;
    END
  END core_wb_adr_o[23]
  PIN core_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 333.920 500.000 334.520 ;
    END
  END core_wb_adr_o[24]
  PIN core_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 345.480 500.000 346.080 ;
    END
  END core_wb_adr_o[25]
  PIN core_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 357.040 500.000 357.640 ;
    END
  END core_wb_adr_o[26]
  PIN core_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 369.280 500.000 369.880 ;
    END
  END core_wb_adr_o[27]
  PIN core_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 64.640 500.000 65.240 ;
    END
  END core_wb_adr_o[2]
  PIN core_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 80.280 500.000 80.880 ;
    END
  END core_wb_adr_o[3]
  PIN core_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 95.920 500.000 96.520 ;
    END
  END core_wb_adr_o[4]
  PIN core_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 108.160 500.000 108.760 ;
    END
  END core_wb_adr_o[5]
  PIN core_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 119.720 500.000 120.320 ;
    END
  END core_wb_adr_o[6]
  PIN core_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 131.960 500.000 132.560 ;
    END
  END core_wb_adr_o[7]
  PIN core_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 143.520 500.000 144.120 ;
    END
  END core_wb_adr_o[8]
  PIN core_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 155.760 500.000 156.360 ;
    END
  END core_wb_adr_o[9]
  PIN core_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 12.960 500.000 13.560 ;
    END
  END core_wb_cyc_o
  PIN core_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 36.760 500.000 37.360 ;
    END
  END core_wb_data_i[0]
  PIN core_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 171.400 500.000 172.000 ;
    END
  END core_wb_data_i[10]
  PIN core_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 182.960 500.000 183.560 ;
    END
  END core_wb_data_i[11]
  PIN core_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 195.200 500.000 195.800 ;
    END
  END core_wb_data_i[12]
  PIN core_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 206.760 500.000 207.360 ;
    END
  END core_wb_data_i[13]
  PIN core_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 219.000 500.000 219.600 ;
    END
  END core_wb_data_i[14]
  PIN core_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 230.560 500.000 231.160 ;
    END
  END core_wb_data_i[15]
  PIN core_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 242.800 500.000 243.400 ;
    END
  END core_wb_data_i[16]
  PIN core_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 254.360 500.000 254.960 ;
    END
  END core_wb_data_i[17]
  PIN core_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 266.600 500.000 267.200 ;
    END
  END core_wb_data_i[18]
  PIN core_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 278.160 500.000 278.760 ;
    END
  END core_wb_data_i[19]
  PIN core_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 52.400 500.000 53.000 ;
    END
  END core_wb_data_i[1]
  PIN core_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 289.720 500.000 290.320 ;
    END
  END core_wb_data_i[20]
  PIN core_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 301.960 500.000 302.560 ;
    END
  END core_wb_data_i[21]
  PIN core_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 313.520 500.000 314.120 ;
    END
  END core_wb_data_i[22]
  PIN core_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 325.760 500.000 326.360 ;
    END
  END core_wb_data_i[23]
  PIN core_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 337.320 500.000 337.920 ;
    END
  END core_wb_data_i[24]
  PIN core_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 349.560 500.000 350.160 ;
    END
  END core_wb_data_i[25]
  PIN core_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 361.120 500.000 361.720 ;
    END
  END core_wb_data_i[26]
  PIN core_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 373.360 500.000 373.960 ;
    END
  END core_wb_data_i[27]
  PIN core_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 380.840 500.000 381.440 ;
    END
  END core_wb_data_i[28]
  PIN core_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 389.000 500.000 389.600 ;
    END
  END core_wb_data_i[29]
  PIN core_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.040 500.000 68.640 ;
    END
  END core_wb_data_i[2]
  PIN core_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 397.160 500.000 397.760 ;
    END
  END core_wb_data_i[30]
  PIN core_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 404.640 500.000 405.240 ;
    END
  END core_wb_data_i[31]
  PIN core_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 84.360 500.000 84.960 ;
    END
  END core_wb_data_i[3]
  PIN core_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 100.000 500.000 100.600 ;
    END
  END core_wb_data_i[4]
  PIN core_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 112.240 500.000 112.840 ;
    END
  END core_wb_data_i[5]
  PIN core_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 123.800 500.000 124.400 ;
    END
  END core_wb_data_i[6]
  PIN core_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 135.360 500.000 135.960 ;
    END
  END core_wb_data_i[7]
  PIN core_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 147.600 500.000 148.200 ;
    END
  END core_wb_data_i[8]
  PIN core_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 159.160 500.000 159.760 ;
    END
  END core_wb_data_i[9]
  PIN core_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 40.840 500.000 41.440 ;
    END
  END core_wb_data_o[0]
  PIN core_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 175.480 500.000 176.080 ;
    END
  END core_wb_data_o[10]
  PIN core_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.040 500.000 187.640 ;
    END
  END core_wb_data_o[11]
  PIN core_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 199.280 500.000 199.880 ;
    END
  END core_wb_data_o[12]
  PIN core_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.840 500.000 211.440 ;
    END
  END core_wb_data_o[13]
  PIN core_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 223.080 500.000 223.680 ;
    END
  END core_wb_data_o[14]
  PIN core_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 234.640 500.000 235.240 ;
    END
  END core_wb_data_o[15]
  PIN core_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 246.200 500.000 246.800 ;
    END
  END core_wb_data_o[16]
  PIN core_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 258.440 500.000 259.040 ;
    END
  END core_wb_data_o[17]
  PIN core_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 270.000 500.000 270.600 ;
    END
  END core_wb_data_o[18]
  PIN core_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 282.240 500.000 282.840 ;
    END
  END core_wb_data_o[19]
  PIN core_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 56.480 500.000 57.080 ;
    END
  END core_wb_data_o[1]
  PIN core_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 293.800 500.000 294.400 ;
    END
  END core_wb_data_o[20]
  PIN core_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 306.040 500.000 306.640 ;
    END
  END core_wb_data_o[21]
  PIN core_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 317.600 500.000 318.200 ;
    END
  END core_wb_data_o[22]
  PIN core_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 329.840 500.000 330.440 ;
    END
  END core_wb_data_o[23]
  PIN core_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 341.400 500.000 342.000 ;
    END
  END core_wb_data_o[24]
  PIN core_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 353.640 500.000 354.240 ;
    END
  END core_wb_data_o[25]
  PIN core_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 365.200 500.000 365.800 ;
    END
  END core_wb_data_o[26]
  PIN core_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 377.440 500.000 378.040 ;
    END
  END core_wb_data_o[27]
  PIN core_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 384.920 500.000 385.520 ;
    END
  END core_wb_data_o[28]
  PIN core_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 393.080 500.000 393.680 ;
    END
  END core_wb_data_o[29]
  PIN core_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 72.120 500.000 72.720 ;
    END
  END core_wb_data_o[2]
  PIN core_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 401.240 500.000 401.840 ;
    END
  END core_wb_data_o[30]
  PIN core_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 408.720 500.000 409.320 ;
    END
  END core_wb_data_o[31]
  PIN core_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 88.440 500.000 89.040 ;
    END
  END core_wb_data_o[3]
  PIN core_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 104.080 500.000 104.680 ;
    END
  END core_wb_data_o[4]
  PIN core_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 115.640 500.000 116.240 ;
    END
  END core_wb_data_o[5]
  PIN core_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 127.880 500.000 128.480 ;
    END
  END core_wb_data_o[6]
  PIN core_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 139.440 500.000 140.040 ;
    END
  END core_wb_data_o[7]
  PIN core_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 151.680 500.000 152.280 ;
    END
  END core_wb_data_o[8]
  PIN core_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 163.240 500.000 163.840 ;
    END
  END core_wb_data_o[9]
  PIN core_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 17.040 500.000 17.640 ;
    END
  END core_wb_error_i
  PIN core_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.920 500.000 45.520 ;
    END
  END core_wb_sel_o[0]
  PIN core_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 60.560 500.000 61.160 ;
    END
  END core_wb_sel_o[1]
  PIN core_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 76.200 500.000 76.800 ;
    END
  END core_wb_sel_o[2]
  PIN core_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 91.840 500.000 92.440 ;
    END
  END core_wb_sel_o[3]
  PIN core_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 21.120 500.000 21.720 ;
    END
  END core_wb_stall_i
  PIN core_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 24.520 500.000 25.120 ;
    END
  END core_wb_stb_o
  PIN core_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 28.600 500.000 29.200 ;
    END
  END core_wb_we_o
  PIN csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END csb0[0]
  PIN csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END csb0[1]
  PIN csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END csb1[0]
  PIN csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END csb1[1]
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END din0[9]
  PIN dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END dout0[32]
  PIN dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END dout0[33]
  PIN dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END dout0[34]
  PIN dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END dout0[35]
  PIN dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END dout0[36]
  PIN dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END dout0[37]
  PIN dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END dout0[38]
  PIN dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END dout0[39]
  PIN dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END dout0[3]
  PIN dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END dout0[40]
  PIN dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END dout0[41]
  PIN dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END dout0[42]
  PIN dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END dout0[43]
  PIN dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END dout0[44]
  PIN dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END dout0[45]
  PIN dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END dout0[46]
  PIN dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END dout0[47]
  PIN dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END dout0[48]
  PIN dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END dout0[49]
  PIN dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END dout0[4]
  PIN dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END dout0[50]
  PIN dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END dout0[51]
  PIN dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END dout0[52]
  PIN dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END dout0[53]
  PIN dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END dout0[54]
  PIN dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END dout0[55]
  PIN dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END dout0[56]
  PIN dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END dout0[57]
  PIN dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.760 4.000 462.360 ;
    END
  END dout0[58]
  PIN dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END dout0[59]
  PIN dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END dout0[5]
  PIN dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END dout0[60]
  PIN dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END dout0[61]
  PIN dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END dout0[62]
  PIN dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END dout0[63]
  PIN dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 577.360 4.000 577.960 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.000 4.000 644.600 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 4.000 648.680 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END dout1[31]
  PIN dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END dout1[32]
  PIN dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END dout1[33]
  PIN dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END dout1[34]
  PIN dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END dout1[35]
  PIN dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 685.480 4.000 686.080 ;
    END
  END dout1[36]
  PIN dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END dout1[37]
  PIN dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END dout1[38]
  PIN dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END dout1[39]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END dout1[3]
  PIN dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END dout1[40]
  PIN dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END dout1[41]
  PIN dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END dout1[42]
  PIN dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.720 4.000 715.320 ;
    END
  END dout1[43]
  PIN dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.800 4.000 719.400 ;
    END
  END dout1[44]
  PIN dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END dout1[45]
  PIN dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.960 4.000 727.560 ;
    END
  END dout1[46]
  PIN dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END dout1[47]
  PIN dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.120 4.000 735.720 ;
    END
  END dout1[48]
  PIN dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.200 4.000 739.800 ;
    END
  END dout1[49]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END dout1[4]
  PIN dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END dout1[50]
  PIN dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 747.360 4.000 747.960 ;
    END
  END dout1[51]
  PIN dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END dout1[52]
  PIN dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END dout1[53]
  PIN dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END dout1[54]
  PIN dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END dout1[55]
  PIN dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END dout1[56]
  PIN dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 772.520 4.000 773.120 ;
    END
  END dout1[57]
  PIN dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END dout1[58]
  PIN dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END dout1[59]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END dout1[5]
  PIN dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END dout1[60]
  PIN dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END dout1[61]
  PIN dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END dout1[62]
  PIN dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END dout1[63]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.120 4.000 565.720 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.200 4.000 569.800 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END dout1[9]
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END irq[0]
  PIN irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 0.000 450.710 4.000 ;
    END
  END irq[10]
  PIN irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END irq[11]
  PIN irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END irq[12]
  PIN irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END irq[13]
  PIN irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END irq[14]
  PIN irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END irq[15]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 0.000 370.210 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END irq[5]
  PIN irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END irq[6]
  PIN irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END irq[7]
  PIN irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END irq[8]
  PIN irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END irq[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END jtag_tms
  PIN localMemory_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 412.800 500.000 413.400 ;
    END
  END localMemory_wb_ack_o
  PIN localMemory_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 436.600 500.000 437.200 ;
    END
  END localMemory_wb_adr_i[0]
  PIN localMemory_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 571.240 500.000 571.840 ;
    END
  END localMemory_wb_adr_i[10]
  PIN localMemory_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 582.800 500.000 583.400 ;
    END
  END localMemory_wb_adr_i[11]
  PIN localMemory_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 595.040 500.000 595.640 ;
    END
  END localMemory_wb_adr_i[12]
  PIN localMemory_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 606.600 500.000 607.200 ;
    END
  END localMemory_wb_adr_i[13]
  PIN localMemory_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 618.840 500.000 619.440 ;
    END
  END localMemory_wb_adr_i[14]
  PIN localMemory_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 630.400 500.000 631.000 ;
    END
  END localMemory_wb_adr_i[15]
  PIN localMemory_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 642.640 500.000 643.240 ;
    END
  END localMemory_wb_adr_i[16]
  PIN localMemory_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 654.200 500.000 654.800 ;
    END
  END localMemory_wb_adr_i[17]
  PIN localMemory_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 666.440 500.000 667.040 ;
    END
  END localMemory_wb_adr_i[18]
  PIN localMemory_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 678.000 500.000 678.600 ;
    END
  END localMemory_wb_adr_i[19]
  PIN localMemory_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 452.240 500.000 452.840 ;
    END
  END localMemory_wb_adr_i[1]
  PIN localMemory_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 689.560 500.000 690.160 ;
    END
  END localMemory_wb_adr_i[20]
  PIN localMemory_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 701.800 500.000 702.400 ;
    END
  END localMemory_wb_adr_i[21]
  PIN localMemory_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 713.360 500.000 713.960 ;
    END
  END localMemory_wb_adr_i[22]
  PIN localMemory_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 725.600 500.000 726.200 ;
    END
  END localMemory_wb_adr_i[23]
  PIN localMemory_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 467.880 500.000 468.480 ;
    END
  END localMemory_wb_adr_i[2]
  PIN localMemory_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 484.200 500.000 484.800 ;
    END
  END localMemory_wb_adr_i[3]
  PIN localMemory_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 499.840 500.000 500.440 ;
    END
  END localMemory_wb_adr_i[4]
  PIN localMemory_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 512.080 500.000 512.680 ;
    END
  END localMemory_wb_adr_i[5]
  PIN localMemory_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 523.640 500.000 524.240 ;
    END
  END localMemory_wb_adr_i[6]
  PIN localMemory_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 535.200 500.000 535.800 ;
    END
  END localMemory_wb_adr_i[7]
  PIN localMemory_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 547.440 500.000 548.040 ;
    END
  END localMemory_wb_adr_i[8]
  PIN localMemory_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 559.000 500.000 559.600 ;
    END
  END localMemory_wb_adr_i[9]
  PIN localMemory_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 416.880 500.000 417.480 ;
    END
  END localMemory_wb_cyc_i
  PIN localMemory_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 440.680 500.000 441.280 ;
    END
  END localMemory_wb_data_i[0]
  PIN localMemory_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 575.320 500.000 575.920 ;
    END
  END localMemory_wb_data_i[10]
  PIN localMemory_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 586.880 500.000 587.480 ;
    END
  END localMemory_wb_data_i[11]
  PIN localMemory_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 599.120 500.000 599.720 ;
    END
  END localMemory_wb_data_i[12]
  PIN localMemory_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 610.680 500.000 611.280 ;
    END
  END localMemory_wb_data_i[13]
  PIN localMemory_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 622.920 500.000 623.520 ;
    END
  END localMemory_wb_data_i[14]
  PIN localMemory_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 634.480 500.000 635.080 ;
    END
  END localMemory_wb_data_i[15]
  PIN localMemory_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 646.040 500.000 646.640 ;
    END
  END localMemory_wb_data_i[16]
  PIN localMemory_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 658.280 500.000 658.880 ;
    END
  END localMemory_wb_data_i[17]
  PIN localMemory_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 669.840 500.000 670.440 ;
    END
  END localMemory_wb_data_i[18]
  PIN localMemory_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 682.080 500.000 682.680 ;
    END
  END localMemory_wb_data_i[19]
  PIN localMemory_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 456.320 500.000 456.920 ;
    END
  END localMemory_wb_data_i[1]
  PIN localMemory_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 693.640 500.000 694.240 ;
    END
  END localMemory_wb_data_i[20]
  PIN localMemory_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 705.880 500.000 706.480 ;
    END
  END localMemory_wb_data_i[21]
  PIN localMemory_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 717.440 500.000 718.040 ;
    END
  END localMemory_wb_data_i[22]
  PIN localMemory_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 729.680 500.000 730.280 ;
    END
  END localMemory_wb_data_i[23]
  PIN localMemory_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 737.160 500.000 737.760 ;
    END
  END localMemory_wb_data_i[24]
  PIN localMemory_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 745.320 500.000 745.920 ;
    END
  END localMemory_wb_data_i[25]
  PIN localMemory_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 753.480 500.000 754.080 ;
    END
  END localMemory_wb_data_i[26]
  PIN localMemory_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 760.960 500.000 761.560 ;
    END
  END localMemory_wb_data_i[27]
  PIN localMemory_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 769.120 500.000 769.720 ;
    END
  END localMemory_wb_data_i[28]
  PIN localMemory_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 777.280 500.000 777.880 ;
    END
  END localMemory_wb_data_i[29]
  PIN localMemory_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 471.960 500.000 472.560 ;
    END
  END localMemory_wb_data_i[2]
  PIN localMemory_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 784.760 500.000 785.360 ;
    END
  END localMemory_wb_data_i[30]
  PIN localMemory_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 792.920 500.000 793.520 ;
    END
  END localMemory_wb_data_i[31]
  PIN localMemory_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 488.280 500.000 488.880 ;
    END
  END localMemory_wb_data_i[3]
  PIN localMemory_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 503.920 500.000 504.520 ;
    END
  END localMemory_wb_data_i[4]
  PIN localMemory_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 515.480 500.000 516.080 ;
    END
  END localMemory_wb_data_i[5]
  PIN localMemory_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 527.720 500.000 528.320 ;
    END
  END localMemory_wb_data_i[6]
  PIN localMemory_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 539.280 500.000 539.880 ;
    END
  END localMemory_wb_data_i[7]
  PIN localMemory_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 551.520 500.000 552.120 ;
    END
  END localMemory_wb_data_i[8]
  PIN localMemory_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 563.080 500.000 563.680 ;
    END
  END localMemory_wb_data_i[9]
  PIN localMemory_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 444.760 500.000 445.360 ;
    END
  END localMemory_wb_data_o[0]
  PIN localMemory_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 578.720 500.000 579.320 ;
    END
  END localMemory_wb_data_o[10]
  PIN localMemory_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 590.960 500.000 591.560 ;
    END
  END localMemory_wb_data_o[11]
  PIN localMemory_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 602.520 500.000 603.120 ;
    END
  END localMemory_wb_data_o[12]
  PIN localMemory_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 614.760 500.000 615.360 ;
    END
  END localMemory_wb_data_o[13]
  PIN localMemory_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 626.320 500.000 626.920 ;
    END
  END localMemory_wb_data_o[14]
  PIN localMemory_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 638.560 500.000 639.160 ;
    END
  END localMemory_wb_data_o[15]
  PIN localMemory_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 650.120 500.000 650.720 ;
    END
  END localMemory_wb_data_o[16]
  PIN localMemory_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 662.360 500.000 662.960 ;
    END
  END localMemory_wb_data_o[17]
  PIN localMemory_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 673.920 500.000 674.520 ;
    END
  END localMemory_wb_data_o[18]
  PIN localMemory_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 686.160 500.000 686.760 ;
    END
  END localMemory_wb_data_o[19]
  PIN localMemory_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 460.400 500.000 461.000 ;
    END
  END localMemory_wb_data_o[1]
  PIN localMemory_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 697.720 500.000 698.320 ;
    END
  END localMemory_wb_data_o[20]
  PIN localMemory_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 709.960 500.000 710.560 ;
    END
  END localMemory_wb_data_o[21]
  PIN localMemory_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 721.520 500.000 722.120 ;
    END
  END localMemory_wb_data_o[22]
  PIN localMemory_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 733.760 500.000 734.360 ;
    END
  END localMemory_wb_data_o[23]
  PIN localMemory_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 741.240 500.000 741.840 ;
    END
  END localMemory_wb_data_o[24]
  PIN localMemory_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 749.400 500.000 750.000 ;
    END
  END localMemory_wb_data_o[25]
  PIN localMemory_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 756.880 500.000 757.480 ;
    END
  END localMemory_wb_data_o[26]
  PIN localMemory_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 765.040 500.000 765.640 ;
    END
  END localMemory_wb_data_o[27]
  PIN localMemory_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 773.200 500.000 773.800 ;
    END
  END localMemory_wb_data_o[28]
  PIN localMemory_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 780.680 500.000 781.280 ;
    END
  END localMemory_wb_data_o[29]
  PIN localMemory_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 476.040 500.000 476.640 ;
    END
  END localMemory_wb_data_o[2]
  PIN localMemory_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 788.840 500.000 789.440 ;
    END
  END localMemory_wb_data_o[30]
  PIN localMemory_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 797.000 500.000 797.600 ;
    END
  END localMemory_wb_data_o[31]
  PIN localMemory_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 491.680 500.000 492.280 ;
    END
  END localMemory_wb_data_o[3]
  PIN localMemory_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 508.000 500.000 508.600 ;
    END
  END localMemory_wb_data_o[4]
  PIN localMemory_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 519.560 500.000 520.160 ;
    END
  END localMemory_wb_data_o[5]
  PIN localMemory_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 531.800 500.000 532.400 ;
    END
  END localMemory_wb_data_o[6]
  PIN localMemory_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 543.360 500.000 543.960 ;
    END
  END localMemory_wb_data_o[7]
  PIN localMemory_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 555.600 500.000 556.200 ;
    END
  END localMemory_wb_data_o[8]
  PIN localMemory_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 567.160 500.000 567.760 ;
    END
  END localMemory_wb_data_o[9]
  PIN localMemory_wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 420.960 500.000 421.560 ;
    END
  END localMemory_wb_error_o
  PIN localMemory_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 448.160 500.000 448.760 ;
    END
  END localMemory_wb_sel_i[0]
  PIN localMemory_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 464.480 500.000 465.080 ;
    END
  END localMemory_wb_sel_i[1]
  PIN localMemory_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 480.120 500.000 480.720 ;
    END
  END localMemory_wb_sel_i[2]
  PIN localMemory_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 495.760 500.000 496.360 ;
    END
  END localMemory_wb_sel_i[3]
  PIN localMemory_wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 424.360 500.000 424.960 ;
    END
  END localMemory_wb_stall_o
  PIN localMemory_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 428.440 500.000 429.040 ;
    END
  END localMemory_wb_stb_i
  PIN localMemory_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 432.520 500.000 433.120 ;
    END
  END localMemory_wb_we_i
  PIN manufacturerID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 796.000 108.470 800.000 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 796.000 236.810 800.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 796.000 121.350 800.000 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 796.000 134.230 800.000 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 796.000 147.110 800.000 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 796.000 159.990 800.000 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 796.000 172.870 800.000 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 796.000 185.750 800.000 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 796.000 198.630 800.000 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 796.000 211.050 800.000 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 796.000 223.930 800.000 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 796.000 249.690 800.000 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 796.000 378.030 800.000 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 796.000 390.910 800.000 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 796.000 403.790 800.000 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 796.000 416.210 800.000 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 796.000 429.090 800.000 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 796.000 441.970 800.000 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 796.000 262.570 800.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 796.000 275.450 800.000 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 796.000 288.330 800.000 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 796.000 301.210 800.000 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 796.000 313.630 800.000 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 796.000 326.510 800.000 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 796.000 339.390 800.000 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 796.000 352.270 800.000 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 796.000 365.150 800.000 ;
    END
  END partID[9]
  PIN probe_env[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END probe_env[0]
  PIN probe_env[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END probe_env[1]
  PIN probe_jtagInstruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END probe_jtagInstruction[0]
  PIN probe_jtagInstruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END probe_jtagInstruction[1]
  PIN probe_jtagInstruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END probe_jtagInstruction[2]
  PIN probe_jtagInstruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END probe_jtagInstruction[3]
  PIN probe_jtagInstruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END probe_jtagInstruction[4]
  PIN probe_programCounter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END probe_programCounter[0]
  PIN probe_programCounter[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END probe_programCounter[10]
  PIN probe_programCounter[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END probe_programCounter[11]
  PIN probe_programCounter[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END probe_programCounter[12]
  PIN probe_programCounter[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END probe_programCounter[13]
  PIN probe_programCounter[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END probe_programCounter[14]
  PIN probe_programCounter[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END probe_programCounter[15]
  PIN probe_programCounter[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END probe_programCounter[16]
  PIN probe_programCounter[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END probe_programCounter[17]
  PIN probe_programCounter[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END probe_programCounter[18]
  PIN probe_programCounter[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END probe_programCounter[19]
  PIN probe_programCounter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END probe_programCounter[1]
  PIN probe_programCounter[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END probe_programCounter[20]
  PIN probe_programCounter[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END probe_programCounter[21]
  PIN probe_programCounter[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END probe_programCounter[22]
  PIN probe_programCounter[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END probe_programCounter[23]
  PIN probe_programCounter[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END probe_programCounter[24]
  PIN probe_programCounter[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END probe_programCounter[25]
  PIN probe_programCounter[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END probe_programCounter[26]
  PIN probe_programCounter[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END probe_programCounter[27]
  PIN probe_programCounter[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END probe_programCounter[28]
  PIN probe_programCounter[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END probe_programCounter[29]
  PIN probe_programCounter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END probe_programCounter[2]
  PIN probe_programCounter[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END probe_programCounter[30]
  PIN probe_programCounter[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END probe_programCounter[31]
  PIN probe_programCounter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END probe_programCounter[3]
  PIN probe_programCounter[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END probe_programCounter[4]
  PIN probe_programCounter[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END probe_programCounter[5]
  PIN probe_programCounter[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END probe_programCounter[6]
  PIN probe_programCounter[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END probe_programCounter[7]
  PIN probe_programCounter[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END probe_programCounter[8]
  PIN probe_programCounter[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END probe_programCounter[9]
  PIN probe_state
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END probe_state
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.570 796.000 454.850 800.000 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 796.000 467.730 800.000 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 796.000 480.610 800.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 796.000 493.490 800.000 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 1.400 500.000 2.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 4.800 500.000 5.400 ;
    END
  END wb_rst_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 788.885 ;
      LAYER met1 ;
        RECT 0.070 6.500 499.950 794.540 ;
      LAYER met2 ;
        RECT 0.090 795.720 5.790 797.485 ;
        RECT 6.630 795.720 18.210 797.485 ;
        RECT 19.050 795.720 31.090 797.485 ;
        RECT 31.930 795.720 43.970 797.485 ;
        RECT 44.810 795.720 56.850 797.485 ;
        RECT 57.690 795.720 69.730 797.485 ;
        RECT 70.570 795.720 82.610 797.485 ;
        RECT 83.450 795.720 95.490 797.485 ;
        RECT 96.330 795.720 107.910 797.485 ;
        RECT 108.750 795.720 120.790 797.485 ;
        RECT 121.630 795.720 133.670 797.485 ;
        RECT 134.510 795.720 146.550 797.485 ;
        RECT 147.390 795.720 159.430 797.485 ;
        RECT 160.270 795.720 172.310 797.485 ;
        RECT 173.150 795.720 185.190 797.485 ;
        RECT 186.030 795.720 198.070 797.485 ;
        RECT 198.910 795.720 210.490 797.485 ;
        RECT 211.330 795.720 223.370 797.485 ;
        RECT 224.210 795.720 236.250 797.485 ;
        RECT 237.090 795.720 249.130 797.485 ;
        RECT 249.970 795.720 262.010 797.485 ;
        RECT 262.850 795.720 274.890 797.485 ;
        RECT 275.730 795.720 287.770 797.485 ;
        RECT 288.610 795.720 300.650 797.485 ;
        RECT 301.490 795.720 313.070 797.485 ;
        RECT 313.910 795.720 325.950 797.485 ;
        RECT 326.790 795.720 338.830 797.485 ;
        RECT 339.670 795.720 351.710 797.485 ;
        RECT 352.550 795.720 364.590 797.485 ;
        RECT 365.430 795.720 377.470 797.485 ;
        RECT 378.310 795.720 390.350 797.485 ;
        RECT 391.190 795.720 403.230 797.485 ;
        RECT 404.070 795.720 415.650 797.485 ;
        RECT 416.490 795.720 428.530 797.485 ;
        RECT 429.370 795.720 441.410 797.485 ;
        RECT 442.250 795.720 454.290 797.485 ;
        RECT 455.130 795.720 467.170 797.485 ;
        RECT 468.010 795.720 480.050 797.485 ;
        RECT 480.890 795.720 492.930 797.485 ;
        RECT 493.770 795.720 499.920 797.485 ;
        RECT 0.090 4.280 499.920 795.720 ;
        RECT 0.090 1.515 3.950 4.280 ;
        RECT 4.790 1.515 12.690 4.280 ;
        RECT 13.530 1.515 21.430 4.280 ;
        RECT 22.270 1.515 30.630 4.280 ;
        RECT 31.470 1.515 39.370 4.280 ;
        RECT 40.210 1.515 48.570 4.280 ;
        RECT 49.410 1.515 57.310 4.280 ;
        RECT 58.150 1.515 66.050 4.280 ;
        RECT 66.890 1.515 75.250 4.280 ;
        RECT 76.090 1.515 83.990 4.280 ;
        RECT 84.830 1.515 93.190 4.280 ;
        RECT 94.030 1.515 101.930 4.280 ;
        RECT 102.770 1.515 110.670 4.280 ;
        RECT 111.510 1.515 119.870 4.280 ;
        RECT 120.710 1.515 128.610 4.280 ;
        RECT 129.450 1.515 137.810 4.280 ;
        RECT 138.650 1.515 146.550 4.280 ;
        RECT 147.390 1.515 155.290 4.280 ;
        RECT 156.130 1.515 164.490 4.280 ;
        RECT 165.330 1.515 173.230 4.280 ;
        RECT 174.070 1.515 182.430 4.280 ;
        RECT 183.270 1.515 191.170 4.280 ;
        RECT 192.010 1.515 200.370 4.280 ;
        RECT 201.210 1.515 209.110 4.280 ;
        RECT 209.950 1.515 217.850 4.280 ;
        RECT 218.690 1.515 227.050 4.280 ;
        RECT 227.890 1.515 235.790 4.280 ;
        RECT 236.630 1.515 244.990 4.280 ;
        RECT 245.830 1.515 253.730 4.280 ;
        RECT 254.570 1.515 262.470 4.280 ;
        RECT 263.310 1.515 271.670 4.280 ;
        RECT 272.510 1.515 280.410 4.280 ;
        RECT 281.250 1.515 289.610 4.280 ;
        RECT 290.450 1.515 298.350 4.280 ;
        RECT 299.190 1.515 307.090 4.280 ;
        RECT 307.930 1.515 316.290 4.280 ;
        RECT 317.130 1.515 325.030 4.280 ;
        RECT 325.870 1.515 334.230 4.280 ;
        RECT 335.070 1.515 342.970 4.280 ;
        RECT 343.810 1.515 352.170 4.280 ;
        RECT 353.010 1.515 360.910 4.280 ;
        RECT 361.750 1.515 369.650 4.280 ;
        RECT 370.490 1.515 378.850 4.280 ;
        RECT 379.690 1.515 387.590 4.280 ;
        RECT 388.430 1.515 396.790 4.280 ;
        RECT 397.630 1.515 405.530 4.280 ;
        RECT 406.370 1.515 414.270 4.280 ;
        RECT 415.110 1.515 423.470 4.280 ;
        RECT 424.310 1.515 432.210 4.280 ;
        RECT 433.050 1.515 441.410 4.280 ;
        RECT 442.250 1.515 450.150 4.280 ;
        RECT 450.990 1.515 458.890 4.280 ;
        RECT 459.730 1.515 468.090 4.280 ;
        RECT 468.930 1.515 476.830 4.280 ;
        RECT 477.670 1.515 486.030 4.280 ;
        RECT 486.870 1.515 494.770 4.280 ;
        RECT 495.610 1.515 499.920 4.280 ;
      LAYER met3 ;
        RECT 4.400 796.600 495.600 797.465 ;
        RECT 0.065 793.920 499.495 796.600 ;
        RECT 4.400 792.520 495.600 793.920 ;
        RECT 0.065 789.840 499.495 792.520 ;
        RECT 4.400 788.440 495.600 789.840 ;
        RECT 0.065 785.760 499.495 788.440 ;
        RECT 4.400 784.360 495.600 785.760 ;
        RECT 0.065 781.680 499.495 784.360 ;
        RECT 4.400 780.280 495.600 781.680 ;
        RECT 0.065 778.280 499.495 780.280 ;
        RECT 0.065 777.600 495.600 778.280 ;
        RECT 4.400 776.880 495.600 777.600 ;
        RECT 4.400 776.200 499.495 776.880 ;
        RECT 0.065 774.200 499.495 776.200 ;
        RECT 0.065 773.520 495.600 774.200 ;
        RECT 4.400 772.800 495.600 773.520 ;
        RECT 4.400 772.120 499.495 772.800 ;
        RECT 0.065 770.120 499.495 772.120 ;
        RECT 0.065 769.440 495.600 770.120 ;
        RECT 4.400 768.720 495.600 769.440 ;
        RECT 4.400 768.040 499.495 768.720 ;
        RECT 0.065 766.040 499.495 768.040 ;
        RECT 0.065 765.360 495.600 766.040 ;
        RECT 4.400 764.640 495.600 765.360 ;
        RECT 4.400 763.960 499.495 764.640 ;
        RECT 0.065 761.960 499.495 763.960 ;
        RECT 0.065 761.280 495.600 761.960 ;
        RECT 4.400 760.560 495.600 761.280 ;
        RECT 4.400 759.880 499.495 760.560 ;
        RECT 0.065 757.880 499.495 759.880 ;
        RECT 0.065 756.520 495.600 757.880 ;
        RECT 4.400 756.480 495.600 756.520 ;
        RECT 4.400 755.120 499.495 756.480 ;
        RECT 0.065 754.480 499.495 755.120 ;
        RECT 0.065 753.080 495.600 754.480 ;
        RECT 0.065 752.440 499.495 753.080 ;
        RECT 4.400 751.040 499.495 752.440 ;
        RECT 0.065 750.400 499.495 751.040 ;
        RECT 0.065 749.000 495.600 750.400 ;
        RECT 0.065 748.360 499.495 749.000 ;
        RECT 4.400 746.960 499.495 748.360 ;
        RECT 0.065 746.320 499.495 746.960 ;
        RECT 0.065 744.920 495.600 746.320 ;
        RECT 0.065 744.280 499.495 744.920 ;
        RECT 4.400 742.880 499.495 744.280 ;
        RECT 0.065 742.240 499.495 742.880 ;
        RECT 0.065 740.840 495.600 742.240 ;
        RECT 0.065 740.200 499.495 740.840 ;
        RECT 4.400 738.800 499.495 740.200 ;
        RECT 0.065 738.160 499.495 738.800 ;
        RECT 0.065 736.760 495.600 738.160 ;
        RECT 0.065 736.120 499.495 736.760 ;
        RECT 4.400 734.760 499.495 736.120 ;
        RECT 4.400 734.720 495.600 734.760 ;
        RECT 0.065 733.360 495.600 734.720 ;
        RECT 0.065 732.040 499.495 733.360 ;
        RECT 4.400 730.680 499.495 732.040 ;
        RECT 4.400 730.640 495.600 730.680 ;
        RECT 0.065 729.280 495.600 730.640 ;
        RECT 0.065 727.960 499.495 729.280 ;
        RECT 4.400 726.600 499.495 727.960 ;
        RECT 4.400 726.560 495.600 726.600 ;
        RECT 0.065 725.200 495.600 726.560 ;
        RECT 0.065 723.880 499.495 725.200 ;
        RECT 4.400 722.520 499.495 723.880 ;
        RECT 4.400 722.480 495.600 722.520 ;
        RECT 0.065 721.120 495.600 722.480 ;
        RECT 0.065 719.800 499.495 721.120 ;
        RECT 4.400 718.440 499.495 719.800 ;
        RECT 4.400 718.400 495.600 718.440 ;
        RECT 0.065 717.040 495.600 718.400 ;
        RECT 0.065 715.720 499.495 717.040 ;
        RECT 4.400 714.360 499.495 715.720 ;
        RECT 4.400 714.320 495.600 714.360 ;
        RECT 0.065 712.960 495.600 714.320 ;
        RECT 0.065 710.960 499.495 712.960 ;
        RECT 4.400 709.560 495.600 710.960 ;
        RECT 0.065 706.880 499.495 709.560 ;
        RECT 4.400 705.480 495.600 706.880 ;
        RECT 0.065 702.800 499.495 705.480 ;
        RECT 4.400 701.400 495.600 702.800 ;
        RECT 0.065 698.720 499.495 701.400 ;
        RECT 4.400 697.320 495.600 698.720 ;
        RECT 0.065 694.640 499.495 697.320 ;
        RECT 4.400 693.240 495.600 694.640 ;
        RECT 0.065 690.560 499.495 693.240 ;
        RECT 4.400 689.160 495.600 690.560 ;
        RECT 0.065 687.160 499.495 689.160 ;
        RECT 0.065 686.480 495.600 687.160 ;
        RECT 4.400 685.760 495.600 686.480 ;
        RECT 4.400 685.080 499.495 685.760 ;
        RECT 0.065 683.080 499.495 685.080 ;
        RECT 0.065 682.400 495.600 683.080 ;
        RECT 4.400 681.680 495.600 682.400 ;
        RECT 4.400 681.000 499.495 681.680 ;
        RECT 0.065 679.000 499.495 681.000 ;
        RECT 0.065 678.320 495.600 679.000 ;
        RECT 4.400 677.600 495.600 678.320 ;
        RECT 4.400 676.920 499.495 677.600 ;
        RECT 0.065 674.920 499.495 676.920 ;
        RECT 0.065 674.240 495.600 674.920 ;
        RECT 4.400 673.520 495.600 674.240 ;
        RECT 4.400 672.840 499.495 673.520 ;
        RECT 0.065 670.840 499.495 672.840 ;
        RECT 0.065 670.160 495.600 670.840 ;
        RECT 4.400 669.440 495.600 670.160 ;
        RECT 4.400 668.760 499.495 669.440 ;
        RECT 0.065 667.440 499.495 668.760 ;
        RECT 0.065 666.040 495.600 667.440 ;
        RECT 0.065 665.400 499.495 666.040 ;
        RECT 4.400 664.000 499.495 665.400 ;
        RECT 0.065 663.360 499.495 664.000 ;
        RECT 0.065 661.960 495.600 663.360 ;
        RECT 0.065 661.320 499.495 661.960 ;
        RECT 4.400 659.920 499.495 661.320 ;
        RECT 0.065 659.280 499.495 659.920 ;
        RECT 0.065 657.880 495.600 659.280 ;
        RECT 0.065 657.240 499.495 657.880 ;
        RECT 4.400 655.840 499.495 657.240 ;
        RECT 0.065 655.200 499.495 655.840 ;
        RECT 0.065 653.800 495.600 655.200 ;
        RECT 0.065 653.160 499.495 653.800 ;
        RECT 4.400 651.760 499.495 653.160 ;
        RECT 0.065 651.120 499.495 651.760 ;
        RECT 0.065 649.720 495.600 651.120 ;
        RECT 0.065 649.080 499.495 649.720 ;
        RECT 4.400 647.680 499.495 649.080 ;
        RECT 0.065 647.040 499.495 647.680 ;
        RECT 0.065 645.640 495.600 647.040 ;
        RECT 0.065 645.000 499.495 645.640 ;
        RECT 4.400 643.640 499.495 645.000 ;
        RECT 4.400 643.600 495.600 643.640 ;
        RECT 0.065 642.240 495.600 643.600 ;
        RECT 0.065 640.920 499.495 642.240 ;
        RECT 4.400 639.560 499.495 640.920 ;
        RECT 4.400 639.520 495.600 639.560 ;
        RECT 0.065 638.160 495.600 639.520 ;
        RECT 0.065 636.840 499.495 638.160 ;
        RECT 4.400 635.480 499.495 636.840 ;
        RECT 4.400 635.440 495.600 635.480 ;
        RECT 0.065 634.080 495.600 635.440 ;
        RECT 0.065 632.760 499.495 634.080 ;
        RECT 4.400 631.400 499.495 632.760 ;
        RECT 4.400 631.360 495.600 631.400 ;
        RECT 0.065 630.000 495.600 631.360 ;
        RECT 0.065 628.680 499.495 630.000 ;
        RECT 4.400 627.320 499.495 628.680 ;
        RECT 4.400 627.280 495.600 627.320 ;
        RECT 0.065 625.920 495.600 627.280 ;
        RECT 0.065 623.920 499.495 625.920 ;
        RECT 4.400 622.520 495.600 623.920 ;
        RECT 0.065 619.840 499.495 622.520 ;
        RECT 4.400 618.440 495.600 619.840 ;
        RECT 0.065 615.760 499.495 618.440 ;
        RECT 4.400 614.360 495.600 615.760 ;
        RECT 0.065 611.680 499.495 614.360 ;
        RECT 4.400 610.280 495.600 611.680 ;
        RECT 0.065 607.600 499.495 610.280 ;
        RECT 4.400 606.200 495.600 607.600 ;
        RECT 0.065 603.520 499.495 606.200 ;
        RECT 4.400 602.120 495.600 603.520 ;
        RECT 0.065 600.120 499.495 602.120 ;
        RECT 0.065 599.440 495.600 600.120 ;
        RECT 4.400 598.720 495.600 599.440 ;
        RECT 4.400 598.040 499.495 598.720 ;
        RECT 0.065 596.040 499.495 598.040 ;
        RECT 0.065 595.360 495.600 596.040 ;
        RECT 4.400 594.640 495.600 595.360 ;
        RECT 4.400 593.960 499.495 594.640 ;
        RECT 0.065 591.960 499.495 593.960 ;
        RECT 0.065 591.280 495.600 591.960 ;
        RECT 4.400 590.560 495.600 591.280 ;
        RECT 4.400 589.880 499.495 590.560 ;
        RECT 0.065 587.880 499.495 589.880 ;
        RECT 0.065 587.200 495.600 587.880 ;
        RECT 4.400 586.480 495.600 587.200 ;
        RECT 4.400 585.800 499.495 586.480 ;
        RECT 0.065 583.800 499.495 585.800 ;
        RECT 0.065 583.120 495.600 583.800 ;
        RECT 4.400 582.400 495.600 583.120 ;
        RECT 4.400 581.720 499.495 582.400 ;
        RECT 0.065 579.720 499.495 581.720 ;
        RECT 0.065 578.360 495.600 579.720 ;
        RECT 4.400 578.320 495.600 578.360 ;
        RECT 4.400 576.960 499.495 578.320 ;
        RECT 0.065 576.320 499.495 576.960 ;
        RECT 0.065 574.920 495.600 576.320 ;
        RECT 0.065 574.280 499.495 574.920 ;
        RECT 4.400 572.880 499.495 574.280 ;
        RECT 0.065 572.240 499.495 572.880 ;
        RECT 0.065 570.840 495.600 572.240 ;
        RECT 0.065 570.200 499.495 570.840 ;
        RECT 4.400 568.800 499.495 570.200 ;
        RECT 0.065 568.160 499.495 568.800 ;
        RECT 0.065 566.760 495.600 568.160 ;
        RECT 0.065 566.120 499.495 566.760 ;
        RECT 4.400 564.720 499.495 566.120 ;
        RECT 0.065 564.080 499.495 564.720 ;
        RECT 0.065 562.680 495.600 564.080 ;
        RECT 0.065 562.040 499.495 562.680 ;
        RECT 4.400 560.640 499.495 562.040 ;
        RECT 0.065 560.000 499.495 560.640 ;
        RECT 0.065 558.600 495.600 560.000 ;
        RECT 0.065 557.960 499.495 558.600 ;
        RECT 4.400 556.600 499.495 557.960 ;
        RECT 4.400 556.560 495.600 556.600 ;
        RECT 0.065 555.200 495.600 556.560 ;
        RECT 0.065 553.880 499.495 555.200 ;
        RECT 4.400 552.520 499.495 553.880 ;
        RECT 4.400 552.480 495.600 552.520 ;
        RECT 0.065 551.120 495.600 552.480 ;
        RECT 0.065 549.800 499.495 551.120 ;
        RECT 4.400 548.440 499.495 549.800 ;
        RECT 4.400 548.400 495.600 548.440 ;
        RECT 0.065 547.040 495.600 548.400 ;
        RECT 0.065 545.720 499.495 547.040 ;
        RECT 4.400 544.360 499.495 545.720 ;
        RECT 4.400 544.320 495.600 544.360 ;
        RECT 0.065 542.960 495.600 544.320 ;
        RECT 0.065 541.640 499.495 542.960 ;
        RECT 4.400 540.280 499.495 541.640 ;
        RECT 4.400 540.240 495.600 540.280 ;
        RECT 0.065 538.880 495.600 540.240 ;
        RECT 0.065 537.560 499.495 538.880 ;
        RECT 4.400 536.200 499.495 537.560 ;
        RECT 4.400 536.160 495.600 536.200 ;
        RECT 0.065 534.800 495.600 536.160 ;
        RECT 0.065 532.800 499.495 534.800 ;
        RECT 4.400 531.400 495.600 532.800 ;
        RECT 0.065 528.720 499.495 531.400 ;
        RECT 4.400 527.320 495.600 528.720 ;
        RECT 0.065 524.640 499.495 527.320 ;
        RECT 4.400 523.240 495.600 524.640 ;
        RECT 0.065 520.560 499.495 523.240 ;
        RECT 4.400 519.160 495.600 520.560 ;
        RECT 0.065 516.480 499.495 519.160 ;
        RECT 4.400 515.080 495.600 516.480 ;
        RECT 0.065 513.080 499.495 515.080 ;
        RECT 0.065 512.400 495.600 513.080 ;
        RECT 4.400 511.680 495.600 512.400 ;
        RECT 4.400 511.000 499.495 511.680 ;
        RECT 0.065 509.000 499.495 511.000 ;
        RECT 0.065 508.320 495.600 509.000 ;
        RECT 4.400 507.600 495.600 508.320 ;
        RECT 4.400 506.920 499.495 507.600 ;
        RECT 0.065 504.920 499.495 506.920 ;
        RECT 0.065 504.240 495.600 504.920 ;
        RECT 4.400 503.520 495.600 504.240 ;
        RECT 4.400 502.840 499.495 503.520 ;
        RECT 0.065 500.840 499.495 502.840 ;
        RECT 0.065 500.160 495.600 500.840 ;
        RECT 4.400 499.440 495.600 500.160 ;
        RECT 4.400 498.760 499.495 499.440 ;
        RECT 0.065 496.760 499.495 498.760 ;
        RECT 0.065 496.080 495.600 496.760 ;
        RECT 4.400 495.360 495.600 496.080 ;
        RECT 4.400 494.680 499.495 495.360 ;
        RECT 0.065 492.680 499.495 494.680 ;
        RECT 0.065 492.000 495.600 492.680 ;
        RECT 4.400 491.280 495.600 492.000 ;
        RECT 4.400 490.600 499.495 491.280 ;
        RECT 0.065 489.280 499.495 490.600 ;
        RECT 0.065 487.880 495.600 489.280 ;
        RECT 0.065 487.240 499.495 487.880 ;
        RECT 4.400 485.840 499.495 487.240 ;
        RECT 0.065 485.200 499.495 485.840 ;
        RECT 0.065 483.800 495.600 485.200 ;
        RECT 0.065 483.160 499.495 483.800 ;
        RECT 4.400 481.760 499.495 483.160 ;
        RECT 0.065 481.120 499.495 481.760 ;
        RECT 0.065 479.720 495.600 481.120 ;
        RECT 0.065 479.080 499.495 479.720 ;
        RECT 4.400 477.680 499.495 479.080 ;
        RECT 0.065 477.040 499.495 477.680 ;
        RECT 0.065 475.640 495.600 477.040 ;
        RECT 0.065 475.000 499.495 475.640 ;
        RECT 4.400 473.600 499.495 475.000 ;
        RECT 0.065 472.960 499.495 473.600 ;
        RECT 0.065 471.560 495.600 472.960 ;
        RECT 0.065 470.920 499.495 471.560 ;
        RECT 4.400 469.520 499.495 470.920 ;
        RECT 0.065 468.880 499.495 469.520 ;
        RECT 0.065 467.480 495.600 468.880 ;
        RECT 0.065 466.840 499.495 467.480 ;
        RECT 4.400 465.480 499.495 466.840 ;
        RECT 4.400 465.440 495.600 465.480 ;
        RECT 0.065 464.080 495.600 465.440 ;
        RECT 0.065 462.760 499.495 464.080 ;
        RECT 4.400 461.400 499.495 462.760 ;
        RECT 4.400 461.360 495.600 461.400 ;
        RECT 0.065 460.000 495.600 461.360 ;
        RECT 0.065 458.680 499.495 460.000 ;
        RECT 4.400 457.320 499.495 458.680 ;
        RECT 4.400 457.280 495.600 457.320 ;
        RECT 0.065 455.920 495.600 457.280 ;
        RECT 0.065 454.600 499.495 455.920 ;
        RECT 4.400 453.240 499.495 454.600 ;
        RECT 4.400 453.200 495.600 453.240 ;
        RECT 0.065 451.840 495.600 453.200 ;
        RECT 0.065 450.520 499.495 451.840 ;
        RECT 4.400 449.160 499.495 450.520 ;
        RECT 4.400 449.120 495.600 449.160 ;
        RECT 0.065 447.760 495.600 449.120 ;
        RECT 0.065 445.760 499.495 447.760 ;
        RECT 4.400 444.360 495.600 445.760 ;
        RECT 0.065 441.680 499.495 444.360 ;
        RECT 4.400 440.280 495.600 441.680 ;
        RECT 0.065 437.600 499.495 440.280 ;
        RECT 4.400 436.200 495.600 437.600 ;
        RECT 0.065 433.520 499.495 436.200 ;
        RECT 4.400 432.120 495.600 433.520 ;
        RECT 0.065 429.440 499.495 432.120 ;
        RECT 4.400 428.040 495.600 429.440 ;
        RECT 0.065 425.360 499.495 428.040 ;
        RECT 4.400 423.960 495.600 425.360 ;
        RECT 0.065 421.960 499.495 423.960 ;
        RECT 0.065 421.280 495.600 421.960 ;
        RECT 4.400 420.560 495.600 421.280 ;
        RECT 4.400 419.880 499.495 420.560 ;
        RECT 0.065 417.880 499.495 419.880 ;
        RECT 0.065 417.200 495.600 417.880 ;
        RECT 4.400 416.480 495.600 417.200 ;
        RECT 4.400 415.800 499.495 416.480 ;
        RECT 0.065 413.800 499.495 415.800 ;
        RECT 0.065 413.120 495.600 413.800 ;
        RECT 4.400 412.400 495.600 413.120 ;
        RECT 4.400 411.720 499.495 412.400 ;
        RECT 0.065 409.720 499.495 411.720 ;
        RECT 0.065 409.040 495.600 409.720 ;
        RECT 4.400 408.320 495.600 409.040 ;
        RECT 4.400 407.640 499.495 408.320 ;
        RECT 0.065 405.640 499.495 407.640 ;
        RECT 0.065 404.960 495.600 405.640 ;
        RECT 4.400 404.240 495.600 404.960 ;
        RECT 4.400 403.560 499.495 404.240 ;
        RECT 0.065 402.240 499.495 403.560 ;
        RECT 0.065 400.840 495.600 402.240 ;
        RECT 0.065 400.200 499.495 400.840 ;
        RECT 4.400 398.800 499.495 400.200 ;
        RECT 0.065 398.160 499.495 398.800 ;
        RECT 0.065 396.760 495.600 398.160 ;
        RECT 0.065 396.120 499.495 396.760 ;
        RECT 4.400 394.720 499.495 396.120 ;
        RECT 0.065 394.080 499.495 394.720 ;
        RECT 0.065 392.680 495.600 394.080 ;
        RECT 0.065 392.040 499.495 392.680 ;
        RECT 4.400 390.640 499.495 392.040 ;
        RECT 0.065 390.000 499.495 390.640 ;
        RECT 0.065 388.600 495.600 390.000 ;
        RECT 0.065 387.960 499.495 388.600 ;
        RECT 4.400 386.560 499.495 387.960 ;
        RECT 0.065 385.920 499.495 386.560 ;
        RECT 0.065 384.520 495.600 385.920 ;
        RECT 0.065 383.880 499.495 384.520 ;
        RECT 4.400 382.480 499.495 383.880 ;
        RECT 0.065 381.840 499.495 382.480 ;
        RECT 0.065 380.440 495.600 381.840 ;
        RECT 0.065 379.800 499.495 380.440 ;
        RECT 4.400 378.440 499.495 379.800 ;
        RECT 4.400 378.400 495.600 378.440 ;
        RECT 0.065 377.040 495.600 378.400 ;
        RECT 0.065 375.720 499.495 377.040 ;
        RECT 4.400 374.360 499.495 375.720 ;
        RECT 4.400 374.320 495.600 374.360 ;
        RECT 0.065 372.960 495.600 374.320 ;
        RECT 0.065 371.640 499.495 372.960 ;
        RECT 4.400 370.280 499.495 371.640 ;
        RECT 4.400 370.240 495.600 370.280 ;
        RECT 0.065 368.880 495.600 370.240 ;
        RECT 0.065 367.560 499.495 368.880 ;
        RECT 4.400 366.200 499.495 367.560 ;
        RECT 4.400 366.160 495.600 366.200 ;
        RECT 0.065 364.800 495.600 366.160 ;
        RECT 0.065 363.480 499.495 364.800 ;
        RECT 4.400 362.120 499.495 363.480 ;
        RECT 4.400 362.080 495.600 362.120 ;
        RECT 0.065 360.720 495.600 362.080 ;
        RECT 0.065 359.400 499.495 360.720 ;
        RECT 4.400 358.040 499.495 359.400 ;
        RECT 4.400 358.000 495.600 358.040 ;
        RECT 0.065 356.640 495.600 358.000 ;
        RECT 0.065 354.640 499.495 356.640 ;
        RECT 4.400 353.240 495.600 354.640 ;
        RECT 0.065 350.560 499.495 353.240 ;
        RECT 4.400 349.160 495.600 350.560 ;
        RECT 0.065 346.480 499.495 349.160 ;
        RECT 4.400 345.080 495.600 346.480 ;
        RECT 0.065 342.400 499.495 345.080 ;
        RECT 4.400 341.000 495.600 342.400 ;
        RECT 0.065 338.320 499.495 341.000 ;
        RECT 4.400 336.920 495.600 338.320 ;
        RECT 0.065 334.920 499.495 336.920 ;
        RECT 0.065 334.240 495.600 334.920 ;
        RECT 4.400 333.520 495.600 334.240 ;
        RECT 4.400 332.840 499.495 333.520 ;
        RECT 0.065 330.840 499.495 332.840 ;
        RECT 0.065 330.160 495.600 330.840 ;
        RECT 4.400 329.440 495.600 330.160 ;
        RECT 4.400 328.760 499.495 329.440 ;
        RECT 0.065 326.760 499.495 328.760 ;
        RECT 0.065 326.080 495.600 326.760 ;
        RECT 4.400 325.360 495.600 326.080 ;
        RECT 4.400 324.680 499.495 325.360 ;
        RECT 0.065 322.680 499.495 324.680 ;
        RECT 0.065 322.000 495.600 322.680 ;
        RECT 4.400 321.280 495.600 322.000 ;
        RECT 4.400 320.600 499.495 321.280 ;
        RECT 0.065 318.600 499.495 320.600 ;
        RECT 0.065 317.920 495.600 318.600 ;
        RECT 4.400 317.200 495.600 317.920 ;
        RECT 4.400 316.520 499.495 317.200 ;
        RECT 0.065 314.520 499.495 316.520 ;
        RECT 0.065 313.160 495.600 314.520 ;
        RECT 4.400 313.120 495.600 313.160 ;
        RECT 4.400 311.760 499.495 313.120 ;
        RECT 0.065 311.120 499.495 311.760 ;
        RECT 0.065 309.720 495.600 311.120 ;
        RECT 0.065 309.080 499.495 309.720 ;
        RECT 4.400 307.680 499.495 309.080 ;
        RECT 0.065 307.040 499.495 307.680 ;
        RECT 0.065 305.640 495.600 307.040 ;
        RECT 0.065 305.000 499.495 305.640 ;
        RECT 4.400 303.600 499.495 305.000 ;
        RECT 0.065 302.960 499.495 303.600 ;
        RECT 0.065 301.560 495.600 302.960 ;
        RECT 0.065 300.920 499.495 301.560 ;
        RECT 4.400 299.520 499.495 300.920 ;
        RECT 0.065 298.880 499.495 299.520 ;
        RECT 0.065 297.480 495.600 298.880 ;
        RECT 0.065 296.840 499.495 297.480 ;
        RECT 4.400 295.440 499.495 296.840 ;
        RECT 0.065 294.800 499.495 295.440 ;
        RECT 0.065 293.400 495.600 294.800 ;
        RECT 0.065 292.760 499.495 293.400 ;
        RECT 4.400 291.360 499.495 292.760 ;
        RECT 0.065 290.720 499.495 291.360 ;
        RECT 0.065 289.320 495.600 290.720 ;
        RECT 0.065 288.680 499.495 289.320 ;
        RECT 4.400 287.320 499.495 288.680 ;
        RECT 4.400 287.280 495.600 287.320 ;
        RECT 0.065 285.920 495.600 287.280 ;
        RECT 0.065 284.600 499.495 285.920 ;
        RECT 4.400 283.240 499.495 284.600 ;
        RECT 4.400 283.200 495.600 283.240 ;
        RECT 0.065 281.840 495.600 283.200 ;
        RECT 0.065 280.520 499.495 281.840 ;
        RECT 4.400 279.160 499.495 280.520 ;
        RECT 4.400 279.120 495.600 279.160 ;
        RECT 0.065 277.760 495.600 279.120 ;
        RECT 0.065 276.440 499.495 277.760 ;
        RECT 4.400 275.080 499.495 276.440 ;
        RECT 4.400 275.040 495.600 275.080 ;
        RECT 0.065 273.680 495.600 275.040 ;
        RECT 0.065 272.360 499.495 273.680 ;
        RECT 4.400 271.000 499.495 272.360 ;
        RECT 4.400 270.960 495.600 271.000 ;
        RECT 0.065 269.600 495.600 270.960 ;
        RECT 0.065 267.600 499.495 269.600 ;
        RECT 4.400 266.200 495.600 267.600 ;
        RECT 0.065 263.520 499.495 266.200 ;
        RECT 4.400 262.120 495.600 263.520 ;
        RECT 0.065 259.440 499.495 262.120 ;
        RECT 4.400 258.040 495.600 259.440 ;
        RECT 0.065 255.360 499.495 258.040 ;
        RECT 4.400 253.960 495.600 255.360 ;
        RECT 0.065 251.280 499.495 253.960 ;
        RECT 4.400 249.880 495.600 251.280 ;
        RECT 0.065 247.200 499.495 249.880 ;
        RECT 4.400 245.800 495.600 247.200 ;
        RECT 0.065 243.800 499.495 245.800 ;
        RECT 0.065 243.120 495.600 243.800 ;
        RECT 4.400 242.400 495.600 243.120 ;
        RECT 4.400 241.720 499.495 242.400 ;
        RECT 0.065 239.720 499.495 241.720 ;
        RECT 0.065 239.040 495.600 239.720 ;
        RECT 4.400 238.320 495.600 239.040 ;
        RECT 4.400 237.640 499.495 238.320 ;
        RECT 0.065 235.640 499.495 237.640 ;
        RECT 0.065 234.960 495.600 235.640 ;
        RECT 4.400 234.240 495.600 234.960 ;
        RECT 4.400 233.560 499.495 234.240 ;
        RECT 0.065 231.560 499.495 233.560 ;
        RECT 0.065 230.880 495.600 231.560 ;
        RECT 4.400 230.160 495.600 230.880 ;
        RECT 4.400 229.480 499.495 230.160 ;
        RECT 0.065 227.480 499.495 229.480 ;
        RECT 0.065 226.800 495.600 227.480 ;
        RECT 4.400 226.080 495.600 226.800 ;
        RECT 4.400 225.400 499.495 226.080 ;
        RECT 0.065 224.080 499.495 225.400 ;
        RECT 0.065 222.680 495.600 224.080 ;
        RECT 0.065 222.040 499.495 222.680 ;
        RECT 4.400 220.640 499.495 222.040 ;
        RECT 0.065 220.000 499.495 220.640 ;
        RECT 0.065 218.600 495.600 220.000 ;
        RECT 0.065 217.960 499.495 218.600 ;
        RECT 4.400 216.560 499.495 217.960 ;
        RECT 0.065 215.920 499.495 216.560 ;
        RECT 0.065 214.520 495.600 215.920 ;
        RECT 0.065 213.880 499.495 214.520 ;
        RECT 4.400 212.480 499.495 213.880 ;
        RECT 0.065 211.840 499.495 212.480 ;
        RECT 0.065 210.440 495.600 211.840 ;
        RECT 0.065 209.800 499.495 210.440 ;
        RECT 4.400 208.400 499.495 209.800 ;
        RECT 0.065 207.760 499.495 208.400 ;
        RECT 0.065 206.360 495.600 207.760 ;
        RECT 0.065 205.720 499.495 206.360 ;
        RECT 4.400 204.320 499.495 205.720 ;
        RECT 0.065 203.680 499.495 204.320 ;
        RECT 0.065 202.280 495.600 203.680 ;
        RECT 0.065 201.640 499.495 202.280 ;
        RECT 4.400 200.280 499.495 201.640 ;
        RECT 4.400 200.240 495.600 200.280 ;
        RECT 0.065 198.880 495.600 200.240 ;
        RECT 0.065 197.560 499.495 198.880 ;
        RECT 4.400 196.200 499.495 197.560 ;
        RECT 4.400 196.160 495.600 196.200 ;
        RECT 0.065 194.800 495.600 196.160 ;
        RECT 0.065 193.480 499.495 194.800 ;
        RECT 4.400 192.120 499.495 193.480 ;
        RECT 4.400 192.080 495.600 192.120 ;
        RECT 0.065 190.720 495.600 192.080 ;
        RECT 0.065 189.400 499.495 190.720 ;
        RECT 4.400 188.040 499.495 189.400 ;
        RECT 4.400 188.000 495.600 188.040 ;
        RECT 0.065 186.640 495.600 188.000 ;
        RECT 0.065 185.320 499.495 186.640 ;
        RECT 4.400 183.960 499.495 185.320 ;
        RECT 4.400 183.920 495.600 183.960 ;
        RECT 0.065 182.560 495.600 183.920 ;
        RECT 0.065 181.240 499.495 182.560 ;
        RECT 4.400 179.880 499.495 181.240 ;
        RECT 4.400 179.840 495.600 179.880 ;
        RECT 0.065 178.480 495.600 179.840 ;
        RECT 0.065 176.480 499.495 178.480 ;
        RECT 4.400 175.080 495.600 176.480 ;
        RECT 0.065 172.400 499.495 175.080 ;
        RECT 4.400 171.000 495.600 172.400 ;
        RECT 0.065 168.320 499.495 171.000 ;
        RECT 4.400 166.920 495.600 168.320 ;
        RECT 0.065 164.240 499.495 166.920 ;
        RECT 4.400 162.840 495.600 164.240 ;
        RECT 0.065 160.160 499.495 162.840 ;
        RECT 4.400 158.760 495.600 160.160 ;
        RECT 0.065 156.760 499.495 158.760 ;
        RECT 0.065 156.080 495.600 156.760 ;
        RECT 4.400 155.360 495.600 156.080 ;
        RECT 4.400 154.680 499.495 155.360 ;
        RECT 0.065 152.680 499.495 154.680 ;
        RECT 0.065 152.000 495.600 152.680 ;
        RECT 4.400 151.280 495.600 152.000 ;
        RECT 4.400 150.600 499.495 151.280 ;
        RECT 0.065 148.600 499.495 150.600 ;
        RECT 0.065 147.920 495.600 148.600 ;
        RECT 4.400 147.200 495.600 147.920 ;
        RECT 4.400 146.520 499.495 147.200 ;
        RECT 0.065 144.520 499.495 146.520 ;
        RECT 0.065 143.840 495.600 144.520 ;
        RECT 4.400 143.120 495.600 143.840 ;
        RECT 4.400 142.440 499.495 143.120 ;
        RECT 0.065 140.440 499.495 142.440 ;
        RECT 0.065 139.760 495.600 140.440 ;
        RECT 4.400 139.040 495.600 139.760 ;
        RECT 4.400 138.360 499.495 139.040 ;
        RECT 0.065 136.360 499.495 138.360 ;
        RECT 0.065 135.000 495.600 136.360 ;
        RECT 4.400 134.960 495.600 135.000 ;
        RECT 4.400 133.600 499.495 134.960 ;
        RECT 0.065 132.960 499.495 133.600 ;
        RECT 0.065 131.560 495.600 132.960 ;
        RECT 0.065 130.920 499.495 131.560 ;
        RECT 4.400 129.520 499.495 130.920 ;
        RECT 0.065 128.880 499.495 129.520 ;
        RECT 0.065 127.480 495.600 128.880 ;
        RECT 0.065 126.840 499.495 127.480 ;
        RECT 4.400 125.440 499.495 126.840 ;
        RECT 0.065 124.800 499.495 125.440 ;
        RECT 0.065 123.400 495.600 124.800 ;
        RECT 0.065 122.760 499.495 123.400 ;
        RECT 4.400 121.360 499.495 122.760 ;
        RECT 0.065 120.720 499.495 121.360 ;
        RECT 0.065 119.320 495.600 120.720 ;
        RECT 0.065 118.680 499.495 119.320 ;
        RECT 4.400 117.280 499.495 118.680 ;
        RECT 0.065 116.640 499.495 117.280 ;
        RECT 0.065 115.240 495.600 116.640 ;
        RECT 0.065 114.600 499.495 115.240 ;
        RECT 4.400 113.240 499.495 114.600 ;
        RECT 4.400 113.200 495.600 113.240 ;
        RECT 0.065 111.840 495.600 113.200 ;
        RECT 0.065 110.520 499.495 111.840 ;
        RECT 4.400 109.160 499.495 110.520 ;
        RECT 4.400 109.120 495.600 109.160 ;
        RECT 0.065 107.760 495.600 109.120 ;
        RECT 0.065 106.440 499.495 107.760 ;
        RECT 4.400 105.080 499.495 106.440 ;
        RECT 4.400 105.040 495.600 105.080 ;
        RECT 0.065 103.680 495.600 105.040 ;
        RECT 0.065 102.360 499.495 103.680 ;
        RECT 4.400 101.000 499.495 102.360 ;
        RECT 4.400 100.960 495.600 101.000 ;
        RECT 0.065 99.600 495.600 100.960 ;
        RECT 0.065 98.280 499.495 99.600 ;
        RECT 4.400 96.920 499.495 98.280 ;
        RECT 4.400 96.880 495.600 96.920 ;
        RECT 0.065 95.520 495.600 96.880 ;
        RECT 0.065 94.200 499.495 95.520 ;
        RECT 4.400 92.840 499.495 94.200 ;
        RECT 4.400 92.800 495.600 92.840 ;
        RECT 0.065 91.440 495.600 92.800 ;
        RECT 0.065 89.440 499.495 91.440 ;
        RECT 4.400 88.040 495.600 89.440 ;
        RECT 0.065 85.360 499.495 88.040 ;
        RECT 4.400 83.960 495.600 85.360 ;
        RECT 0.065 81.280 499.495 83.960 ;
        RECT 4.400 79.880 495.600 81.280 ;
        RECT 0.065 77.200 499.495 79.880 ;
        RECT 4.400 75.800 495.600 77.200 ;
        RECT 0.065 73.120 499.495 75.800 ;
        RECT 4.400 71.720 495.600 73.120 ;
        RECT 0.065 69.040 499.495 71.720 ;
        RECT 4.400 67.640 495.600 69.040 ;
        RECT 0.065 65.640 499.495 67.640 ;
        RECT 0.065 64.960 495.600 65.640 ;
        RECT 4.400 64.240 495.600 64.960 ;
        RECT 4.400 63.560 499.495 64.240 ;
        RECT 0.065 61.560 499.495 63.560 ;
        RECT 0.065 60.880 495.600 61.560 ;
        RECT 4.400 60.160 495.600 60.880 ;
        RECT 4.400 59.480 499.495 60.160 ;
        RECT 0.065 57.480 499.495 59.480 ;
        RECT 0.065 56.800 495.600 57.480 ;
        RECT 4.400 56.080 495.600 56.800 ;
        RECT 4.400 55.400 499.495 56.080 ;
        RECT 0.065 53.400 499.495 55.400 ;
        RECT 0.065 52.720 495.600 53.400 ;
        RECT 4.400 52.000 495.600 52.720 ;
        RECT 4.400 51.320 499.495 52.000 ;
        RECT 0.065 49.320 499.495 51.320 ;
        RECT 0.065 48.640 495.600 49.320 ;
        RECT 4.400 47.920 495.600 48.640 ;
        RECT 4.400 47.240 499.495 47.920 ;
        RECT 0.065 45.920 499.495 47.240 ;
        RECT 0.065 44.520 495.600 45.920 ;
        RECT 0.065 43.880 499.495 44.520 ;
        RECT 4.400 42.480 499.495 43.880 ;
        RECT 0.065 41.840 499.495 42.480 ;
        RECT 0.065 40.440 495.600 41.840 ;
        RECT 0.065 39.800 499.495 40.440 ;
        RECT 4.400 38.400 499.495 39.800 ;
        RECT 0.065 37.760 499.495 38.400 ;
        RECT 0.065 36.360 495.600 37.760 ;
        RECT 0.065 35.720 499.495 36.360 ;
        RECT 4.400 34.320 499.495 35.720 ;
        RECT 0.065 33.680 499.495 34.320 ;
        RECT 0.065 32.280 495.600 33.680 ;
        RECT 0.065 31.640 499.495 32.280 ;
        RECT 4.400 30.240 499.495 31.640 ;
        RECT 0.065 29.600 499.495 30.240 ;
        RECT 0.065 28.200 495.600 29.600 ;
        RECT 0.065 27.560 499.495 28.200 ;
        RECT 4.400 26.160 499.495 27.560 ;
        RECT 0.065 25.520 499.495 26.160 ;
        RECT 0.065 24.120 495.600 25.520 ;
        RECT 0.065 23.480 499.495 24.120 ;
        RECT 4.400 22.120 499.495 23.480 ;
        RECT 4.400 22.080 495.600 22.120 ;
        RECT 0.065 20.720 495.600 22.080 ;
        RECT 0.065 19.400 499.495 20.720 ;
        RECT 4.400 18.040 499.495 19.400 ;
        RECT 4.400 18.000 495.600 18.040 ;
        RECT 0.065 16.640 495.600 18.000 ;
        RECT 0.065 15.320 499.495 16.640 ;
        RECT 4.400 13.960 499.495 15.320 ;
        RECT 4.400 13.920 495.600 13.960 ;
        RECT 0.065 12.560 495.600 13.920 ;
        RECT 0.065 11.240 499.495 12.560 ;
        RECT 4.400 9.880 499.495 11.240 ;
        RECT 4.400 9.840 495.600 9.880 ;
        RECT 0.065 8.480 495.600 9.840 ;
        RECT 0.065 7.160 499.495 8.480 ;
        RECT 4.400 5.800 499.495 7.160 ;
        RECT 4.400 5.760 495.600 5.800 ;
        RECT 0.065 4.400 495.600 5.760 ;
        RECT 0.065 3.080 499.495 4.400 ;
        RECT 4.400 2.400 499.495 3.080 ;
        RECT 4.400 1.680 495.600 2.400 ;
        RECT 0.065 1.535 495.600 1.680 ;
      LAYER met4 ;
        RECT 10.415 23.975 20.640 775.705 ;
        RECT 23.040 23.975 97.440 775.705 ;
        RECT 99.840 23.975 174.240 775.705 ;
        RECT 176.640 23.975 251.040 775.705 ;
        RECT 253.440 23.975 327.840 775.705 ;
        RECT 330.240 23.975 404.640 775.705 ;
        RECT 407.040 23.975 481.440 775.705 ;
        RECT 483.840 23.975 495.585 775.705 ;
  END
END ExperiarCore
END LIBRARY

