VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ExperiarCore
  CLASS BLOCK ;
  FOREIGN ExperiarCore ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 900.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END addr0[8]
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.760 4.000 564.360 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 577.360 4.000 577.960 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.880 4.000 587.480 ;
    END
  END addr1[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END clk0
  PIN clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END clk1
  PIN coreIndex[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 896.000 5.430 900.000 ;
    END
  END coreIndex[0]
  PIN coreIndex[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 896.000 16.010 900.000 ;
    END
  END coreIndex[1]
  PIN coreIndex[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 896.000 26.590 900.000 ;
    END
  END coreIndex[2]
  PIN coreIndex[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 896.000 37.170 900.000 ;
    END
  END coreIndex[3]
  PIN coreIndex[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 896.000 48.210 900.000 ;
    END
  END coreIndex[4]
  PIN coreIndex[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 896.000 58.790 900.000 ;
    END
  END coreIndex[5]
  PIN coreIndex[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 896.000 69.370 900.000 ;
    END
  END coreIndex[6]
  PIN coreIndex[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 896.000 80.410 900.000 ;
    END
  END coreIndex[7]
  PIN core_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 10.240 450.000 10.840 ;
    END
  END core_wb_ack_i
  PIN core_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 36.760 450.000 37.360 ;
    END
  END core_wb_adr_o[0]
  PIN core_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 185.000 450.000 185.600 ;
    END
  END core_wb_adr_o[10]
  PIN core_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 198.600 450.000 199.200 ;
    END
  END core_wb_adr_o[11]
  PIN core_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 211.520 450.000 212.120 ;
    END
  END core_wb_adr_o[12]
  PIN core_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 224.440 450.000 225.040 ;
    END
  END core_wb_adr_o[13]
  PIN core_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 238.040 450.000 238.640 ;
    END
  END core_wb_adr_o[14]
  PIN core_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 250.960 450.000 251.560 ;
    END
  END core_wb_adr_o[15]
  PIN core_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 263.880 450.000 264.480 ;
    END
  END core_wb_adr_o[16]
  PIN core_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 276.800 450.000 277.400 ;
    END
  END core_wb_adr_o[17]
  PIN core_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 290.400 450.000 291.000 ;
    END
  END core_wb_adr_o[18]
  PIN core_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 303.320 450.000 303.920 ;
    END
  END core_wb_adr_o[19]
  PIN core_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 54.440 450.000 55.040 ;
    END
  END core_wb_adr_o[1]
  PIN core_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 316.240 450.000 316.840 ;
    END
  END core_wb_adr_o[20]
  PIN core_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 329.840 450.000 330.440 ;
    END
  END core_wb_adr_o[21]
  PIN core_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 342.760 450.000 343.360 ;
    END
  END core_wb_adr_o[22]
  PIN core_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 355.680 450.000 356.280 ;
    END
  END core_wb_adr_o[23]
  PIN core_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 368.600 450.000 369.200 ;
    END
  END core_wb_adr_o[24]
  PIN core_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 382.200 450.000 382.800 ;
    END
  END core_wb_adr_o[25]
  PIN core_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 395.120 450.000 395.720 ;
    END
  END core_wb_adr_o[26]
  PIN core_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 408.040 450.000 408.640 ;
    END
  END core_wb_adr_o[27]
  PIN core_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 71.440 450.000 72.040 ;
    END
  END core_wb_adr_o[2]
  PIN core_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 89.120 450.000 89.720 ;
    END
  END core_wb_adr_o[3]
  PIN core_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 106.800 450.000 107.400 ;
    END
  END core_wb_adr_o[4]
  PIN core_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 119.720 450.000 120.320 ;
    END
  END core_wb_adr_o[5]
  PIN core_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 132.640 450.000 133.240 ;
    END
  END core_wb_adr_o[6]
  PIN core_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 146.240 450.000 146.840 ;
    END
  END core_wb_adr_o[7]
  PIN core_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 159.160 450.000 159.760 ;
    END
  END core_wb_adr_o[8]
  PIN core_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 172.080 450.000 172.680 ;
    END
  END core_wb_adr_o[9]
  PIN core_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 15.000 450.000 15.600 ;
    END
  END core_wb_cyc_o
  PIN core_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 40.840 450.000 41.440 ;
    END
  END core_wb_data_i[0]
  PIN core_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 189.760 450.000 190.360 ;
    END
  END core_wb_data_i[10]
  PIN core_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 202.680 450.000 203.280 ;
    END
  END core_wb_data_i[11]
  PIN core_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 215.600 450.000 216.200 ;
    END
  END core_wb_data_i[12]
  PIN core_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 229.200 450.000 229.800 ;
    END
  END core_wb_data_i[13]
  PIN core_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 242.120 450.000 242.720 ;
    END
  END core_wb_data_i[14]
  PIN core_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 255.040 450.000 255.640 ;
    END
  END core_wb_data_i[15]
  PIN core_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 268.640 450.000 269.240 ;
    END
  END core_wb_data_i[16]
  PIN core_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 281.560 450.000 282.160 ;
    END
  END core_wb_data_i[17]
  PIN core_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 294.480 450.000 295.080 ;
    END
  END core_wb_data_i[18]
  PIN core_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 307.400 450.000 308.000 ;
    END
  END core_wb_data_i[19]
  PIN core_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 58.520 450.000 59.120 ;
    END
  END core_wb_data_i[1]
  PIN core_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 321.000 450.000 321.600 ;
    END
  END core_wb_data_i[20]
  PIN core_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 333.920 450.000 334.520 ;
    END
  END core_wb_data_i[21]
  PIN core_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 346.840 450.000 347.440 ;
    END
  END core_wb_data_i[22]
  PIN core_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 360.440 450.000 361.040 ;
    END
  END core_wb_data_i[23]
  PIN core_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 373.360 450.000 373.960 ;
    END
  END core_wb_data_i[24]
  PIN core_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 386.280 450.000 386.880 ;
    END
  END core_wb_data_i[25]
  PIN core_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 399.200 450.000 399.800 ;
    END
  END core_wb_data_i[26]
  PIN core_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 412.800 450.000 413.400 ;
    END
  END core_wb_data_i[27]
  PIN core_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 421.640 450.000 422.240 ;
    END
  END core_wb_data_i[28]
  PIN core_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 429.800 450.000 430.400 ;
    END
  END core_wb_data_i[29]
  PIN core_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 76.200 450.000 76.800 ;
    END
  END core_wb_data_i[2]
  PIN core_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 438.640 450.000 439.240 ;
    END
  END core_wb_data_i[30]
  PIN core_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 447.480 450.000 448.080 ;
    END
  END core_wb_data_i[31]
  PIN core_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 93.200 450.000 93.800 ;
    END
  END core_wb_data_i[3]
  PIN core_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 110.880 450.000 111.480 ;
    END
  END core_wb_data_i[4]
  PIN core_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 123.800 450.000 124.400 ;
    END
  END core_wb_data_i[5]
  PIN core_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 137.400 450.000 138.000 ;
    END
  END core_wb_data_i[6]
  PIN core_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 150.320 450.000 150.920 ;
    END
  END core_wb_data_i[7]
  PIN core_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 163.240 450.000 163.840 ;
    END
  END core_wb_data_i[8]
  PIN core_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 176.840 450.000 177.440 ;
    END
  END core_wb_data_i[9]
  PIN core_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 45.600 450.000 46.200 ;
    END
  END core_wb_data_o[0]
  PIN core_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 193.840 450.000 194.440 ;
    END
  END core_wb_data_o[10]
  PIN core_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 207.440 450.000 208.040 ;
    END
  END core_wb_data_o[11]
  PIN core_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 220.360 450.000 220.960 ;
    END
  END core_wb_data_o[12]
  PIN core_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 233.280 450.000 233.880 ;
    END
  END core_wb_data_o[13]
  PIN core_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 246.200 450.000 246.800 ;
    END
  END core_wb_data_o[14]
  PIN core_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 259.800 450.000 260.400 ;
    END
  END core_wb_data_o[15]
  PIN core_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 272.720 450.000 273.320 ;
    END
  END core_wb_data_o[16]
  PIN core_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 285.640 450.000 286.240 ;
    END
  END core_wb_data_o[17]
  PIN core_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 299.240 450.000 299.840 ;
    END
  END core_wb_data_o[18]
  PIN core_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 312.160 450.000 312.760 ;
    END
  END core_wb_data_o[19]
  PIN core_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 62.600 450.000 63.200 ;
    END
  END core_wb_data_o[1]
  PIN core_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 325.080 450.000 325.680 ;
    END
  END core_wb_data_o[20]
  PIN core_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 338.000 450.000 338.600 ;
    END
  END core_wb_data_o[21]
  PIN core_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 351.600 450.000 352.200 ;
    END
  END core_wb_data_o[22]
  PIN core_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 364.520 450.000 365.120 ;
    END
  END core_wb_data_o[23]
  PIN core_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 377.440 450.000 378.040 ;
    END
  END core_wb_data_o[24]
  PIN core_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 391.040 450.000 391.640 ;
    END
  END core_wb_data_o[25]
  PIN core_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 403.960 450.000 404.560 ;
    END
  END core_wb_data_o[26]
  PIN core_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 416.880 450.000 417.480 ;
    END
  END core_wb_data_o[27]
  PIN core_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 425.720 450.000 426.320 ;
    END
  END core_wb_data_o[28]
  PIN core_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 434.560 450.000 435.160 ;
    END
  END core_wb_data_o[29]
  PIN core_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 80.280 450.000 80.880 ;
    END
  END core_wb_data_o[2]
  PIN core_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 443.400 450.000 444.000 ;
    END
  END core_wb_data_o[30]
  PIN core_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 452.240 450.000 452.840 ;
    END
  END core_wb_data_o[31]
  PIN core_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 97.960 450.000 98.560 ;
    END
  END core_wb_data_o[3]
  PIN core_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 115.640 450.000 116.240 ;
    END
  END core_wb_data_o[4]
  PIN core_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 128.560 450.000 129.160 ;
    END
  END core_wb_data_o[5]
  PIN core_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 141.480 450.000 142.080 ;
    END
  END core_wb_data_o[6]
  PIN core_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 154.400 450.000 155.000 ;
    END
  END core_wb_data_o[7]
  PIN core_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 168.000 450.000 168.600 ;
    END
  END core_wb_data_o[8]
  PIN core_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 180.920 450.000 181.520 ;
    END
  END core_wb_data_o[9]
  PIN core_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 19.080 450.000 19.680 ;
    END
  END core_wb_error_i
  PIN core_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 49.680 450.000 50.280 ;
    END
  END core_wb_sel_o[0]
  PIN core_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 67.360 450.000 67.960 ;
    END
  END core_wb_sel_o[1]
  PIN core_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 85.040 450.000 85.640 ;
    END
  END core_wb_sel_o[2]
  PIN core_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 102.040 450.000 102.640 ;
    END
  END core_wb_sel_o[3]
  PIN core_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 23.840 450.000 24.440 ;
    END
  END core_wb_stall_i
  PIN core_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 27.920 450.000 28.520 ;
    END
  END core_wb_stb_o
  PIN core_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 32.000 450.000 32.600 ;
    END
  END core_wb_we_o
  PIN csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END csb0[0]
  PIN csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END csb0[1]
  PIN csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END csb1[0]
  PIN csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END csb1[1]
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END din0[9]
  PIN dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.000 4.000 372.600 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END dout0[32]
  PIN dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END dout0[33]
  PIN dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END dout0[34]
  PIN dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END dout0[35]
  PIN dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END dout0[36]
  PIN dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END dout0[37]
  PIN dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END dout0[38]
  PIN dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 422.320 4.000 422.920 ;
    END
  END dout0[39]
  PIN dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END dout0[3]
  PIN dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END dout0[40]
  PIN dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END dout0[41]
  PIN dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END dout0[42]
  PIN dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END dout0[43]
  PIN dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END dout0[44]
  PIN dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END dout0[45]
  PIN dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END dout0[46]
  PIN dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END dout0[47]
  PIN dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END dout0[48]
  PIN dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END dout0[49]
  PIN dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END dout0[4]
  PIN dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END dout0[50]
  PIN dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END dout0[51]
  PIN dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END dout0[52]
  PIN dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END dout0[53]
  PIN dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END dout0[54]
  PIN dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END dout0[55]
  PIN dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END dout0[56]
  PIN dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END dout0[57]
  PIN dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 509.360 4.000 509.960 ;
    END
  END dout0[58]
  PIN dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END dout0[59]
  PIN dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END dout0[5]
  PIN dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END dout0[60]
  PIN dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.960 4.000 523.560 ;
    END
  END dout0[61]
  PIN dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END dout0[62]
  PIN dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END dout0[63]
  PIN dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.200 4.000 637.800 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.280 4.000 641.880 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 687.520 4.000 688.120 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.120 4.000 701.720 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.720 4.000 715.320 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 723.560 4.000 724.160 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 600.480 4.000 601.080 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 728.320 4.000 728.920 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END dout1[31]
  PIN dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END dout1[32]
  PIN dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.920 4.000 742.520 ;
    END
  END dout1[33]
  PIN dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END dout1[34]
  PIN dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END dout1[35]
  PIN dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END dout1[36]
  PIN dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END dout1[37]
  PIN dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END dout1[38]
  PIN dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END dout1[39]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END dout1[3]
  PIN dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.880 4.000 774.480 ;
    END
  END dout1[40]
  PIN dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END dout1[41]
  PIN dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 783.400 4.000 784.000 ;
    END
  END dout1[42]
  PIN dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END dout1[43]
  PIN dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END dout1[44]
  PIN dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END dout1[45]
  PIN dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.760 4.000 802.360 ;
    END
  END dout1[46]
  PIN dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END dout1[47]
  PIN dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END dout1[48]
  PIN dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END dout1[49]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END dout1[4]
  PIN dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END dout1[50]
  PIN dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.200 4.000 824.800 ;
    END
  END dout1[51]
  PIN dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.960 4.000 829.560 ;
    END
  END dout1[52]
  PIN dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.720 4.000 834.320 ;
    END
  END dout1[53]
  PIN dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END dout1[54]
  PIN dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 842.560 4.000 843.160 ;
    END
  END dout1[55]
  PIN dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 847.320 4.000 847.920 ;
    END
  END dout1[56]
  PIN dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 852.080 4.000 852.680 ;
    END
  END dout1[57]
  PIN dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.160 4.000 856.760 ;
    END
  END dout1[58]
  PIN dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.920 4.000 861.520 ;
    END
  END dout1[59]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.080 4.000 614.680 ;
    END
  END dout1[5]
  PIN dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.680 4.000 866.280 ;
    END
  END dout1[60]
  PIN dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 869.760 4.000 870.360 ;
    END
  END dout1[61]
  PIN dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 874.520 4.000 875.120 ;
    END
  END dout1[62]
  PIN dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.280 4.000 879.880 ;
    END
  END dout1[63]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END dout1[9]
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END irq[0]
  PIN irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 888.800 450.000 889.400 ;
    END
  END irq[10]
  PIN irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 896.000 444.270 900.000 ;
    END
  END irq[11]
  PIN irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 893.560 450.000 894.160 ;
    END
  END irq[12]
  PIN irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END irq[13]
  PIN irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END irq[14]
  PIN irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 897.640 450.000 898.240 ;
    END
  END irq[15]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 896.000 423.110 900.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 884.720 450.000 885.320 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 896.000 433.690 900.000 ;
    END
  END irq[5]
  PIN irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END irq[6]
  PIN irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END irq[7]
  PIN irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END irq[8]
  PIN irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.880 4.000 893.480 ;
    END
  END irq[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END jtag_tms
  PIN localMemory_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 456.320 450.000 456.920 ;
    END
  END localMemory_wb_ack_o
  PIN localMemory_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 482.160 450.000 482.760 ;
    END
  END localMemory_wb_adr_i[0]
  PIN localMemory_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 631.080 450.000 631.680 ;
    END
  END localMemory_wb_adr_i[10]
  PIN localMemory_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 644.000 450.000 644.600 ;
    END
  END localMemory_wb_adr_i[11]
  PIN localMemory_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 657.600 450.000 658.200 ;
    END
  END localMemory_wb_adr_i[12]
  PIN localMemory_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 670.520 450.000 671.120 ;
    END
  END localMemory_wb_adr_i[13]
  PIN localMemory_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 683.440 450.000 684.040 ;
    END
  END localMemory_wb_adr_i[14]
  PIN localMemory_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 696.360 450.000 696.960 ;
    END
  END localMemory_wb_adr_i[15]
  PIN localMemory_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 709.960 450.000 710.560 ;
    END
  END localMemory_wb_adr_i[16]
  PIN localMemory_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 722.880 450.000 723.480 ;
    END
  END localMemory_wb_adr_i[17]
  PIN localMemory_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 735.800 450.000 736.400 ;
    END
  END localMemory_wb_adr_i[18]
  PIN localMemory_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 749.400 450.000 750.000 ;
    END
  END localMemory_wb_adr_i[19]
  PIN localMemory_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 499.840 450.000 500.440 ;
    END
  END localMemory_wb_adr_i[1]
  PIN localMemory_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 762.320 450.000 762.920 ;
    END
  END localMemory_wb_adr_i[20]
  PIN localMemory_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 775.240 450.000 775.840 ;
    END
  END localMemory_wb_adr_i[21]
  PIN localMemory_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 788.160 450.000 788.760 ;
    END
  END localMemory_wb_adr_i[22]
  PIN localMemory_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 801.760 450.000 802.360 ;
    END
  END localMemory_wb_adr_i[23]
  PIN localMemory_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 517.520 450.000 518.120 ;
    END
  END localMemory_wb_adr_i[2]
  PIN localMemory_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 535.200 450.000 535.800 ;
    END
  END localMemory_wb_adr_i[3]
  PIN localMemory_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 552.200 450.000 552.800 ;
    END
  END localMemory_wb_adr_i[4]
  PIN localMemory_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 565.800 450.000 566.400 ;
    END
  END localMemory_wb_adr_i[5]
  PIN localMemory_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 578.720 450.000 579.320 ;
    END
  END localMemory_wb_adr_i[6]
  PIN localMemory_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 591.640 450.000 592.240 ;
    END
  END localMemory_wb_adr_i[7]
  PIN localMemory_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 604.560 450.000 605.160 ;
    END
  END localMemory_wb_adr_i[8]
  PIN localMemory_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 618.160 450.000 618.760 ;
    END
  END localMemory_wb_adr_i[9]
  PIN localMemory_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 460.400 450.000 461.000 ;
    END
  END localMemory_wb_cyc_i
  PIN localMemory_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 486.920 450.000 487.520 ;
    END
  END localMemory_wb_data_i[0]
  PIN localMemory_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 635.160 450.000 635.760 ;
    END
  END localMemory_wb_data_i[10]
  PIN localMemory_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 648.760 450.000 649.360 ;
    END
  END localMemory_wb_data_i[11]
  PIN localMemory_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 661.680 450.000 662.280 ;
    END
  END localMemory_wb_data_i[12]
  PIN localMemory_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 674.600 450.000 675.200 ;
    END
  END localMemory_wb_data_i[13]
  PIN localMemory_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 688.200 450.000 688.800 ;
    END
  END localMemory_wb_data_i[14]
  PIN localMemory_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 701.120 450.000 701.720 ;
    END
  END localMemory_wb_data_i[15]
  PIN localMemory_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 714.040 450.000 714.640 ;
    END
  END localMemory_wb_data_i[16]
  PIN localMemory_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 726.960 450.000 727.560 ;
    END
  END localMemory_wb_data_i[17]
  PIN localMemory_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 740.560 450.000 741.160 ;
    END
  END localMemory_wb_data_i[18]
  PIN localMemory_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 753.480 450.000 754.080 ;
    END
  END localMemory_wb_data_i[19]
  PIN localMemory_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 504.600 450.000 505.200 ;
    END
  END localMemory_wb_data_i[1]
  PIN localMemory_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 766.400 450.000 767.000 ;
    END
  END localMemory_wb_data_i[20]
  PIN localMemory_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 780.000 450.000 780.600 ;
    END
  END localMemory_wb_data_i[21]
  PIN localMemory_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 792.920 450.000 793.520 ;
    END
  END localMemory_wb_data_i[22]
  PIN localMemory_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 805.840 450.000 806.440 ;
    END
  END localMemory_wb_data_i[23]
  PIN localMemory_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 814.680 450.000 815.280 ;
    END
  END localMemory_wb_data_i[24]
  PIN localMemory_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 823.520 450.000 824.120 ;
    END
  END localMemory_wb_data_i[25]
  PIN localMemory_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 832.360 450.000 832.960 ;
    END
  END localMemory_wb_data_i[26]
  PIN localMemory_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 841.200 450.000 841.800 ;
    END
  END localMemory_wb_data_i[27]
  PIN localMemory_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 849.360 450.000 849.960 ;
    END
  END localMemory_wb_data_i[28]
  PIN localMemory_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 858.200 450.000 858.800 ;
    END
  END localMemory_wb_data_i[29]
  PIN localMemory_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 521.600 450.000 522.200 ;
    END
  END localMemory_wb_data_i[2]
  PIN localMemory_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 867.040 450.000 867.640 ;
    END
  END localMemory_wb_data_i[30]
  PIN localMemory_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 875.880 450.000 876.480 ;
    END
  END localMemory_wb_data_i[31]
  PIN localMemory_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 539.280 450.000 539.880 ;
    END
  END localMemory_wb_data_i[3]
  PIN localMemory_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 556.960 450.000 557.560 ;
    END
  END localMemory_wb_data_i[4]
  PIN localMemory_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 569.880 450.000 570.480 ;
    END
  END localMemory_wb_data_i[5]
  PIN localMemory_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 582.800 450.000 583.400 ;
    END
  END localMemory_wb_data_i[6]
  PIN localMemory_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 596.400 450.000 597.000 ;
    END
  END localMemory_wb_data_i[7]
  PIN localMemory_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 609.320 450.000 609.920 ;
    END
  END localMemory_wb_data_i[8]
  PIN localMemory_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 622.240 450.000 622.840 ;
    END
  END localMemory_wb_data_i[9]
  PIN localMemory_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 491.000 450.000 491.600 ;
    END
  END localMemory_wb_data_o[0]
  PIN localMemory_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 639.920 450.000 640.520 ;
    END
  END localMemory_wb_data_o[10]
  PIN localMemory_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 652.840 450.000 653.440 ;
    END
  END localMemory_wb_data_o[11]
  PIN localMemory_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 665.760 450.000 666.360 ;
    END
  END localMemory_wb_data_o[12]
  PIN localMemory_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 679.360 450.000 679.960 ;
    END
  END localMemory_wb_data_o[13]
  PIN localMemory_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 692.280 450.000 692.880 ;
    END
  END localMemory_wb_data_o[14]
  PIN localMemory_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 705.200 450.000 705.800 ;
    END
  END localMemory_wb_data_o[15]
  PIN localMemory_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 718.800 450.000 719.400 ;
    END
  END localMemory_wb_data_o[16]
  PIN localMemory_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 731.720 450.000 732.320 ;
    END
  END localMemory_wb_data_o[17]
  PIN localMemory_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 744.640 450.000 745.240 ;
    END
  END localMemory_wb_data_o[18]
  PIN localMemory_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 757.560 450.000 758.160 ;
    END
  END localMemory_wb_data_o[19]
  PIN localMemory_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 508.680 450.000 509.280 ;
    END
  END localMemory_wb_data_o[1]
  PIN localMemory_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 771.160 450.000 771.760 ;
    END
  END localMemory_wb_data_o[20]
  PIN localMemory_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 784.080 450.000 784.680 ;
    END
  END localMemory_wb_data_o[21]
  PIN localMemory_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 797.000 450.000 797.600 ;
    END
  END localMemory_wb_data_o[22]
  PIN localMemory_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 810.600 450.000 811.200 ;
    END
  END localMemory_wb_data_o[23]
  PIN localMemory_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 818.760 450.000 819.360 ;
    END
  END localMemory_wb_data_o[24]
  PIN localMemory_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 827.600 450.000 828.200 ;
    END
  END localMemory_wb_data_o[25]
  PIN localMemory_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 836.440 450.000 837.040 ;
    END
  END localMemory_wb_data_o[26]
  PIN localMemory_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 845.280 450.000 845.880 ;
    END
  END localMemory_wb_data_o[27]
  PIN localMemory_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 854.120 450.000 854.720 ;
    END
  END localMemory_wb_data_o[28]
  PIN localMemory_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 862.960 450.000 863.560 ;
    END
  END localMemory_wb_data_o[29]
  PIN localMemory_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 526.360 450.000 526.960 ;
    END
  END localMemory_wb_data_o[2]
  PIN localMemory_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 871.800 450.000 872.400 ;
    END
  END localMemory_wb_data_o[30]
  PIN localMemory_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 879.960 450.000 880.560 ;
    END
  END localMemory_wb_data_o[31]
  PIN localMemory_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 543.360 450.000 543.960 ;
    END
  END localMemory_wb_data_o[3]
  PIN localMemory_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 561.040 450.000 561.640 ;
    END
  END localMemory_wb_data_o[4]
  PIN localMemory_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 573.960 450.000 574.560 ;
    END
  END localMemory_wb_data_o[5]
  PIN localMemory_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 587.560 450.000 588.160 ;
    END
  END localMemory_wb_data_o[6]
  PIN localMemory_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 600.480 450.000 601.080 ;
    END
  END localMemory_wb_data_o[7]
  PIN localMemory_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 613.400 450.000 614.000 ;
    END
  END localMemory_wb_data_o[8]
  PIN localMemory_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 627.000 450.000 627.600 ;
    END
  END localMemory_wb_data_o[9]
  PIN localMemory_wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 465.160 450.000 465.760 ;
    END
  END localMemory_wb_error_o
  PIN localMemory_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 495.760 450.000 496.360 ;
    END
  END localMemory_wb_sel_i[0]
  PIN localMemory_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 512.760 450.000 513.360 ;
    END
  END localMemory_wb_sel_i[1]
  PIN localMemory_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 530.440 450.000 531.040 ;
    END
  END localMemory_wb_sel_i[2]
  PIN localMemory_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 548.120 450.000 548.720 ;
    END
  END localMemory_wb_sel_i[3]
  PIN localMemory_wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 469.240 450.000 469.840 ;
    END
  END localMemory_wb_stall_o
  PIN localMemory_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 474.000 450.000 474.600 ;
    END
  END localMemory_wb_stb_i
  PIN localMemory_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 478.080 450.000 478.680 ;
    END
  END localMemory_wb_we_i
  PIN manufacturerID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 896.000 90.990 900.000 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 896.000 198.170 900.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 896.000 101.570 900.000 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 896.000 112.150 900.000 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 896.000 123.190 900.000 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 896.000 133.770 900.000 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 896.000 144.350 900.000 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 896.000 155.390 900.000 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 896.000 165.970 900.000 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 896.000 176.550 900.000 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 896.000 187.130 900.000 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 896.000 208.750 900.000 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 896.000 315.930 900.000 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 896.000 326.510 900.000 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 896.000 337.090 900.000 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 896.000 348.130 900.000 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 896.000 358.710 900.000 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 896.000 369.290 900.000 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 896.000 219.330 900.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 896.000 230.370 900.000 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 896.000 240.950 900.000 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 896.000 251.530 900.000 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 896.000 262.110 900.000 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 896.000 273.150 900.000 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 896.000 283.730 900.000 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 896.000 294.310 900.000 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 896.000 305.350 900.000 ;
    END
  END partID[9]
  PIN probe_env[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END probe_env[0]
  PIN probe_env[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END probe_env[1]
  PIN probe_errorCode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END probe_errorCode[0]
  PIN probe_errorCode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END probe_errorCode[1]
  PIN probe_isBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END probe_isBranch
  PIN probe_isCompressed
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END probe_isCompressed
  PIN probe_isLoad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END probe_isLoad
  PIN probe_isStore
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END probe_isStore
  PIN probe_jtagInstruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END probe_jtagInstruction[0]
  PIN probe_jtagInstruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END probe_jtagInstruction[1]
  PIN probe_jtagInstruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END probe_jtagInstruction[2]
  PIN probe_jtagInstruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END probe_jtagInstruction[3]
  PIN probe_jtagInstruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END probe_jtagInstruction[4]
  PIN probe_opcode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END probe_opcode[0]
  PIN probe_opcode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END probe_opcode[1]
  PIN probe_opcode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END probe_opcode[2]
  PIN probe_opcode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END probe_opcode[3]
  PIN probe_opcode[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END probe_opcode[4]
  PIN probe_opcode[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END probe_opcode[5]
  PIN probe_opcode[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END probe_opcode[6]
  PIN probe_programCounter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END probe_programCounter[0]
  PIN probe_programCounter[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END probe_programCounter[10]
  PIN probe_programCounter[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END probe_programCounter[11]
  PIN probe_programCounter[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END probe_programCounter[12]
  PIN probe_programCounter[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END probe_programCounter[13]
  PIN probe_programCounter[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END probe_programCounter[14]
  PIN probe_programCounter[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END probe_programCounter[15]
  PIN probe_programCounter[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END probe_programCounter[16]
  PIN probe_programCounter[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END probe_programCounter[17]
  PIN probe_programCounter[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END probe_programCounter[18]
  PIN probe_programCounter[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END probe_programCounter[19]
  PIN probe_programCounter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END probe_programCounter[1]
  PIN probe_programCounter[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END probe_programCounter[20]
  PIN probe_programCounter[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END probe_programCounter[21]
  PIN probe_programCounter[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END probe_programCounter[22]
  PIN probe_programCounter[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 0.000 348.590 4.000 ;
    END
  END probe_programCounter[23]
  PIN probe_programCounter[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END probe_programCounter[24]
  PIN probe_programCounter[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END probe_programCounter[25]
  PIN probe_programCounter[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END probe_programCounter[26]
  PIN probe_programCounter[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END probe_programCounter[27]
  PIN probe_programCounter[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END probe_programCounter[28]
  PIN probe_programCounter[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END probe_programCounter[29]
  PIN probe_programCounter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END probe_programCounter[2]
  PIN probe_programCounter[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END probe_programCounter[30]
  PIN probe_programCounter[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END probe_programCounter[31]
  PIN probe_programCounter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END probe_programCounter[3]
  PIN probe_programCounter[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END probe_programCounter[4]
  PIN probe_programCounter[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END probe_programCounter[5]
  PIN probe_programCounter[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END probe_programCounter[6]
  PIN probe_programCounter[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END probe_programCounter[7]
  PIN probe_programCounter[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END probe_programCounter[8]
  PIN probe_programCounter[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END probe_programCounter[9]
  PIN probe_state[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END probe_state[0]
  PIN probe_state[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END probe_state[1]
  PIN probe_takeBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END probe_takeBranch
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 886.960 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 896.000 380.330 900.000 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 896.000 390.910 900.000 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 896.000 401.490 900.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 896.000 412.070 900.000 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 886.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 886.960 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 2.080 450.000 2.680 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 6.160 450.000 6.760 ;
    END
  END wb_rst_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 444.360 886.805 ;
      LAYER met1 ;
        RECT 0.070 3.440 449.810 889.400 ;
      LAYER met2 ;
        RECT 0.090 895.720 4.870 898.125 ;
        RECT 5.710 895.720 15.450 898.125 ;
        RECT 16.290 895.720 26.030 898.125 ;
        RECT 26.870 895.720 36.610 898.125 ;
        RECT 37.450 895.720 47.650 898.125 ;
        RECT 48.490 895.720 58.230 898.125 ;
        RECT 59.070 895.720 68.810 898.125 ;
        RECT 69.650 895.720 79.850 898.125 ;
        RECT 80.690 895.720 90.430 898.125 ;
        RECT 91.270 895.720 101.010 898.125 ;
        RECT 101.850 895.720 111.590 898.125 ;
        RECT 112.430 895.720 122.630 898.125 ;
        RECT 123.470 895.720 133.210 898.125 ;
        RECT 134.050 895.720 143.790 898.125 ;
        RECT 144.630 895.720 154.830 898.125 ;
        RECT 155.670 895.720 165.410 898.125 ;
        RECT 166.250 895.720 175.990 898.125 ;
        RECT 176.830 895.720 186.570 898.125 ;
        RECT 187.410 895.720 197.610 898.125 ;
        RECT 198.450 895.720 208.190 898.125 ;
        RECT 209.030 895.720 218.770 898.125 ;
        RECT 219.610 895.720 229.810 898.125 ;
        RECT 230.650 895.720 240.390 898.125 ;
        RECT 241.230 895.720 250.970 898.125 ;
        RECT 251.810 895.720 261.550 898.125 ;
        RECT 262.390 895.720 272.590 898.125 ;
        RECT 273.430 895.720 283.170 898.125 ;
        RECT 284.010 895.720 293.750 898.125 ;
        RECT 294.590 895.720 304.790 898.125 ;
        RECT 305.630 895.720 315.370 898.125 ;
        RECT 316.210 895.720 325.950 898.125 ;
        RECT 326.790 895.720 336.530 898.125 ;
        RECT 337.370 895.720 347.570 898.125 ;
        RECT 348.410 895.720 358.150 898.125 ;
        RECT 358.990 895.720 368.730 898.125 ;
        RECT 369.570 895.720 379.770 898.125 ;
        RECT 380.610 895.720 390.350 898.125 ;
        RECT 391.190 895.720 400.930 898.125 ;
        RECT 401.770 895.720 411.510 898.125 ;
        RECT 412.350 895.720 422.550 898.125 ;
        RECT 423.390 895.720 433.130 898.125 ;
        RECT 433.970 895.720 443.710 898.125 ;
        RECT 444.550 895.720 449.790 898.125 ;
        RECT 0.090 4.280 449.790 895.720 ;
        RECT 0.090 2.195 3.490 4.280 ;
        RECT 4.330 2.195 10.850 4.280 ;
        RECT 11.690 2.195 18.210 4.280 ;
        RECT 19.050 2.195 25.570 4.280 ;
        RECT 26.410 2.195 33.390 4.280 ;
        RECT 34.230 2.195 40.750 4.280 ;
        RECT 41.590 2.195 48.110 4.280 ;
        RECT 48.950 2.195 55.930 4.280 ;
        RECT 56.770 2.195 63.290 4.280 ;
        RECT 64.130 2.195 70.650 4.280 ;
        RECT 71.490 2.195 78.470 4.280 ;
        RECT 79.310 2.195 85.830 4.280 ;
        RECT 86.670 2.195 93.190 4.280 ;
        RECT 94.030 2.195 100.550 4.280 ;
        RECT 101.390 2.195 108.370 4.280 ;
        RECT 109.210 2.195 115.730 4.280 ;
        RECT 116.570 2.195 123.090 4.280 ;
        RECT 123.930 2.195 130.910 4.280 ;
        RECT 131.750 2.195 138.270 4.280 ;
        RECT 139.110 2.195 145.630 4.280 ;
        RECT 146.470 2.195 153.450 4.280 ;
        RECT 154.290 2.195 160.810 4.280 ;
        RECT 161.650 2.195 168.170 4.280 ;
        RECT 169.010 2.195 175.530 4.280 ;
        RECT 176.370 2.195 183.350 4.280 ;
        RECT 184.190 2.195 190.710 4.280 ;
        RECT 191.550 2.195 198.070 4.280 ;
        RECT 198.910 2.195 205.890 4.280 ;
        RECT 206.730 2.195 213.250 4.280 ;
        RECT 214.090 2.195 220.610 4.280 ;
        RECT 221.450 2.195 228.430 4.280 ;
        RECT 229.270 2.195 235.790 4.280 ;
        RECT 236.630 2.195 243.150 4.280 ;
        RECT 243.990 2.195 250.510 4.280 ;
        RECT 251.350 2.195 258.330 4.280 ;
        RECT 259.170 2.195 265.690 4.280 ;
        RECT 266.530 2.195 273.050 4.280 ;
        RECT 273.890 2.195 280.870 4.280 ;
        RECT 281.710 2.195 288.230 4.280 ;
        RECT 289.070 2.195 295.590 4.280 ;
        RECT 296.430 2.195 303.410 4.280 ;
        RECT 304.250 2.195 310.770 4.280 ;
        RECT 311.610 2.195 318.130 4.280 ;
        RECT 318.970 2.195 325.490 4.280 ;
        RECT 326.330 2.195 333.310 4.280 ;
        RECT 334.150 2.195 340.670 4.280 ;
        RECT 341.510 2.195 348.030 4.280 ;
        RECT 348.870 2.195 355.850 4.280 ;
        RECT 356.690 2.195 363.210 4.280 ;
        RECT 364.050 2.195 370.570 4.280 ;
        RECT 371.410 2.195 378.390 4.280 ;
        RECT 379.230 2.195 385.750 4.280 ;
        RECT 386.590 2.195 393.110 4.280 ;
        RECT 393.950 2.195 400.470 4.280 ;
        RECT 401.310 2.195 408.290 4.280 ;
        RECT 409.130 2.195 415.650 4.280 ;
        RECT 416.490 2.195 423.010 4.280 ;
        RECT 423.850 2.195 430.830 4.280 ;
        RECT 431.670 2.195 438.190 4.280 ;
        RECT 439.030 2.195 445.550 4.280 ;
        RECT 446.390 2.195 449.790 4.280 ;
      LAYER met3 ;
        RECT 4.400 897.240 445.600 898.105 ;
        RECT 0.065 894.560 449.815 897.240 ;
        RECT 0.065 893.880 445.600 894.560 ;
        RECT 4.400 893.160 445.600 893.880 ;
        RECT 4.400 892.480 449.815 893.160 ;
        RECT 0.065 889.800 449.815 892.480 ;
        RECT 0.065 889.120 445.600 889.800 ;
        RECT 4.400 888.400 445.600 889.120 ;
        RECT 4.400 887.720 449.815 888.400 ;
        RECT 0.065 885.720 449.815 887.720 ;
        RECT 0.065 885.040 445.600 885.720 ;
        RECT 4.400 884.320 445.600 885.040 ;
        RECT 4.400 883.640 449.815 884.320 ;
        RECT 0.065 880.960 449.815 883.640 ;
        RECT 0.065 880.280 445.600 880.960 ;
        RECT 4.400 879.560 445.600 880.280 ;
        RECT 4.400 878.880 449.815 879.560 ;
        RECT 0.065 876.880 449.815 878.880 ;
        RECT 0.065 875.520 445.600 876.880 ;
        RECT 4.400 875.480 445.600 875.520 ;
        RECT 4.400 874.120 449.815 875.480 ;
        RECT 0.065 872.800 449.815 874.120 ;
        RECT 0.065 871.400 445.600 872.800 ;
        RECT 0.065 870.760 449.815 871.400 ;
        RECT 4.400 869.360 449.815 870.760 ;
        RECT 0.065 868.040 449.815 869.360 ;
        RECT 0.065 866.680 445.600 868.040 ;
        RECT 4.400 866.640 445.600 866.680 ;
        RECT 4.400 865.280 449.815 866.640 ;
        RECT 0.065 863.960 449.815 865.280 ;
        RECT 0.065 862.560 445.600 863.960 ;
        RECT 0.065 861.920 449.815 862.560 ;
        RECT 4.400 860.520 449.815 861.920 ;
        RECT 0.065 859.200 449.815 860.520 ;
        RECT 0.065 857.800 445.600 859.200 ;
        RECT 0.065 857.160 449.815 857.800 ;
        RECT 4.400 855.760 449.815 857.160 ;
        RECT 0.065 855.120 449.815 855.760 ;
        RECT 0.065 853.720 445.600 855.120 ;
        RECT 0.065 853.080 449.815 853.720 ;
        RECT 4.400 851.680 449.815 853.080 ;
        RECT 0.065 850.360 449.815 851.680 ;
        RECT 0.065 848.960 445.600 850.360 ;
        RECT 0.065 848.320 449.815 848.960 ;
        RECT 4.400 846.920 449.815 848.320 ;
        RECT 0.065 846.280 449.815 846.920 ;
        RECT 0.065 844.880 445.600 846.280 ;
        RECT 0.065 843.560 449.815 844.880 ;
        RECT 4.400 842.200 449.815 843.560 ;
        RECT 4.400 842.160 445.600 842.200 ;
        RECT 0.065 840.800 445.600 842.160 ;
        RECT 0.065 838.800 449.815 840.800 ;
        RECT 4.400 837.440 449.815 838.800 ;
        RECT 4.400 837.400 445.600 837.440 ;
        RECT 0.065 836.040 445.600 837.400 ;
        RECT 0.065 834.720 449.815 836.040 ;
        RECT 4.400 833.360 449.815 834.720 ;
        RECT 4.400 833.320 445.600 833.360 ;
        RECT 0.065 831.960 445.600 833.320 ;
        RECT 0.065 829.960 449.815 831.960 ;
        RECT 4.400 828.600 449.815 829.960 ;
        RECT 4.400 828.560 445.600 828.600 ;
        RECT 0.065 827.200 445.600 828.560 ;
        RECT 0.065 825.200 449.815 827.200 ;
        RECT 4.400 824.520 449.815 825.200 ;
        RECT 4.400 823.800 445.600 824.520 ;
        RECT 0.065 823.120 445.600 823.800 ;
        RECT 0.065 821.120 449.815 823.120 ;
        RECT 4.400 819.760 449.815 821.120 ;
        RECT 4.400 819.720 445.600 819.760 ;
        RECT 0.065 818.360 445.600 819.720 ;
        RECT 0.065 816.360 449.815 818.360 ;
        RECT 4.400 815.680 449.815 816.360 ;
        RECT 4.400 814.960 445.600 815.680 ;
        RECT 0.065 814.280 445.600 814.960 ;
        RECT 0.065 811.600 449.815 814.280 ;
        RECT 4.400 810.200 445.600 811.600 ;
        RECT 0.065 806.840 449.815 810.200 ;
        RECT 4.400 805.440 445.600 806.840 ;
        RECT 0.065 802.760 449.815 805.440 ;
        RECT 4.400 801.360 445.600 802.760 ;
        RECT 0.065 798.000 449.815 801.360 ;
        RECT 4.400 796.600 445.600 798.000 ;
        RECT 0.065 793.920 449.815 796.600 ;
        RECT 0.065 793.240 445.600 793.920 ;
        RECT 4.400 792.520 445.600 793.240 ;
        RECT 4.400 791.840 449.815 792.520 ;
        RECT 0.065 789.160 449.815 791.840 ;
        RECT 0.065 788.480 445.600 789.160 ;
        RECT 4.400 787.760 445.600 788.480 ;
        RECT 4.400 787.080 449.815 787.760 ;
        RECT 0.065 785.080 449.815 787.080 ;
        RECT 0.065 784.400 445.600 785.080 ;
        RECT 4.400 783.680 445.600 784.400 ;
        RECT 4.400 783.000 449.815 783.680 ;
        RECT 0.065 781.000 449.815 783.000 ;
        RECT 0.065 779.640 445.600 781.000 ;
        RECT 4.400 779.600 445.600 779.640 ;
        RECT 4.400 778.240 449.815 779.600 ;
        RECT 0.065 776.240 449.815 778.240 ;
        RECT 0.065 774.880 445.600 776.240 ;
        RECT 4.400 774.840 445.600 774.880 ;
        RECT 4.400 773.480 449.815 774.840 ;
        RECT 0.065 772.160 449.815 773.480 ;
        RECT 0.065 770.800 445.600 772.160 ;
        RECT 4.400 770.760 445.600 770.800 ;
        RECT 4.400 769.400 449.815 770.760 ;
        RECT 0.065 767.400 449.815 769.400 ;
        RECT 0.065 766.040 445.600 767.400 ;
        RECT 4.400 766.000 445.600 766.040 ;
        RECT 4.400 764.640 449.815 766.000 ;
        RECT 0.065 763.320 449.815 764.640 ;
        RECT 0.065 761.920 445.600 763.320 ;
        RECT 0.065 761.280 449.815 761.920 ;
        RECT 4.400 759.880 449.815 761.280 ;
        RECT 0.065 758.560 449.815 759.880 ;
        RECT 0.065 757.160 445.600 758.560 ;
        RECT 0.065 756.520 449.815 757.160 ;
        RECT 4.400 755.120 449.815 756.520 ;
        RECT 0.065 754.480 449.815 755.120 ;
        RECT 0.065 753.080 445.600 754.480 ;
        RECT 0.065 752.440 449.815 753.080 ;
        RECT 4.400 751.040 449.815 752.440 ;
        RECT 0.065 750.400 449.815 751.040 ;
        RECT 0.065 749.000 445.600 750.400 ;
        RECT 0.065 747.680 449.815 749.000 ;
        RECT 4.400 746.280 449.815 747.680 ;
        RECT 0.065 745.640 449.815 746.280 ;
        RECT 0.065 744.240 445.600 745.640 ;
        RECT 0.065 742.920 449.815 744.240 ;
        RECT 4.400 741.560 449.815 742.920 ;
        RECT 4.400 741.520 445.600 741.560 ;
        RECT 0.065 740.160 445.600 741.520 ;
        RECT 0.065 738.840 449.815 740.160 ;
        RECT 4.400 737.440 449.815 738.840 ;
        RECT 0.065 736.800 449.815 737.440 ;
        RECT 0.065 735.400 445.600 736.800 ;
        RECT 0.065 734.080 449.815 735.400 ;
        RECT 4.400 732.720 449.815 734.080 ;
        RECT 4.400 732.680 445.600 732.720 ;
        RECT 0.065 731.320 445.600 732.680 ;
        RECT 0.065 729.320 449.815 731.320 ;
        RECT 4.400 727.960 449.815 729.320 ;
        RECT 4.400 727.920 445.600 727.960 ;
        RECT 0.065 726.560 445.600 727.920 ;
        RECT 0.065 724.560 449.815 726.560 ;
        RECT 4.400 723.880 449.815 724.560 ;
        RECT 4.400 723.160 445.600 723.880 ;
        RECT 0.065 722.480 445.600 723.160 ;
        RECT 0.065 720.480 449.815 722.480 ;
        RECT 4.400 719.800 449.815 720.480 ;
        RECT 4.400 719.080 445.600 719.800 ;
        RECT 0.065 718.400 445.600 719.080 ;
        RECT 0.065 715.720 449.815 718.400 ;
        RECT 4.400 715.040 449.815 715.720 ;
        RECT 4.400 714.320 445.600 715.040 ;
        RECT 0.065 713.640 445.600 714.320 ;
        RECT 0.065 710.960 449.815 713.640 ;
        RECT 4.400 709.560 445.600 710.960 ;
        RECT 0.065 706.880 449.815 709.560 ;
        RECT 4.400 706.200 449.815 706.880 ;
        RECT 4.400 705.480 445.600 706.200 ;
        RECT 0.065 704.800 445.600 705.480 ;
        RECT 0.065 702.120 449.815 704.800 ;
        RECT 4.400 700.720 445.600 702.120 ;
        RECT 0.065 697.360 449.815 700.720 ;
        RECT 4.400 695.960 445.600 697.360 ;
        RECT 0.065 693.280 449.815 695.960 ;
        RECT 0.065 692.600 445.600 693.280 ;
        RECT 4.400 691.880 445.600 692.600 ;
        RECT 4.400 691.200 449.815 691.880 ;
        RECT 0.065 689.200 449.815 691.200 ;
        RECT 0.065 688.520 445.600 689.200 ;
        RECT 4.400 687.800 445.600 688.520 ;
        RECT 4.400 687.120 449.815 687.800 ;
        RECT 0.065 684.440 449.815 687.120 ;
        RECT 0.065 683.760 445.600 684.440 ;
        RECT 4.400 683.040 445.600 683.760 ;
        RECT 4.400 682.360 449.815 683.040 ;
        RECT 0.065 680.360 449.815 682.360 ;
        RECT 0.065 679.000 445.600 680.360 ;
        RECT 4.400 678.960 445.600 679.000 ;
        RECT 4.400 677.600 449.815 678.960 ;
        RECT 0.065 675.600 449.815 677.600 ;
        RECT 0.065 674.240 445.600 675.600 ;
        RECT 4.400 674.200 445.600 674.240 ;
        RECT 4.400 672.840 449.815 674.200 ;
        RECT 0.065 671.520 449.815 672.840 ;
        RECT 0.065 670.160 445.600 671.520 ;
        RECT 4.400 670.120 445.600 670.160 ;
        RECT 4.400 668.760 449.815 670.120 ;
        RECT 0.065 666.760 449.815 668.760 ;
        RECT 0.065 665.400 445.600 666.760 ;
        RECT 4.400 665.360 445.600 665.400 ;
        RECT 4.400 664.000 449.815 665.360 ;
        RECT 0.065 662.680 449.815 664.000 ;
        RECT 0.065 661.280 445.600 662.680 ;
        RECT 0.065 660.640 449.815 661.280 ;
        RECT 4.400 659.240 449.815 660.640 ;
        RECT 0.065 658.600 449.815 659.240 ;
        RECT 0.065 657.200 445.600 658.600 ;
        RECT 0.065 656.560 449.815 657.200 ;
        RECT 4.400 655.160 449.815 656.560 ;
        RECT 0.065 653.840 449.815 655.160 ;
        RECT 0.065 652.440 445.600 653.840 ;
        RECT 0.065 651.800 449.815 652.440 ;
        RECT 4.400 650.400 449.815 651.800 ;
        RECT 0.065 649.760 449.815 650.400 ;
        RECT 0.065 648.360 445.600 649.760 ;
        RECT 0.065 647.040 449.815 648.360 ;
        RECT 4.400 645.640 449.815 647.040 ;
        RECT 0.065 645.000 449.815 645.640 ;
        RECT 0.065 643.600 445.600 645.000 ;
        RECT 0.065 642.280 449.815 643.600 ;
        RECT 4.400 640.920 449.815 642.280 ;
        RECT 4.400 640.880 445.600 640.920 ;
        RECT 0.065 639.520 445.600 640.880 ;
        RECT 0.065 638.200 449.815 639.520 ;
        RECT 4.400 636.800 449.815 638.200 ;
        RECT 0.065 636.160 449.815 636.800 ;
        RECT 0.065 634.760 445.600 636.160 ;
        RECT 0.065 633.440 449.815 634.760 ;
        RECT 4.400 632.080 449.815 633.440 ;
        RECT 4.400 632.040 445.600 632.080 ;
        RECT 0.065 630.680 445.600 632.040 ;
        RECT 0.065 628.680 449.815 630.680 ;
        RECT 4.400 628.000 449.815 628.680 ;
        RECT 4.400 627.280 445.600 628.000 ;
        RECT 0.065 626.600 445.600 627.280 ;
        RECT 0.065 624.600 449.815 626.600 ;
        RECT 4.400 623.240 449.815 624.600 ;
        RECT 4.400 623.200 445.600 623.240 ;
        RECT 0.065 621.840 445.600 623.200 ;
        RECT 0.065 619.840 449.815 621.840 ;
        RECT 4.400 619.160 449.815 619.840 ;
        RECT 4.400 618.440 445.600 619.160 ;
        RECT 0.065 617.760 445.600 618.440 ;
        RECT 0.065 615.080 449.815 617.760 ;
        RECT 4.400 614.400 449.815 615.080 ;
        RECT 4.400 613.680 445.600 614.400 ;
        RECT 0.065 613.000 445.600 613.680 ;
        RECT 0.065 610.320 449.815 613.000 ;
        RECT 4.400 608.920 445.600 610.320 ;
        RECT 0.065 606.240 449.815 608.920 ;
        RECT 4.400 605.560 449.815 606.240 ;
        RECT 4.400 604.840 445.600 605.560 ;
        RECT 0.065 604.160 445.600 604.840 ;
        RECT 0.065 601.480 449.815 604.160 ;
        RECT 4.400 600.080 445.600 601.480 ;
        RECT 0.065 597.400 449.815 600.080 ;
        RECT 0.065 596.720 445.600 597.400 ;
        RECT 4.400 596.000 445.600 596.720 ;
        RECT 4.400 595.320 449.815 596.000 ;
        RECT 0.065 592.640 449.815 595.320 ;
        RECT 0.065 591.960 445.600 592.640 ;
        RECT 4.400 591.240 445.600 591.960 ;
        RECT 4.400 590.560 449.815 591.240 ;
        RECT 0.065 588.560 449.815 590.560 ;
        RECT 0.065 587.880 445.600 588.560 ;
        RECT 4.400 587.160 445.600 587.880 ;
        RECT 4.400 586.480 449.815 587.160 ;
        RECT 0.065 583.800 449.815 586.480 ;
        RECT 0.065 583.120 445.600 583.800 ;
        RECT 4.400 582.400 445.600 583.120 ;
        RECT 4.400 581.720 449.815 582.400 ;
        RECT 0.065 579.720 449.815 581.720 ;
        RECT 0.065 578.360 445.600 579.720 ;
        RECT 4.400 578.320 445.600 578.360 ;
        RECT 4.400 576.960 449.815 578.320 ;
        RECT 0.065 574.960 449.815 576.960 ;
        RECT 0.065 574.280 445.600 574.960 ;
        RECT 4.400 573.560 445.600 574.280 ;
        RECT 4.400 572.880 449.815 573.560 ;
        RECT 0.065 570.880 449.815 572.880 ;
        RECT 0.065 569.520 445.600 570.880 ;
        RECT 4.400 569.480 445.600 569.520 ;
        RECT 4.400 568.120 449.815 569.480 ;
        RECT 0.065 566.800 449.815 568.120 ;
        RECT 0.065 565.400 445.600 566.800 ;
        RECT 0.065 564.760 449.815 565.400 ;
        RECT 4.400 563.360 449.815 564.760 ;
        RECT 0.065 562.040 449.815 563.360 ;
        RECT 0.065 560.640 445.600 562.040 ;
        RECT 0.065 560.000 449.815 560.640 ;
        RECT 4.400 558.600 449.815 560.000 ;
        RECT 0.065 557.960 449.815 558.600 ;
        RECT 0.065 556.560 445.600 557.960 ;
        RECT 0.065 555.920 449.815 556.560 ;
        RECT 4.400 554.520 449.815 555.920 ;
        RECT 0.065 553.200 449.815 554.520 ;
        RECT 0.065 551.800 445.600 553.200 ;
        RECT 0.065 551.160 449.815 551.800 ;
        RECT 4.400 549.760 449.815 551.160 ;
        RECT 0.065 549.120 449.815 549.760 ;
        RECT 0.065 547.720 445.600 549.120 ;
        RECT 0.065 546.400 449.815 547.720 ;
        RECT 4.400 545.000 449.815 546.400 ;
        RECT 0.065 544.360 449.815 545.000 ;
        RECT 0.065 542.960 445.600 544.360 ;
        RECT 0.065 542.320 449.815 542.960 ;
        RECT 4.400 540.920 449.815 542.320 ;
        RECT 0.065 540.280 449.815 540.920 ;
        RECT 0.065 538.880 445.600 540.280 ;
        RECT 0.065 537.560 449.815 538.880 ;
        RECT 4.400 536.200 449.815 537.560 ;
        RECT 4.400 536.160 445.600 536.200 ;
        RECT 0.065 534.800 445.600 536.160 ;
        RECT 0.065 532.800 449.815 534.800 ;
        RECT 4.400 531.440 449.815 532.800 ;
        RECT 4.400 531.400 445.600 531.440 ;
        RECT 0.065 530.040 445.600 531.400 ;
        RECT 0.065 528.040 449.815 530.040 ;
        RECT 4.400 527.360 449.815 528.040 ;
        RECT 4.400 526.640 445.600 527.360 ;
        RECT 0.065 525.960 445.600 526.640 ;
        RECT 0.065 523.960 449.815 525.960 ;
        RECT 4.400 522.600 449.815 523.960 ;
        RECT 4.400 522.560 445.600 522.600 ;
        RECT 0.065 521.200 445.600 522.560 ;
        RECT 0.065 519.200 449.815 521.200 ;
        RECT 4.400 518.520 449.815 519.200 ;
        RECT 4.400 517.800 445.600 518.520 ;
        RECT 0.065 517.120 445.600 517.800 ;
        RECT 0.065 514.440 449.815 517.120 ;
        RECT 4.400 513.760 449.815 514.440 ;
        RECT 4.400 513.040 445.600 513.760 ;
        RECT 0.065 512.360 445.600 513.040 ;
        RECT 0.065 510.360 449.815 512.360 ;
        RECT 4.400 509.680 449.815 510.360 ;
        RECT 4.400 508.960 445.600 509.680 ;
        RECT 0.065 508.280 445.600 508.960 ;
        RECT 0.065 505.600 449.815 508.280 ;
        RECT 4.400 504.200 445.600 505.600 ;
        RECT 0.065 500.840 449.815 504.200 ;
        RECT 4.400 499.440 445.600 500.840 ;
        RECT 0.065 496.760 449.815 499.440 ;
        RECT 0.065 496.080 445.600 496.760 ;
        RECT 4.400 495.360 445.600 496.080 ;
        RECT 4.400 494.680 449.815 495.360 ;
        RECT 0.065 492.000 449.815 494.680 ;
        RECT 4.400 490.600 445.600 492.000 ;
        RECT 0.065 487.920 449.815 490.600 ;
        RECT 0.065 487.240 445.600 487.920 ;
        RECT 4.400 486.520 445.600 487.240 ;
        RECT 4.400 485.840 449.815 486.520 ;
        RECT 0.065 483.160 449.815 485.840 ;
        RECT 0.065 482.480 445.600 483.160 ;
        RECT 4.400 481.760 445.600 482.480 ;
        RECT 4.400 481.080 449.815 481.760 ;
        RECT 0.065 479.080 449.815 481.080 ;
        RECT 0.065 477.720 445.600 479.080 ;
        RECT 4.400 477.680 445.600 477.720 ;
        RECT 4.400 476.320 449.815 477.680 ;
        RECT 0.065 475.000 449.815 476.320 ;
        RECT 0.065 473.640 445.600 475.000 ;
        RECT 4.400 473.600 445.600 473.640 ;
        RECT 4.400 472.240 449.815 473.600 ;
        RECT 0.065 470.240 449.815 472.240 ;
        RECT 0.065 468.880 445.600 470.240 ;
        RECT 4.400 468.840 445.600 468.880 ;
        RECT 4.400 467.480 449.815 468.840 ;
        RECT 0.065 466.160 449.815 467.480 ;
        RECT 0.065 464.760 445.600 466.160 ;
        RECT 0.065 464.120 449.815 464.760 ;
        RECT 4.400 462.720 449.815 464.120 ;
        RECT 0.065 461.400 449.815 462.720 ;
        RECT 0.065 460.040 445.600 461.400 ;
        RECT 4.400 460.000 445.600 460.040 ;
        RECT 4.400 458.640 449.815 460.000 ;
        RECT 0.065 457.320 449.815 458.640 ;
        RECT 0.065 455.920 445.600 457.320 ;
        RECT 0.065 455.280 449.815 455.920 ;
        RECT 4.400 453.880 449.815 455.280 ;
        RECT 0.065 453.240 449.815 453.880 ;
        RECT 0.065 451.840 445.600 453.240 ;
        RECT 0.065 450.520 449.815 451.840 ;
        RECT 4.400 449.120 449.815 450.520 ;
        RECT 0.065 448.480 449.815 449.120 ;
        RECT 0.065 447.080 445.600 448.480 ;
        RECT 0.065 445.760 449.815 447.080 ;
        RECT 4.400 444.400 449.815 445.760 ;
        RECT 4.400 444.360 445.600 444.400 ;
        RECT 0.065 443.000 445.600 444.360 ;
        RECT 0.065 441.680 449.815 443.000 ;
        RECT 4.400 440.280 449.815 441.680 ;
        RECT 0.065 439.640 449.815 440.280 ;
        RECT 0.065 438.240 445.600 439.640 ;
        RECT 0.065 436.920 449.815 438.240 ;
        RECT 4.400 435.560 449.815 436.920 ;
        RECT 4.400 435.520 445.600 435.560 ;
        RECT 0.065 434.160 445.600 435.520 ;
        RECT 0.065 432.160 449.815 434.160 ;
        RECT 4.400 430.800 449.815 432.160 ;
        RECT 4.400 430.760 445.600 430.800 ;
        RECT 0.065 429.400 445.600 430.760 ;
        RECT 0.065 428.080 449.815 429.400 ;
        RECT 4.400 426.720 449.815 428.080 ;
        RECT 4.400 426.680 445.600 426.720 ;
        RECT 0.065 425.320 445.600 426.680 ;
        RECT 0.065 423.320 449.815 425.320 ;
        RECT 4.400 422.640 449.815 423.320 ;
        RECT 4.400 421.920 445.600 422.640 ;
        RECT 0.065 421.240 445.600 421.920 ;
        RECT 0.065 418.560 449.815 421.240 ;
        RECT 4.400 417.880 449.815 418.560 ;
        RECT 4.400 417.160 445.600 417.880 ;
        RECT 0.065 416.480 445.600 417.160 ;
        RECT 0.065 413.800 449.815 416.480 ;
        RECT 4.400 412.400 445.600 413.800 ;
        RECT 0.065 409.720 449.815 412.400 ;
        RECT 4.400 409.040 449.815 409.720 ;
        RECT 4.400 408.320 445.600 409.040 ;
        RECT 0.065 407.640 445.600 408.320 ;
        RECT 0.065 404.960 449.815 407.640 ;
        RECT 4.400 403.560 445.600 404.960 ;
        RECT 0.065 400.200 449.815 403.560 ;
        RECT 4.400 398.800 445.600 400.200 ;
        RECT 0.065 396.120 449.815 398.800 ;
        RECT 0.065 395.440 445.600 396.120 ;
        RECT 4.400 394.720 445.600 395.440 ;
        RECT 4.400 394.040 449.815 394.720 ;
        RECT 0.065 392.040 449.815 394.040 ;
        RECT 0.065 391.360 445.600 392.040 ;
        RECT 4.400 390.640 445.600 391.360 ;
        RECT 4.400 389.960 449.815 390.640 ;
        RECT 0.065 387.280 449.815 389.960 ;
        RECT 0.065 386.600 445.600 387.280 ;
        RECT 4.400 385.880 445.600 386.600 ;
        RECT 4.400 385.200 449.815 385.880 ;
        RECT 0.065 383.200 449.815 385.200 ;
        RECT 0.065 381.840 445.600 383.200 ;
        RECT 4.400 381.800 445.600 381.840 ;
        RECT 4.400 380.440 449.815 381.800 ;
        RECT 0.065 378.440 449.815 380.440 ;
        RECT 0.065 377.760 445.600 378.440 ;
        RECT 4.400 377.040 445.600 377.760 ;
        RECT 4.400 376.360 449.815 377.040 ;
        RECT 0.065 374.360 449.815 376.360 ;
        RECT 0.065 373.000 445.600 374.360 ;
        RECT 4.400 372.960 445.600 373.000 ;
        RECT 4.400 371.600 449.815 372.960 ;
        RECT 0.065 369.600 449.815 371.600 ;
        RECT 0.065 368.240 445.600 369.600 ;
        RECT 4.400 368.200 445.600 368.240 ;
        RECT 4.400 366.840 449.815 368.200 ;
        RECT 0.065 365.520 449.815 366.840 ;
        RECT 0.065 364.120 445.600 365.520 ;
        RECT 0.065 363.480 449.815 364.120 ;
        RECT 4.400 362.080 449.815 363.480 ;
        RECT 0.065 361.440 449.815 362.080 ;
        RECT 0.065 360.040 445.600 361.440 ;
        RECT 0.065 359.400 449.815 360.040 ;
        RECT 4.400 358.000 449.815 359.400 ;
        RECT 0.065 356.680 449.815 358.000 ;
        RECT 0.065 355.280 445.600 356.680 ;
        RECT 0.065 354.640 449.815 355.280 ;
        RECT 4.400 353.240 449.815 354.640 ;
        RECT 0.065 352.600 449.815 353.240 ;
        RECT 0.065 351.200 445.600 352.600 ;
        RECT 0.065 349.880 449.815 351.200 ;
        RECT 4.400 348.480 449.815 349.880 ;
        RECT 0.065 347.840 449.815 348.480 ;
        RECT 0.065 346.440 445.600 347.840 ;
        RECT 0.065 345.800 449.815 346.440 ;
        RECT 4.400 344.400 449.815 345.800 ;
        RECT 0.065 343.760 449.815 344.400 ;
        RECT 0.065 342.360 445.600 343.760 ;
        RECT 0.065 341.040 449.815 342.360 ;
        RECT 4.400 339.640 449.815 341.040 ;
        RECT 0.065 339.000 449.815 339.640 ;
        RECT 0.065 337.600 445.600 339.000 ;
        RECT 0.065 336.280 449.815 337.600 ;
        RECT 4.400 334.920 449.815 336.280 ;
        RECT 4.400 334.880 445.600 334.920 ;
        RECT 0.065 333.520 445.600 334.880 ;
        RECT 0.065 331.520 449.815 333.520 ;
        RECT 4.400 330.840 449.815 331.520 ;
        RECT 4.400 330.120 445.600 330.840 ;
        RECT 0.065 329.440 445.600 330.120 ;
        RECT 0.065 327.440 449.815 329.440 ;
        RECT 4.400 326.080 449.815 327.440 ;
        RECT 4.400 326.040 445.600 326.080 ;
        RECT 0.065 324.680 445.600 326.040 ;
        RECT 0.065 322.680 449.815 324.680 ;
        RECT 4.400 322.000 449.815 322.680 ;
        RECT 4.400 321.280 445.600 322.000 ;
        RECT 0.065 320.600 445.600 321.280 ;
        RECT 0.065 317.920 449.815 320.600 ;
        RECT 4.400 317.240 449.815 317.920 ;
        RECT 4.400 316.520 445.600 317.240 ;
        RECT 0.065 315.840 445.600 316.520 ;
        RECT 0.065 313.840 449.815 315.840 ;
        RECT 4.400 313.160 449.815 313.840 ;
        RECT 4.400 312.440 445.600 313.160 ;
        RECT 0.065 311.760 445.600 312.440 ;
        RECT 0.065 309.080 449.815 311.760 ;
        RECT 4.400 308.400 449.815 309.080 ;
        RECT 4.400 307.680 445.600 308.400 ;
        RECT 0.065 307.000 445.600 307.680 ;
        RECT 0.065 304.320 449.815 307.000 ;
        RECT 4.400 302.920 445.600 304.320 ;
        RECT 0.065 300.240 449.815 302.920 ;
        RECT 0.065 299.560 445.600 300.240 ;
        RECT 4.400 298.840 445.600 299.560 ;
        RECT 4.400 298.160 449.815 298.840 ;
        RECT 0.065 295.480 449.815 298.160 ;
        RECT 4.400 294.080 445.600 295.480 ;
        RECT 0.065 291.400 449.815 294.080 ;
        RECT 0.065 290.720 445.600 291.400 ;
        RECT 4.400 290.000 445.600 290.720 ;
        RECT 4.400 289.320 449.815 290.000 ;
        RECT 0.065 286.640 449.815 289.320 ;
        RECT 0.065 285.960 445.600 286.640 ;
        RECT 4.400 285.240 445.600 285.960 ;
        RECT 4.400 284.560 449.815 285.240 ;
        RECT 0.065 282.560 449.815 284.560 ;
        RECT 0.065 281.200 445.600 282.560 ;
        RECT 4.400 281.160 445.600 281.200 ;
        RECT 4.400 279.800 449.815 281.160 ;
        RECT 0.065 277.800 449.815 279.800 ;
        RECT 0.065 277.120 445.600 277.800 ;
        RECT 4.400 276.400 445.600 277.120 ;
        RECT 4.400 275.720 449.815 276.400 ;
        RECT 0.065 273.720 449.815 275.720 ;
        RECT 0.065 272.360 445.600 273.720 ;
        RECT 4.400 272.320 445.600 272.360 ;
        RECT 4.400 270.960 449.815 272.320 ;
        RECT 0.065 269.640 449.815 270.960 ;
        RECT 0.065 268.240 445.600 269.640 ;
        RECT 0.065 267.600 449.815 268.240 ;
        RECT 4.400 266.200 449.815 267.600 ;
        RECT 0.065 264.880 449.815 266.200 ;
        RECT 0.065 263.520 445.600 264.880 ;
        RECT 4.400 263.480 445.600 263.520 ;
        RECT 4.400 262.120 449.815 263.480 ;
        RECT 0.065 260.800 449.815 262.120 ;
        RECT 0.065 259.400 445.600 260.800 ;
        RECT 0.065 258.760 449.815 259.400 ;
        RECT 4.400 257.360 449.815 258.760 ;
        RECT 0.065 256.040 449.815 257.360 ;
        RECT 0.065 254.640 445.600 256.040 ;
        RECT 0.065 254.000 449.815 254.640 ;
        RECT 4.400 252.600 449.815 254.000 ;
        RECT 0.065 251.960 449.815 252.600 ;
        RECT 0.065 250.560 445.600 251.960 ;
        RECT 0.065 249.240 449.815 250.560 ;
        RECT 4.400 247.840 449.815 249.240 ;
        RECT 0.065 247.200 449.815 247.840 ;
        RECT 0.065 245.800 445.600 247.200 ;
        RECT 0.065 245.160 449.815 245.800 ;
        RECT 4.400 243.760 449.815 245.160 ;
        RECT 0.065 243.120 449.815 243.760 ;
        RECT 0.065 241.720 445.600 243.120 ;
        RECT 0.065 240.400 449.815 241.720 ;
        RECT 4.400 239.040 449.815 240.400 ;
        RECT 4.400 239.000 445.600 239.040 ;
        RECT 0.065 237.640 445.600 239.000 ;
        RECT 0.065 235.640 449.815 237.640 ;
        RECT 4.400 234.280 449.815 235.640 ;
        RECT 4.400 234.240 445.600 234.280 ;
        RECT 0.065 232.880 445.600 234.240 ;
        RECT 0.065 231.560 449.815 232.880 ;
        RECT 4.400 230.200 449.815 231.560 ;
        RECT 4.400 230.160 445.600 230.200 ;
        RECT 0.065 228.800 445.600 230.160 ;
        RECT 0.065 226.800 449.815 228.800 ;
        RECT 4.400 225.440 449.815 226.800 ;
        RECT 4.400 225.400 445.600 225.440 ;
        RECT 0.065 224.040 445.600 225.400 ;
        RECT 0.065 222.040 449.815 224.040 ;
        RECT 4.400 221.360 449.815 222.040 ;
        RECT 4.400 220.640 445.600 221.360 ;
        RECT 0.065 219.960 445.600 220.640 ;
        RECT 0.065 217.280 449.815 219.960 ;
        RECT 4.400 216.600 449.815 217.280 ;
        RECT 4.400 215.880 445.600 216.600 ;
        RECT 0.065 215.200 445.600 215.880 ;
        RECT 0.065 213.200 449.815 215.200 ;
        RECT 4.400 212.520 449.815 213.200 ;
        RECT 4.400 211.800 445.600 212.520 ;
        RECT 0.065 211.120 445.600 211.800 ;
        RECT 0.065 208.440 449.815 211.120 ;
        RECT 4.400 207.040 445.600 208.440 ;
        RECT 0.065 203.680 449.815 207.040 ;
        RECT 4.400 202.280 445.600 203.680 ;
        RECT 0.065 199.600 449.815 202.280 ;
        RECT 0.065 198.920 445.600 199.600 ;
        RECT 4.400 198.200 445.600 198.920 ;
        RECT 4.400 197.520 449.815 198.200 ;
        RECT 0.065 194.840 449.815 197.520 ;
        RECT 4.400 193.440 445.600 194.840 ;
        RECT 0.065 190.760 449.815 193.440 ;
        RECT 0.065 190.080 445.600 190.760 ;
        RECT 4.400 189.360 445.600 190.080 ;
        RECT 4.400 188.680 449.815 189.360 ;
        RECT 0.065 186.000 449.815 188.680 ;
        RECT 0.065 185.320 445.600 186.000 ;
        RECT 4.400 184.600 445.600 185.320 ;
        RECT 4.400 183.920 449.815 184.600 ;
        RECT 0.065 181.920 449.815 183.920 ;
        RECT 0.065 181.240 445.600 181.920 ;
        RECT 4.400 180.520 445.600 181.240 ;
        RECT 4.400 179.840 449.815 180.520 ;
        RECT 0.065 177.840 449.815 179.840 ;
        RECT 0.065 176.480 445.600 177.840 ;
        RECT 4.400 176.440 445.600 176.480 ;
        RECT 4.400 175.080 449.815 176.440 ;
        RECT 0.065 173.080 449.815 175.080 ;
        RECT 0.065 171.720 445.600 173.080 ;
        RECT 4.400 171.680 445.600 171.720 ;
        RECT 4.400 170.320 449.815 171.680 ;
        RECT 0.065 169.000 449.815 170.320 ;
        RECT 0.065 167.600 445.600 169.000 ;
        RECT 0.065 166.960 449.815 167.600 ;
        RECT 4.400 165.560 449.815 166.960 ;
        RECT 0.065 164.240 449.815 165.560 ;
        RECT 0.065 162.880 445.600 164.240 ;
        RECT 4.400 162.840 445.600 162.880 ;
        RECT 4.400 161.480 449.815 162.840 ;
        RECT 0.065 160.160 449.815 161.480 ;
        RECT 0.065 158.760 445.600 160.160 ;
        RECT 0.065 158.120 449.815 158.760 ;
        RECT 4.400 156.720 449.815 158.120 ;
        RECT 0.065 155.400 449.815 156.720 ;
        RECT 0.065 154.000 445.600 155.400 ;
        RECT 0.065 153.360 449.815 154.000 ;
        RECT 4.400 151.960 449.815 153.360 ;
        RECT 0.065 151.320 449.815 151.960 ;
        RECT 0.065 149.920 445.600 151.320 ;
        RECT 0.065 149.280 449.815 149.920 ;
        RECT 4.400 147.880 449.815 149.280 ;
        RECT 0.065 147.240 449.815 147.880 ;
        RECT 0.065 145.840 445.600 147.240 ;
        RECT 0.065 144.520 449.815 145.840 ;
        RECT 4.400 143.120 449.815 144.520 ;
        RECT 0.065 142.480 449.815 143.120 ;
        RECT 0.065 141.080 445.600 142.480 ;
        RECT 0.065 139.760 449.815 141.080 ;
        RECT 4.400 138.400 449.815 139.760 ;
        RECT 4.400 138.360 445.600 138.400 ;
        RECT 0.065 137.000 445.600 138.360 ;
        RECT 0.065 135.000 449.815 137.000 ;
        RECT 4.400 133.640 449.815 135.000 ;
        RECT 4.400 133.600 445.600 133.640 ;
        RECT 0.065 132.240 445.600 133.600 ;
        RECT 0.065 130.920 449.815 132.240 ;
        RECT 4.400 129.560 449.815 130.920 ;
        RECT 4.400 129.520 445.600 129.560 ;
        RECT 0.065 128.160 445.600 129.520 ;
        RECT 0.065 126.160 449.815 128.160 ;
        RECT 4.400 124.800 449.815 126.160 ;
        RECT 4.400 124.760 445.600 124.800 ;
        RECT 0.065 123.400 445.600 124.760 ;
        RECT 0.065 121.400 449.815 123.400 ;
        RECT 4.400 120.720 449.815 121.400 ;
        RECT 4.400 120.000 445.600 120.720 ;
        RECT 0.065 119.320 445.600 120.000 ;
        RECT 0.065 117.320 449.815 119.320 ;
        RECT 4.400 116.640 449.815 117.320 ;
        RECT 4.400 115.920 445.600 116.640 ;
        RECT 0.065 115.240 445.600 115.920 ;
        RECT 0.065 112.560 449.815 115.240 ;
        RECT 4.400 111.880 449.815 112.560 ;
        RECT 4.400 111.160 445.600 111.880 ;
        RECT 0.065 110.480 445.600 111.160 ;
        RECT 0.065 107.800 449.815 110.480 ;
        RECT 4.400 106.400 445.600 107.800 ;
        RECT 0.065 103.040 449.815 106.400 ;
        RECT 4.400 101.640 445.600 103.040 ;
        RECT 0.065 98.960 449.815 101.640 ;
        RECT 4.400 97.560 445.600 98.960 ;
        RECT 0.065 94.200 449.815 97.560 ;
        RECT 4.400 92.800 445.600 94.200 ;
        RECT 0.065 90.120 449.815 92.800 ;
        RECT 0.065 89.440 445.600 90.120 ;
        RECT 4.400 88.720 445.600 89.440 ;
        RECT 4.400 88.040 449.815 88.720 ;
        RECT 0.065 86.040 449.815 88.040 ;
        RECT 0.065 84.680 445.600 86.040 ;
        RECT 4.400 84.640 445.600 84.680 ;
        RECT 4.400 83.280 449.815 84.640 ;
        RECT 0.065 81.280 449.815 83.280 ;
        RECT 0.065 80.600 445.600 81.280 ;
        RECT 4.400 79.880 445.600 80.600 ;
        RECT 4.400 79.200 449.815 79.880 ;
        RECT 0.065 77.200 449.815 79.200 ;
        RECT 0.065 75.840 445.600 77.200 ;
        RECT 4.400 75.800 445.600 75.840 ;
        RECT 4.400 74.440 449.815 75.800 ;
        RECT 0.065 72.440 449.815 74.440 ;
        RECT 0.065 71.080 445.600 72.440 ;
        RECT 4.400 71.040 445.600 71.080 ;
        RECT 4.400 69.680 449.815 71.040 ;
        RECT 0.065 68.360 449.815 69.680 ;
        RECT 0.065 67.000 445.600 68.360 ;
        RECT 4.400 66.960 445.600 67.000 ;
        RECT 4.400 65.600 449.815 66.960 ;
        RECT 0.065 63.600 449.815 65.600 ;
        RECT 0.065 62.240 445.600 63.600 ;
        RECT 4.400 62.200 445.600 62.240 ;
        RECT 4.400 60.840 449.815 62.200 ;
        RECT 0.065 59.520 449.815 60.840 ;
        RECT 0.065 58.120 445.600 59.520 ;
        RECT 0.065 57.480 449.815 58.120 ;
        RECT 4.400 56.080 449.815 57.480 ;
        RECT 0.065 55.440 449.815 56.080 ;
        RECT 0.065 54.040 445.600 55.440 ;
        RECT 0.065 52.720 449.815 54.040 ;
        RECT 4.400 51.320 449.815 52.720 ;
        RECT 0.065 50.680 449.815 51.320 ;
        RECT 0.065 49.280 445.600 50.680 ;
        RECT 0.065 48.640 449.815 49.280 ;
        RECT 4.400 47.240 449.815 48.640 ;
        RECT 0.065 46.600 449.815 47.240 ;
        RECT 0.065 45.200 445.600 46.600 ;
        RECT 0.065 43.880 449.815 45.200 ;
        RECT 4.400 42.480 449.815 43.880 ;
        RECT 0.065 41.840 449.815 42.480 ;
        RECT 0.065 40.440 445.600 41.840 ;
        RECT 0.065 39.120 449.815 40.440 ;
        RECT 4.400 37.760 449.815 39.120 ;
        RECT 4.400 37.720 445.600 37.760 ;
        RECT 0.065 36.360 445.600 37.720 ;
        RECT 0.065 35.040 449.815 36.360 ;
        RECT 4.400 33.640 449.815 35.040 ;
        RECT 0.065 33.000 449.815 33.640 ;
        RECT 0.065 31.600 445.600 33.000 ;
        RECT 0.065 30.280 449.815 31.600 ;
        RECT 4.400 28.920 449.815 30.280 ;
        RECT 4.400 28.880 445.600 28.920 ;
        RECT 0.065 27.520 445.600 28.880 ;
        RECT 0.065 25.520 449.815 27.520 ;
        RECT 4.400 24.840 449.815 25.520 ;
        RECT 4.400 24.120 445.600 24.840 ;
        RECT 0.065 23.440 445.600 24.120 ;
        RECT 0.065 20.760 449.815 23.440 ;
        RECT 4.400 20.080 449.815 20.760 ;
        RECT 4.400 19.360 445.600 20.080 ;
        RECT 0.065 18.680 445.600 19.360 ;
        RECT 0.065 16.680 449.815 18.680 ;
        RECT 4.400 16.000 449.815 16.680 ;
        RECT 4.400 15.280 445.600 16.000 ;
        RECT 0.065 14.600 445.600 15.280 ;
        RECT 0.065 11.920 449.815 14.600 ;
        RECT 4.400 11.240 449.815 11.920 ;
        RECT 4.400 10.520 445.600 11.240 ;
        RECT 0.065 9.840 445.600 10.520 ;
        RECT 0.065 7.160 449.815 9.840 ;
        RECT 4.400 5.760 445.600 7.160 ;
        RECT 0.065 3.080 449.815 5.760 ;
        RECT 4.400 2.215 445.600 3.080 ;
      LAYER met4 ;
        RECT 0.295 12.415 20.640 883.825 ;
        RECT 23.040 12.415 97.440 883.825 ;
        RECT 99.840 12.415 174.240 883.825 ;
        RECT 176.640 12.415 251.040 883.825 ;
        RECT 253.440 12.415 327.840 883.825 ;
        RECT 330.240 12.415 404.640 883.825 ;
        RECT 407.040 12.415 449.585 883.825 ;
  END
END ExperiarCore
END LIBRARY

