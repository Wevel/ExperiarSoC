VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ExperiarCore
  CLASS BLOCK ;
  FOREIGN ExperiarCore ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 500.000 ;
  PIN addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 496.000 27.970 500.000 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 496.000 32.110 500.000 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 496.000 36.250 500.000 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 496.000 40.850 500.000 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 496.000 44.990 500.000 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 496.000 49.130 500.000 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 496.000 53.730 500.000 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 496.000 57.870 500.000 ;
    END
  END addr0[7]
  PIN addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 496.000 62.010 500.000 ;
    END
  END addr0[8]
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 496.000 483.830 500.000 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 496.000 487.970 500.000 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 496.000 492.110 500.000 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 496.000 496.710 500.000 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 496.000 500.850 500.000 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 496.000 504.990 500.000 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 496.000 509.590 500.000 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 496.000 513.730 500.000 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 496.000 517.870 500.000 ;
    END
  END addr1[8]
  PIN clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 496.000 2.210 500.000 ;
    END
  END clk0
  PIN clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 496.000 479.230 500.000 ;
    END
  END clk1
  PIN coreIndex[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END coreIndex[0]
  PIN coreIndex[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END coreIndex[1]
  PIN coreIndex[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END coreIndex[2]
  PIN coreIndex[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END coreIndex[3]
  PIN coreIndex[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END coreIndex[4]
  PIN coreIndex[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END coreIndex[5]
  PIN coreIndex[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END coreIndex[6]
  PIN coreIndex[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END coreIndex[7]
  PIN core_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 5.480 800.000 6.080 ;
    END
  END core_wb_ack_i
  PIN core_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 19.760 800.000 20.360 ;
    END
  END core_wb_adr_o[0]
  PIN core_wb_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 102.040 800.000 102.640 ;
    END
  END core_wb_adr_o[10]
  PIN core_wb_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 108.840 800.000 109.440 ;
    END
  END core_wb_adr_o[11]
  PIN core_wb_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 116.320 800.000 116.920 ;
    END
  END core_wb_adr_o[12]
  PIN core_wb_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 123.800 800.000 124.400 ;
    END
  END core_wb_adr_o[13]
  PIN core_wb_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 130.600 800.000 131.200 ;
    END
  END core_wb_adr_o[14]
  PIN core_wb_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 138.080 800.000 138.680 ;
    END
  END core_wb_adr_o[15]
  PIN core_wb_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 145.560 800.000 146.160 ;
    END
  END core_wb_adr_o[16]
  PIN core_wb_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 152.360 800.000 152.960 ;
    END
  END core_wb_adr_o[17]
  PIN core_wb_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 159.840 800.000 160.440 ;
    END
  END core_wb_adr_o[18]
  PIN core_wb_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 167.320 800.000 167.920 ;
    END
  END core_wb_adr_o[19]
  PIN core_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 29.280 800.000 29.880 ;
    END
  END core_wb_adr_o[1]
  PIN core_wb_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 174.120 800.000 174.720 ;
    END
  END core_wb_adr_o[20]
  PIN core_wb_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 181.600 800.000 182.200 ;
    END
  END core_wb_adr_o[21]
  PIN core_wb_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 188.400 800.000 189.000 ;
    END
  END core_wb_adr_o[22]
  PIN core_wb_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 195.880 800.000 196.480 ;
    END
  END core_wb_adr_o[23]
  PIN core_wb_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 203.360 800.000 203.960 ;
    END
  END core_wb_adr_o[24]
  PIN core_wb_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 210.160 800.000 210.760 ;
    END
  END core_wb_adr_o[25]
  PIN core_wb_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 217.640 800.000 218.240 ;
    END
  END core_wb_adr_o[26]
  PIN core_wb_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 225.120 800.000 225.720 ;
    END
  END core_wb_adr_o[27]
  PIN core_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 38.800 800.000 39.400 ;
    END
  END core_wb_adr_o[2]
  PIN core_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 49.000 800.000 49.600 ;
    END
  END core_wb_adr_o[3]
  PIN core_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 58.520 800.000 59.120 ;
    END
  END core_wb_adr_o[4]
  PIN core_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 65.320 800.000 65.920 ;
    END
  END core_wb_adr_o[5]
  PIN core_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 72.800 800.000 73.400 ;
    END
  END core_wb_adr_o[6]
  PIN core_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 80.280 800.000 80.880 ;
    END
  END core_wb_adr_o[7]
  PIN core_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 87.080 800.000 87.680 ;
    END
  END core_wb_adr_o[8]
  PIN core_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 94.560 800.000 95.160 ;
    END
  END core_wb_adr_o[9]
  PIN core_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 7.520 800.000 8.120 ;
    END
  END core_wb_cyc_o
  PIN core_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 21.800 800.000 22.400 ;
    END
  END core_wb_data_i[0]
  PIN core_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 104.080 800.000 104.680 ;
    END
  END core_wb_data_i[10]
  PIN core_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 111.560 800.000 112.160 ;
    END
  END core_wb_data_i[11]
  PIN core_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 118.360 800.000 118.960 ;
    END
  END core_wb_data_i[12]
  PIN core_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 125.840 800.000 126.440 ;
    END
  END core_wb_data_i[13]
  PIN core_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 133.320 800.000 133.920 ;
    END
  END core_wb_data_i[14]
  PIN core_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 140.120 800.000 140.720 ;
    END
  END core_wb_data_i[15]
  PIN core_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 147.600 800.000 148.200 ;
    END
  END core_wb_data_i[16]
  PIN core_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 155.080 800.000 155.680 ;
    END
  END core_wb_data_i[17]
  PIN core_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 161.880 800.000 162.480 ;
    END
  END core_wb_data_i[18]
  PIN core_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 169.360 800.000 169.960 ;
    END
  END core_wb_data_i[19]
  PIN core_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 32.000 800.000 32.600 ;
    END
  END core_wb_data_i[1]
  PIN core_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 176.840 800.000 177.440 ;
    END
  END core_wb_data_i[20]
  PIN core_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 183.640 800.000 184.240 ;
    END
  END core_wb_data_i[21]
  PIN core_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 191.120 800.000 191.720 ;
    END
  END core_wb_data_i[22]
  PIN core_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 198.600 800.000 199.200 ;
    END
  END core_wb_data_i[23]
  PIN core_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 205.400 800.000 206.000 ;
    END
  END core_wb_data_i[24]
  PIN core_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 212.880 800.000 213.480 ;
    END
  END core_wb_data_i[25]
  PIN core_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 220.360 800.000 220.960 ;
    END
  END core_wb_data_i[26]
  PIN core_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 227.160 800.000 227.760 ;
    END
  END core_wb_data_i[27]
  PIN core_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 231.920 800.000 232.520 ;
    END
  END core_wb_data_i[28]
  PIN core_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 236.680 800.000 237.280 ;
    END
  END core_wb_data_i[29]
  PIN core_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 41.520 800.000 42.120 ;
    END
  END core_wb_data_i[2]
  PIN core_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 242.120 800.000 242.720 ;
    END
  END core_wb_data_i[30]
  PIN core_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 246.880 800.000 247.480 ;
    END
  END core_wb_data_i[31]
  PIN core_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 51.040 800.000 51.640 ;
    END
  END core_wb_data_i[3]
  PIN core_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 60.560 800.000 61.160 ;
    END
  END core_wb_data_i[4]
  PIN core_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 68.040 800.000 68.640 ;
    END
  END core_wb_data_i[5]
  PIN core_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 75.520 800.000 76.120 ;
    END
  END core_wb_data_i[6]
  PIN core_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 82.320 800.000 82.920 ;
    END
  END core_wb_data_i[7]
  PIN core_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 89.800 800.000 90.400 ;
    END
  END core_wb_data_i[8]
  PIN core_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 97.280 800.000 97.880 ;
    END
  END core_wb_data_i[9]
  PIN core_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 24.520 800.000 25.120 ;
    END
  END core_wb_data_o[0]
  PIN core_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 106.800 800.000 107.400 ;
    END
  END core_wb_data_o[10]
  PIN core_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 113.600 800.000 114.200 ;
    END
  END core_wb_data_o[11]
  PIN core_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 121.080 800.000 121.680 ;
    END
  END core_wb_data_o[12]
  PIN core_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 128.560 800.000 129.160 ;
    END
  END core_wb_data_o[13]
  PIN core_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 135.360 800.000 135.960 ;
    END
  END core_wb_data_o[14]
  PIN core_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 142.840 800.000 143.440 ;
    END
  END core_wb_data_o[15]
  PIN core_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 150.320 800.000 150.920 ;
    END
  END core_wb_data_o[16]
  PIN core_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 157.120 800.000 157.720 ;
    END
  END core_wb_data_o[17]
  PIN core_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 164.600 800.000 165.200 ;
    END
  END core_wb_data_o[18]
  PIN core_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 172.080 800.000 172.680 ;
    END
  END core_wb_data_o[19]
  PIN core_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 34.040 800.000 34.640 ;
    END
  END core_wb_data_o[1]
  PIN core_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 178.880 800.000 179.480 ;
    END
  END core_wb_data_o[20]
  PIN core_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 186.360 800.000 186.960 ;
    END
  END core_wb_data_o[21]
  PIN core_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 193.840 800.000 194.440 ;
    END
  END core_wb_data_o[22]
  PIN core_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 200.640 800.000 201.240 ;
    END
  END core_wb_data_o[23]
  PIN core_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 208.120 800.000 208.720 ;
    END
  END core_wb_data_o[24]
  PIN core_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 215.600 800.000 216.200 ;
    END
  END core_wb_data_o[25]
  PIN core_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 222.400 800.000 223.000 ;
    END
  END core_wb_data_o[26]
  PIN core_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 229.880 800.000 230.480 ;
    END
  END core_wb_data_o[27]
  PIN core_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 234.640 800.000 235.240 ;
    END
  END core_wb_data_o[28]
  PIN core_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 239.400 800.000 240.000 ;
    END
  END core_wb_data_o[29]
  PIN core_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 43.560 800.000 44.160 ;
    END
  END core_wb_data_o[2]
  PIN core_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 244.160 800.000 244.760 ;
    END
  END core_wb_data_o[30]
  PIN core_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 248.920 800.000 249.520 ;
    END
  END core_wb_data_o[31]
  PIN core_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 53.760 800.000 54.360 ;
    END
  END core_wb_data_o[3]
  PIN core_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 63.280 800.000 63.880 ;
    END
  END core_wb_data_o[4]
  PIN core_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 70.080 800.000 70.680 ;
    END
  END core_wb_data_o[5]
  PIN core_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 77.560 800.000 78.160 ;
    END
  END core_wb_data_o[6]
  PIN core_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 85.040 800.000 85.640 ;
    END
  END core_wb_data_o[7]
  PIN core_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 91.840 800.000 92.440 ;
    END
  END core_wb_data_o[8]
  PIN core_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 99.320 800.000 99.920 ;
    END
  END core_wb_data_o[9]
  PIN core_wb_error_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 10.240 800.000 10.840 ;
    END
  END core_wb_error_i
  PIN core_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 27.240 800.000 27.840 ;
    END
  END core_wb_sel_o[0]
  PIN core_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 36.760 800.000 37.360 ;
    END
  END core_wb_sel_o[1]
  PIN core_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 46.280 800.000 46.880 ;
    END
  END core_wb_sel_o[2]
  PIN core_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 55.800 800.000 56.400 ;
    END
  END core_wb_sel_o[3]
  PIN core_wb_stall_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 12.280 800.000 12.880 ;
    END
  END core_wb_stall_i
  PIN core_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 15.000 800.000 15.600 ;
    END
  END core_wb_stb_o
  PIN core_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 17.040 800.000 17.640 ;
    END
  END core_wb_we_o
  PIN csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 493.040 800.000 493.640 ;
    END
  END csb0[0]
  PIN csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 495.080 800.000 495.680 ;
    END
  END csb0[1]
  PIN csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 494.400 4.000 495.000 ;
    END
  END csb1[0]
  PIN csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 497.800 800.000 498.400 ;
    END
  END csb1[1]
  PIN din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 496.000 66.610 500.000 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 496.000 109.390 500.000 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 496.000 113.990 500.000 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 496.000 118.130 500.000 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 496.000 122.270 500.000 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 496.000 126.870 500.000 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 496.000 131.010 500.000 ;
    END
  END din0[15]
  PIN din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 496.000 135.150 500.000 ;
    END
  END din0[16]
  PIN din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 496.000 139.750 500.000 ;
    END
  END din0[17]
  PIN din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 496.000 143.890 500.000 ;
    END
  END din0[18]
  PIN din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 496.000 148.030 500.000 ;
    END
  END din0[19]
  PIN din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 496.000 70.750 500.000 ;
    END
  END din0[1]
  PIN din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 496.000 152.630 500.000 ;
    END
  END din0[20]
  PIN din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 496.000 156.770 500.000 ;
    END
  END din0[21]
  PIN din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 496.000 160.910 500.000 ;
    END
  END din0[22]
  PIN din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 496.000 165.510 500.000 ;
    END
  END din0[23]
  PIN din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 496.000 169.650 500.000 ;
    END
  END din0[24]
  PIN din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 496.000 173.790 500.000 ;
    END
  END din0[25]
  PIN din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 496.000 178.390 500.000 ;
    END
  END din0[26]
  PIN din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 496.000 182.530 500.000 ;
    END
  END din0[27]
  PIN din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 496.000 187.130 500.000 ;
    END
  END din0[28]
  PIN din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 496.000 191.270 500.000 ;
    END
  END din0[29]
  PIN din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 496.000 74.890 500.000 ;
    END
  END din0[2]
  PIN din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 496.000 195.410 500.000 ;
    END
  END din0[30]
  PIN din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 496.000 200.010 500.000 ;
    END
  END din0[31]
  PIN din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 496.000 79.490 500.000 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 496.000 83.630 500.000 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 496.000 87.770 500.000 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 496.000 92.370 500.000 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 496.000 96.510 500.000 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 496.000 101.110 500.000 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 496.000 105.250 500.000 ;
    END
  END din0[9]
  PIN dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 496.000 204.150 500.000 ;
    END
  END dout0[0]
  PIN dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 496.000 246.930 500.000 ;
    END
  END dout0[10]
  PIN dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 496.000 251.530 500.000 ;
    END
  END dout0[11]
  PIN dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 496.000 255.670 500.000 ;
    END
  END dout0[12]
  PIN dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 496.000 259.810 500.000 ;
    END
  END dout0[13]
  PIN dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 496.000 264.410 500.000 ;
    END
  END dout0[14]
  PIN dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 496.000 268.550 500.000 ;
    END
  END dout0[15]
  PIN dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 496.000 273.150 500.000 ;
    END
  END dout0[16]
  PIN dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 496.000 277.290 500.000 ;
    END
  END dout0[17]
  PIN dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 496.000 281.430 500.000 ;
    END
  END dout0[18]
  PIN dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 496.000 286.030 500.000 ;
    END
  END dout0[19]
  PIN dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 496.000 208.290 500.000 ;
    END
  END dout0[1]
  PIN dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 496.000 290.170 500.000 ;
    END
  END dout0[20]
  PIN dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 496.000 294.310 500.000 ;
    END
  END dout0[21]
  PIN dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 496.000 298.910 500.000 ;
    END
  END dout0[22]
  PIN dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 496.000 303.050 500.000 ;
    END
  END dout0[23]
  PIN dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 496.000 307.190 500.000 ;
    END
  END dout0[24]
  PIN dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 496.000 311.790 500.000 ;
    END
  END dout0[25]
  PIN dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 496.000 315.930 500.000 ;
    END
  END dout0[26]
  PIN dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 496.000 320.070 500.000 ;
    END
  END dout0[27]
  PIN dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 496.000 324.670 500.000 ;
    END
  END dout0[28]
  PIN dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 496.000 328.810 500.000 ;
    END
  END dout0[29]
  PIN dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 496.000 212.890 500.000 ;
    END
  END dout0[2]
  PIN dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 496.000 332.950 500.000 ;
    END
  END dout0[30]
  PIN dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 496.000 337.550 500.000 ;
    END
  END dout0[31]
  PIN dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 496.000 341.690 500.000 ;
    END
  END dout0[32]
  PIN dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 496.000 345.830 500.000 ;
    END
  END dout0[33]
  PIN dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 496.000 350.430 500.000 ;
    END
  END dout0[34]
  PIN dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 496.000 354.570 500.000 ;
    END
  END dout0[35]
  PIN dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 496.000 359.170 500.000 ;
    END
  END dout0[36]
  PIN dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 496.000 363.310 500.000 ;
    END
  END dout0[37]
  PIN dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 496.000 367.450 500.000 ;
    END
  END dout0[38]
  PIN dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 496.000 372.050 500.000 ;
    END
  END dout0[39]
  PIN dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 496.000 217.030 500.000 ;
    END
  END dout0[3]
  PIN dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 496.000 376.190 500.000 ;
    END
  END dout0[40]
  PIN dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 496.000 380.330 500.000 ;
    END
  END dout0[41]
  PIN dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 496.000 384.930 500.000 ;
    END
  END dout0[42]
  PIN dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 496.000 389.070 500.000 ;
    END
  END dout0[43]
  PIN dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 496.000 393.210 500.000 ;
    END
  END dout0[44]
  PIN dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 496.000 397.810 500.000 ;
    END
  END dout0[45]
  PIN dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 496.000 401.950 500.000 ;
    END
  END dout0[46]
  PIN dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 496.000 406.090 500.000 ;
    END
  END dout0[47]
  PIN dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 496.000 410.690 500.000 ;
    END
  END dout0[48]
  PIN dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 496.000 414.830 500.000 ;
    END
  END dout0[49]
  PIN dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 496.000 221.170 500.000 ;
    END
  END dout0[4]
  PIN dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 496.000 418.970 500.000 ;
    END
  END dout0[50]
  PIN dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 496.000 423.570 500.000 ;
    END
  END dout0[51]
  PIN dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 496.000 427.710 500.000 ;
    END
  END dout0[52]
  PIN dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 496.000 431.850 500.000 ;
    END
  END dout0[53]
  PIN dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 496.000 436.450 500.000 ;
    END
  END dout0[54]
  PIN dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 496.000 440.590 500.000 ;
    END
  END dout0[55]
  PIN dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 496.000 444.730 500.000 ;
    END
  END dout0[56]
  PIN dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 496.000 449.330 500.000 ;
    END
  END dout0[57]
  PIN dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 496.000 453.470 500.000 ;
    END
  END dout0[58]
  PIN dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 496.000 458.070 500.000 ;
    END
  END dout0[59]
  PIN dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 496.000 225.770 500.000 ;
    END
  END dout0[5]
  PIN dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 496.000 462.210 500.000 ;
    END
  END dout0[60]
  PIN dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 496.000 466.350 500.000 ;
    END
  END dout0[61]
  PIN dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 496.000 470.950 500.000 ;
    END
  END dout0[62]
  PIN dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 496.000 475.090 500.000 ;
    END
  END dout0[63]
  PIN dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 496.000 229.910 500.000 ;
    END
  END dout0[6]
  PIN dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 496.000 234.050 500.000 ;
    END
  END dout0[7]
  PIN dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 496.000 238.650 500.000 ;
    END
  END dout0[8]
  PIN dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 496.000 242.790 500.000 ;
    END
  END dout0[9]
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 496.000 522.470 500.000 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 496.000 565.250 500.000 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 496.000 569.850 500.000 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 496.000 573.990 500.000 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 496.000 578.130 500.000 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 496.000 582.730 500.000 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 496.000 586.870 500.000 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 496.000 591.010 500.000 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 496.000 595.610 500.000 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 496.000 599.750 500.000 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 496.000 603.890 500.000 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 496.000 526.610 500.000 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 496.000 608.490 500.000 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 496.000 612.630 500.000 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 496.000 616.770 500.000 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 496.000 621.370 500.000 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 496.000 625.510 500.000 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 496.000 630.110 500.000 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 496.000 634.250 500.000 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.110 496.000 638.390 500.000 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 496.000 642.990 500.000 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 496.000 647.130 500.000 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 496.000 530.750 500.000 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 496.000 651.270 500.000 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 496.000 655.870 500.000 ;
    END
  END dout1[31]
  PIN dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 496.000 660.010 500.000 ;
    END
  END dout1[32]
  PIN dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 496.000 664.150 500.000 ;
    END
  END dout1[33]
  PIN dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 496.000 668.750 500.000 ;
    END
  END dout1[34]
  PIN dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 496.000 672.890 500.000 ;
    END
  END dout1[35]
  PIN dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 496.000 677.030 500.000 ;
    END
  END dout1[36]
  PIN dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 496.000 681.630 500.000 ;
    END
  END dout1[37]
  PIN dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 496.000 685.770 500.000 ;
    END
  END dout1[38]
  PIN dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 496.000 689.910 500.000 ;
    END
  END dout1[39]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 496.000 535.350 500.000 ;
    END
  END dout1[3]
  PIN dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 496.000 694.510 500.000 ;
    END
  END dout1[40]
  PIN dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 496.000 698.650 500.000 ;
    END
  END dout1[41]
  PIN dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 496.000 702.790 500.000 ;
    END
  END dout1[42]
  PIN dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 496.000 707.390 500.000 ;
    END
  END dout1[43]
  PIN dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 496.000 711.530 500.000 ;
    END
  END dout1[44]
  PIN dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 496.000 716.130 500.000 ;
    END
  END dout1[45]
  PIN dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 496.000 720.270 500.000 ;
    END
  END dout1[46]
  PIN dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 496.000 724.410 500.000 ;
    END
  END dout1[47]
  PIN dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 496.000 729.010 500.000 ;
    END
  END dout1[48]
  PIN dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 496.000 733.150 500.000 ;
    END
  END dout1[49]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 496.000 539.490 500.000 ;
    END
  END dout1[4]
  PIN dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 496.000 737.290 500.000 ;
    END
  END dout1[50]
  PIN dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 496.000 741.890 500.000 ;
    END
  END dout1[51]
  PIN dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 496.000 746.030 500.000 ;
    END
  END dout1[52]
  PIN dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 496.000 750.170 500.000 ;
    END
  END dout1[53]
  PIN dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 496.000 754.770 500.000 ;
    END
  END dout1[54]
  PIN dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.630 496.000 758.910 500.000 ;
    END
  END dout1[55]
  PIN dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 496.000 763.050 500.000 ;
    END
  END dout1[56]
  PIN dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 496.000 767.650 500.000 ;
    END
  END dout1[57]
  PIN dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 496.000 771.790 500.000 ;
    END
  END dout1[58]
  PIN dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 496.000 775.930 500.000 ;
    END
  END dout1[59]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 496.000 544.090 500.000 ;
    END
  END dout1[5]
  PIN dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 496.000 780.530 500.000 ;
    END
  END dout1[60]
  PIN dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 496.000 784.670 500.000 ;
    END
  END dout1[61]
  PIN dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.530 496.000 788.810 500.000 ;
    END
  END dout1[62]
  PIN dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 496.000 793.410 500.000 ;
    END
  END dout1[63]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 496.000 548.230 500.000 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 496.000 552.370 500.000 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 496.000 556.970 500.000 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 496.000 561.110 500.000 ;
    END
  END dout1[9]
  PIN jtag_tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END jtag_tck
  PIN jtag_tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 496.000 797.550 500.000 ;
    END
  END jtag_tdi
  PIN jtag_tdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 488.280 800.000 488.880 ;
    END
  END jtag_tdo
  PIN jtag_tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 490.320 800.000 490.920 ;
    END
  END jtag_tms
  PIN localMemory_wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 251.640 800.000 252.240 ;
    END
  END localMemory_wb_ack_o
  PIN localMemory_wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 265.920 800.000 266.520 ;
    END
  END localMemory_wb_adr_i[0]
  PIN localMemory_wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 348.200 800.000 348.800 ;
    END
  END localMemory_wb_adr_i[10]
  PIN localMemory_wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 355.000 800.000 355.600 ;
    END
  END localMemory_wb_adr_i[11]
  PIN localMemory_wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 362.480 800.000 363.080 ;
    END
  END localMemory_wb_adr_i[12]
  PIN localMemory_wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 369.960 800.000 370.560 ;
    END
  END localMemory_wb_adr_i[13]
  PIN localMemory_wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 376.760 800.000 377.360 ;
    END
  END localMemory_wb_adr_i[14]
  PIN localMemory_wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 384.240 800.000 384.840 ;
    END
  END localMemory_wb_adr_i[15]
  PIN localMemory_wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 391.720 800.000 392.320 ;
    END
  END localMemory_wb_adr_i[16]
  PIN localMemory_wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 398.520 800.000 399.120 ;
    END
  END localMemory_wb_adr_i[17]
  PIN localMemory_wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 406.000 800.000 406.600 ;
    END
  END localMemory_wb_adr_i[18]
  PIN localMemory_wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 413.480 800.000 414.080 ;
    END
  END localMemory_wb_adr_i[19]
  PIN localMemory_wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 275.440 800.000 276.040 ;
    END
  END localMemory_wb_adr_i[1]
  PIN localMemory_wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 420.280 800.000 420.880 ;
    END
  END localMemory_wb_adr_i[20]
  PIN localMemory_wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 427.760 800.000 428.360 ;
    END
  END localMemory_wb_adr_i[21]
  PIN localMemory_wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 435.240 800.000 435.840 ;
    END
  END localMemory_wb_adr_i[22]
  PIN localMemory_wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 442.040 800.000 442.640 ;
    END
  END localMemory_wb_adr_i[23]
  PIN localMemory_wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 284.960 800.000 285.560 ;
    END
  END localMemory_wb_adr_i[2]
  PIN localMemory_wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 295.160 800.000 295.760 ;
    END
  END localMemory_wb_adr_i[3]
  PIN localMemory_wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 304.680 800.000 305.280 ;
    END
  END localMemory_wb_adr_i[4]
  PIN localMemory_wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 312.160 800.000 312.760 ;
    END
  END localMemory_wb_adr_i[5]
  PIN localMemory_wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 318.960 800.000 319.560 ;
    END
  END localMemory_wb_adr_i[6]
  PIN localMemory_wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 326.440 800.000 327.040 ;
    END
  END localMemory_wb_adr_i[7]
  PIN localMemory_wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 333.920 800.000 334.520 ;
    END
  END localMemory_wb_adr_i[8]
  PIN localMemory_wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 340.720 800.000 341.320 ;
    END
  END localMemory_wb_adr_i[9]
  PIN localMemory_wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 253.680 800.000 254.280 ;
    END
  END localMemory_wb_cyc_i
  PIN localMemory_wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 268.640 800.000 269.240 ;
    END
  END localMemory_wb_data_i[0]
  PIN localMemory_wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 350.240 800.000 350.840 ;
    END
  END localMemory_wb_data_i[10]
  PIN localMemory_wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 357.720 800.000 358.320 ;
    END
  END localMemory_wb_data_i[11]
  PIN localMemory_wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 365.200 800.000 365.800 ;
    END
  END localMemory_wb_data_i[12]
  PIN localMemory_wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 372.000 800.000 372.600 ;
    END
  END localMemory_wb_data_i[13]
  PIN localMemory_wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 379.480 800.000 380.080 ;
    END
  END localMemory_wb_data_i[14]
  PIN localMemory_wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 386.960 800.000 387.560 ;
    END
  END localMemory_wb_data_i[15]
  PIN localMemory_wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 393.760 800.000 394.360 ;
    END
  END localMemory_wb_data_i[16]
  PIN localMemory_wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 401.240 800.000 401.840 ;
    END
  END localMemory_wb_data_i[17]
  PIN localMemory_wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 408.720 800.000 409.320 ;
    END
  END localMemory_wb_data_i[18]
  PIN localMemory_wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 415.520 800.000 416.120 ;
    END
  END localMemory_wb_data_i[19]
  PIN localMemory_wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 278.160 800.000 278.760 ;
    END
  END localMemory_wb_data_i[1]
  PIN localMemory_wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 423.000 800.000 423.600 ;
    END
  END localMemory_wb_data_i[20]
  PIN localMemory_wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 430.480 800.000 431.080 ;
    END
  END localMemory_wb_data_i[21]
  PIN localMemory_wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 437.280 800.000 437.880 ;
    END
  END localMemory_wb_data_i[22]
  PIN localMemory_wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 444.760 800.000 445.360 ;
    END
  END localMemory_wb_data_i[23]
  PIN localMemory_wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 449.520 800.000 450.120 ;
    END
  END localMemory_wb_data_i[24]
  PIN localMemory_wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 454.280 800.000 454.880 ;
    END
  END localMemory_wb_data_i[25]
  PIN localMemory_wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 459.040 800.000 459.640 ;
    END
  END localMemory_wb_data_i[26]
  PIN localMemory_wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 463.800 800.000 464.400 ;
    END
  END localMemory_wb_data_i[27]
  PIN localMemory_wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 468.560 800.000 469.160 ;
    END
  END localMemory_wb_data_i[28]
  PIN localMemory_wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 473.320 800.000 473.920 ;
    END
  END localMemory_wb_data_i[29]
  PIN localMemory_wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 287.680 800.000 288.280 ;
    END
  END localMemory_wb_data_i[2]
  PIN localMemory_wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 478.760 800.000 479.360 ;
    END
  END localMemory_wb_data_i[30]
  PIN localMemory_wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 483.520 800.000 484.120 ;
    END
  END localMemory_wb_data_i[31]
  PIN localMemory_wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 297.200 800.000 297.800 ;
    END
  END localMemory_wb_data_i[3]
  PIN localMemory_wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 306.720 800.000 307.320 ;
    END
  END localMemory_wb_data_i[4]
  PIN localMemory_wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 314.200 800.000 314.800 ;
    END
  END localMemory_wb_data_i[5]
  PIN localMemory_wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 321.680 800.000 322.280 ;
    END
  END localMemory_wb_data_i[6]
  PIN localMemory_wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 328.480 800.000 329.080 ;
    END
  END localMemory_wb_data_i[7]
  PIN localMemory_wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 335.960 800.000 336.560 ;
    END
  END localMemory_wb_data_i[8]
  PIN localMemory_wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 343.440 800.000 344.040 ;
    END
  END localMemory_wb_data_i[9]
  PIN localMemory_wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 270.680 800.000 271.280 ;
    END
  END localMemory_wb_data_o[0]
  PIN localMemory_wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 352.960 800.000 353.560 ;
    END
  END localMemory_wb_data_o[10]
  PIN localMemory_wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 360.440 800.000 361.040 ;
    END
  END localMemory_wb_data_o[11]
  PIN localMemory_wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 367.240 800.000 367.840 ;
    END
  END localMemory_wb_data_o[12]
  PIN localMemory_wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 374.720 800.000 375.320 ;
    END
  END localMemory_wb_data_o[13]
  PIN localMemory_wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 382.200 800.000 382.800 ;
    END
  END localMemory_wb_data_o[14]
  PIN localMemory_wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 389.000 800.000 389.600 ;
    END
  END localMemory_wb_data_o[15]
  PIN localMemory_wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 396.480 800.000 397.080 ;
    END
  END localMemory_wb_data_o[16]
  PIN localMemory_wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 403.280 800.000 403.880 ;
    END
  END localMemory_wb_data_o[17]
  PIN localMemory_wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 410.760 800.000 411.360 ;
    END
  END localMemory_wb_data_o[18]
  PIN localMemory_wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 418.240 800.000 418.840 ;
    END
  END localMemory_wb_data_o[19]
  PIN localMemory_wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 280.200 800.000 280.800 ;
    END
  END localMemory_wb_data_o[1]
  PIN localMemory_wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 425.040 800.000 425.640 ;
    END
  END localMemory_wb_data_o[20]
  PIN localMemory_wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 432.520 800.000 433.120 ;
    END
  END localMemory_wb_data_o[21]
  PIN localMemory_wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 440.000 800.000 440.600 ;
    END
  END localMemory_wb_data_o[22]
  PIN localMemory_wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 446.800 800.000 447.400 ;
    END
  END localMemory_wb_data_o[23]
  PIN localMemory_wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 451.560 800.000 452.160 ;
    END
  END localMemory_wb_data_o[24]
  PIN localMemory_wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 457.000 800.000 457.600 ;
    END
  END localMemory_wb_data_o[25]
  PIN localMemory_wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 461.760 800.000 462.360 ;
    END
  END localMemory_wb_data_o[26]
  PIN localMemory_wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 466.520 800.000 467.120 ;
    END
  END localMemory_wb_data_o[27]
  PIN localMemory_wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 471.280 800.000 471.880 ;
    END
  END localMemory_wb_data_o[28]
  PIN localMemory_wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 476.040 800.000 476.640 ;
    END
  END localMemory_wb_data_o[29]
  PIN localMemory_wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 290.400 800.000 291.000 ;
    END
  END localMemory_wb_data_o[2]
  PIN localMemory_wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 480.800 800.000 481.400 ;
    END
  END localMemory_wb_data_o[30]
  PIN localMemory_wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 485.560 800.000 486.160 ;
    END
  END localMemory_wb_data_o[31]
  PIN localMemory_wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 299.920 800.000 300.520 ;
    END
  END localMemory_wb_data_o[3]
  PIN localMemory_wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 309.440 800.000 310.040 ;
    END
  END localMemory_wb_data_o[4]
  PIN localMemory_wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 316.920 800.000 317.520 ;
    END
  END localMemory_wb_data_o[5]
  PIN localMemory_wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 323.720 800.000 324.320 ;
    END
  END localMemory_wb_data_o[6]
  PIN localMemory_wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 331.200 800.000 331.800 ;
    END
  END localMemory_wb_data_o[7]
  PIN localMemory_wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 338.680 800.000 339.280 ;
    END
  END localMemory_wb_data_o[8]
  PIN localMemory_wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 345.480 800.000 346.080 ;
    END
  END localMemory_wb_data_o[9]
  PIN localMemory_wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 256.400 800.000 257.000 ;
    END
  END localMemory_wb_error_o
  PIN localMemory_wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 273.400 800.000 274.000 ;
    END
  END localMemory_wb_sel_i[0]
  PIN localMemory_wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 282.920 800.000 283.520 ;
    END
  END localMemory_wb_sel_i[1]
  PIN localMemory_wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 292.440 800.000 293.040 ;
    END
  END localMemory_wb_sel_i[2]
  PIN localMemory_wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 301.960 800.000 302.560 ;
    END
  END localMemory_wb_sel_i[3]
  PIN localMemory_wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 258.440 800.000 259.040 ;
    END
  END localMemory_wb_stall_o
  PIN localMemory_wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 261.160 800.000 261.760 ;
    END
  END localMemory_wb_stb_i
  PIN localMemory_wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 263.880 800.000 264.480 ;
    END
  END localMemory_wb_we_i
  PIN manufacturerID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END manufacturerID[0]
  PIN manufacturerID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END manufacturerID[10]
  PIN manufacturerID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END manufacturerID[1]
  PIN manufacturerID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END manufacturerID[2]
  PIN manufacturerID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END manufacturerID[3]
  PIN manufacturerID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END manufacturerID[4]
  PIN manufacturerID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END manufacturerID[5]
  PIN manufacturerID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END manufacturerID[6]
  PIN manufacturerID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END manufacturerID[7]
  PIN manufacturerID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END manufacturerID[8]
  PIN manufacturerID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END manufacturerID[9]
  PIN partID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END partID[0]
  PIN partID[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END partID[10]
  PIN partID[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END partID[11]
  PIN partID[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 0.000 629.650 4.000 ;
    END
  END partID[12]
  PIN partID[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END partID[13]
  PIN partID[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 0.000 669.670 4.000 ;
    END
  END partID[14]
  PIN partID[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END partID[15]
  PIN partID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END partID[1]
  PIN partID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END partID[2]
  PIN partID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END partID[3]
  PIN partID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END partID[4]
  PIN partID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END partID[5]
  PIN partID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END partID[6]
  PIN partID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END partID[7]
  PIN partID[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END partID[8]
  PIN partID[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END partID[9]
  PIN probe_errorCode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END probe_errorCode[0]
  PIN probe_errorCode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END probe_errorCode[1]
  PIN probe_errorCode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END probe_errorCode[2]
  PIN probe_errorCode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END probe_errorCode[3]
  PIN probe_isBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END probe_isBranch
  PIN probe_isCompressed
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END probe_isCompressed
  PIN probe_isLoad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END probe_isLoad
  PIN probe_isStore
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END probe_isStore
  PIN probe_jtagInstruction[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END probe_jtagInstruction[0]
  PIN probe_jtagInstruction[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END probe_jtagInstruction[1]
  PIN probe_jtagInstruction[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END probe_jtagInstruction[2]
  PIN probe_jtagInstruction[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END probe_jtagInstruction[3]
  PIN probe_jtagInstruction[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END probe_jtagInstruction[4]
  PIN probe_opcode[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END probe_opcode[0]
  PIN probe_opcode[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END probe_opcode[1]
  PIN probe_opcode[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END probe_opcode[2]
  PIN probe_opcode[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END probe_opcode[3]
  PIN probe_opcode[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END probe_opcode[4]
  PIN probe_opcode[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END probe_opcode[5]
  PIN probe_opcode[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END probe_opcode[6]
  PIN probe_programCounter[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END probe_programCounter[0]
  PIN probe_programCounter[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END probe_programCounter[10]
  PIN probe_programCounter[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END probe_programCounter[11]
  PIN probe_programCounter[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END probe_programCounter[12]
  PIN probe_programCounter[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END probe_programCounter[13]
  PIN probe_programCounter[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END probe_programCounter[14]
  PIN probe_programCounter[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END probe_programCounter[15]
  PIN probe_programCounter[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END probe_programCounter[16]
  PIN probe_programCounter[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END probe_programCounter[17]
  PIN probe_programCounter[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END probe_programCounter[18]
  PIN probe_programCounter[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END probe_programCounter[19]
  PIN probe_programCounter[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END probe_programCounter[1]
  PIN probe_programCounter[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END probe_programCounter[20]
  PIN probe_programCounter[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END probe_programCounter[21]
  PIN probe_programCounter[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END probe_programCounter[22]
  PIN probe_programCounter[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.160 4.000 414.760 ;
    END
  END probe_programCounter[23]
  PIN probe_programCounter[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END probe_programCounter[24]
  PIN probe_programCounter[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END probe_programCounter[25]
  PIN probe_programCounter[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END probe_programCounter[26]
  PIN probe_programCounter[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END probe_programCounter[27]
  PIN probe_programCounter[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END probe_programCounter[28]
  PIN probe_programCounter[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END probe_programCounter[29]
  PIN probe_programCounter[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END probe_programCounter[2]
  PIN probe_programCounter[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END probe_programCounter[30]
  PIN probe_programCounter[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END probe_programCounter[31]
  PIN probe_programCounter[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END probe_programCounter[3]
  PIN probe_programCounter[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END probe_programCounter[4]
  PIN probe_programCounter[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END probe_programCounter[5]
  PIN probe_programCounter[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END probe_programCounter[6]
  PIN probe_programCounter[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END probe_programCounter[7]
  PIN probe_programCounter[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END probe_programCounter[8]
  PIN probe_programCounter[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END probe_programCounter[9]
  PIN probe_state[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END probe_state[0]
  PIN probe_state[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END probe_state[1]
  PIN probe_takeBranch
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END probe_takeBranch
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 487.120 ;
    END
  END vccd1
  PIN versionID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END versionID[0]
  PIN versionID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END versionID[1]
  PIN versionID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END versionID[2]
  PIN versionID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END versionID[3]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 487.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 0.720 800.000 1.320 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 2.760 800.000 3.360 ;
    END
  END wb_rst_i
  PIN web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 496.000 6.350 500.000 ;
    END
  END web0
  PIN wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 496.000 10.490 500.000 ;
    END
  END wmask0[0]
  PIN wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 496.000 15.090 500.000 ;
    END
  END wmask0[1]
  PIN wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 496.000 19.230 500.000 ;
    END
  END wmask0[2]
  PIN wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 496.000 23.370 500.000 ;
    END
  END wmask0[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 486.965 ;
      LAYER met1 ;
        RECT 1.910 7.860 797.570 490.240 ;
      LAYER met2 ;
        RECT 2.490 495.720 5.790 498.285 ;
        RECT 6.630 495.720 9.930 498.285 ;
        RECT 10.770 495.720 14.530 498.285 ;
        RECT 15.370 495.720 18.670 498.285 ;
        RECT 19.510 495.720 22.810 498.285 ;
        RECT 23.650 495.720 27.410 498.285 ;
        RECT 28.250 495.720 31.550 498.285 ;
        RECT 32.390 495.720 35.690 498.285 ;
        RECT 36.530 495.720 40.290 498.285 ;
        RECT 41.130 495.720 44.430 498.285 ;
        RECT 45.270 495.720 48.570 498.285 ;
        RECT 49.410 495.720 53.170 498.285 ;
        RECT 54.010 495.720 57.310 498.285 ;
        RECT 58.150 495.720 61.450 498.285 ;
        RECT 62.290 495.720 66.050 498.285 ;
        RECT 66.890 495.720 70.190 498.285 ;
        RECT 71.030 495.720 74.330 498.285 ;
        RECT 75.170 495.720 78.930 498.285 ;
        RECT 79.770 495.720 83.070 498.285 ;
        RECT 83.910 495.720 87.210 498.285 ;
        RECT 88.050 495.720 91.810 498.285 ;
        RECT 92.650 495.720 95.950 498.285 ;
        RECT 96.790 495.720 100.550 498.285 ;
        RECT 101.390 495.720 104.690 498.285 ;
        RECT 105.530 495.720 108.830 498.285 ;
        RECT 109.670 495.720 113.430 498.285 ;
        RECT 114.270 495.720 117.570 498.285 ;
        RECT 118.410 495.720 121.710 498.285 ;
        RECT 122.550 495.720 126.310 498.285 ;
        RECT 127.150 495.720 130.450 498.285 ;
        RECT 131.290 495.720 134.590 498.285 ;
        RECT 135.430 495.720 139.190 498.285 ;
        RECT 140.030 495.720 143.330 498.285 ;
        RECT 144.170 495.720 147.470 498.285 ;
        RECT 148.310 495.720 152.070 498.285 ;
        RECT 152.910 495.720 156.210 498.285 ;
        RECT 157.050 495.720 160.350 498.285 ;
        RECT 161.190 495.720 164.950 498.285 ;
        RECT 165.790 495.720 169.090 498.285 ;
        RECT 169.930 495.720 173.230 498.285 ;
        RECT 174.070 495.720 177.830 498.285 ;
        RECT 178.670 495.720 181.970 498.285 ;
        RECT 182.810 495.720 186.570 498.285 ;
        RECT 187.410 495.720 190.710 498.285 ;
        RECT 191.550 495.720 194.850 498.285 ;
        RECT 195.690 495.720 199.450 498.285 ;
        RECT 200.290 495.720 203.590 498.285 ;
        RECT 204.430 495.720 207.730 498.285 ;
        RECT 208.570 495.720 212.330 498.285 ;
        RECT 213.170 495.720 216.470 498.285 ;
        RECT 217.310 495.720 220.610 498.285 ;
        RECT 221.450 495.720 225.210 498.285 ;
        RECT 226.050 495.720 229.350 498.285 ;
        RECT 230.190 495.720 233.490 498.285 ;
        RECT 234.330 495.720 238.090 498.285 ;
        RECT 238.930 495.720 242.230 498.285 ;
        RECT 243.070 495.720 246.370 498.285 ;
        RECT 247.210 495.720 250.970 498.285 ;
        RECT 251.810 495.720 255.110 498.285 ;
        RECT 255.950 495.720 259.250 498.285 ;
        RECT 260.090 495.720 263.850 498.285 ;
        RECT 264.690 495.720 267.990 498.285 ;
        RECT 268.830 495.720 272.590 498.285 ;
        RECT 273.430 495.720 276.730 498.285 ;
        RECT 277.570 495.720 280.870 498.285 ;
        RECT 281.710 495.720 285.470 498.285 ;
        RECT 286.310 495.720 289.610 498.285 ;
        RECT 290.450 495.720 293.750 498.285 ;
        RECT 294.590 495.720 298.350 498.285 ;
        RECT 299.190 495.720 302.490 498.285 ;
        RECT 303.330 495.720 306.630 498.285 ;
        RECT 307.470 495.720 311.230 498.285 ;
        RECT 312.070 495.720 315.370 498.285 ;
        RECT 316.210 495.720 319.510 498.285 ;
        RECT 320.350 495.720 324.110 498.285 ;
        RECT 324.950 495.720 328.250 498.285 ;
        RECT 329.090 495.720 332.390 498.285 ;
        RECT 333.230 495.720 336.990 498.285 ;
        RECT 337.830 495.720 341.130 498.285 ;
        RECT 341.970 495.720 345.270 498.285 ;
        RECT 346.110 495.720 349.870 498.285 ;
        RECT 350.710 495.720 354.010 498.285 ;
        RECT 354.850 495.720 358.610 498.285 ;
        RECT 359.450 495.720 362.750 498.285 ;
        RECT 363.590 495.720 366.890 498.285 ;
        RECT 367.730 495.720 371.490 498.285 ;
        RECT 372.330 495.720 375.630 498.285 ;
        RECT 376.470 495.720 379.770 498.285 ;
        RECT 380.610 495.720 384.370 498.285 ;
        RECT 385.210 495.720 388.510 498.285 ;
        RECT 389.350 495.720 392.650 498.285 ;
        RECT 393.490 495.720 397.250 498.285 ;
        RECT 398.090 495.720 401.390 498.285 ;
        RECT 402.230 495.720 405.530 498.285 ;
        RECT 406.370 495.720 410.130 498.285 ;
        RECT 410.970 495.720 414.270 498.285 ;
        RECT 415.110 495.720 418.410 498.285 ;
        RECT 419.250 495.720 423.010 498.285 ;
        RECT 423.850 495.720 427.150 498.285 ;
        RECT 427.990 495.720 431.290 498.285 ;
        RECT 432.130 495.720 435.890 498.285 ;
        RECT 436.730 495.720 440.030 498.285 ;
        RECT 440.870 495.720 444.170 498.285 ;
        RECT 445.010 495.720 448.770 498.285 ;
        RECT 449.610 495.720 452.910 498.285 ;
        RECT 453.750 495.720 457.510 498.285 ;
        RECT 458.350 495.720 461.650 498.285 ;
        RECT 462.490 495.720 465.790 498.285 ;
        RECT 466.630 495.720 470.390 498.285 ;
        RECT 471.230 495.720 474.530 498.285 ;
        RECT 475.370 495.720 478.670 498.285 ;
        RECT 479.510 495.720 483.270 498.285 ;
        RECT 484.110 495.720 487.410 498.285 ;
        RECT 488.250 495.720 491.550 498.285 ;
        RECT 492.390 495.720 496.150 498.285 ;
        RECT 496.990 495.720 500.290 498.285 ;
        RECT 501.130 495.720 504.430 498.285 ;
        RECT 505.270 495.720 509.030 498.285 ;
        RECT 509.870 495.720 513.170 498.285 ;
        RECT 514.010 495.720 517.310 498.285 ;
        RECT 518.150 495.720 521.910 498.285 ;
        RECT 522.750 495.720 526.050 498.285 ;
        RECT 526.890 495.720 530.190 498.285 ;
        RECT 531.030 495.720 534.790 498.285 ;
        RECT 535.630 495.720 538.930 498.285 ;
        RECT 539.770 495.720 543.530 498.285 ;
        RECT 544.370 495.720 547.670 498.285 ;
        RECT 548.510 495.720 551.810 498.285 ;
        RECT 552.650 495.720 556.410 498.285 ;
        RECT 557.250 495.720 560.550 498.285 ;
        RECT 561.390 495.720 564.690 498.285 ;
        RECT 565.530 495.720 569.290 498.285 ;
        RECT 570.130 495.720 573.430 498.285 ;
        RECT 574.270 495.720 577.570 498.285 ;
        RECT 578.410 495.720 582.170 498.285 ;
        RECT 583.010 495.720 586.310 498.285 ;
        RECT 587.150 495.720 590.450 498.285 ;
        RECT 591.290 495.720 595.050 498.285 ;
        RECT 595.890 495.720 599.190 498.285 ;
        RECT 600.030 495.720 603.330 498.285 ;
        RECT 604.170 495.720 607.930 498.285 ;
        RECT 608.770 495.720 612.070 498.285 ;
        RECT 612.910 495.720 616.210 498.285 ;
        RECT 617.050 495.720 620.810 498.285 ;
        RECT 621.650 495.720 624.950 498.285 ;
        RECT 625.790 495.720 629.550 498.285 ;
        RECT 630.390 495.720 633.690 498.285 ;
        RECT 634.530 495.720 637.830 498.285 ;
        RECT 638.670 495.720 642.430 498.285 ;
        RECT 643.270 495.720 646.570 498.285 ;
        RECT 647.410 495.720 650.710 498.285 ;
        RECT 651.550 495.720 655.310 498.285 ;
        RECT 656.150 495.720 659.450 498.285 ;
        RECT 660.290 495.720 663.590 498.285 ;
        RECT 664.430 495.720 668.190 498.285 ;
        RECT 669.030 495.720 672.330 498.285 ;
        RECT 673.170 495.720 676.470 498.285 ;
        RECT 677.310 495.720 681.070 498.285 ;
        RECT 681.910 495.720 685.210 498.285 ;
        RECT 686.050 495.720 689.350 498.285 ;
        RECT 690.190 495.720 693.950 498.285 ;
        RECT 694.790 495.720 698.090 498.285 ;
        RECT 698.930 495.720 702.230 498.285 ;
        RECT 703.070 495.720 706.830 498.285 ;
        RECT 707.670 495.720 710.970 498.285 ;
        RECT 711.810 495.720 715.570 498.285 ;
        RECT 716.410 495.720 719.710 498.285 ;
        RECT 720.550 495.720 723.850 498.285 ;
        RECT 724.690 495.720 728.450 498.285 ;
        RECT 729.290 495.720 732.590 498.285 ;
        RECT 733.430 495.720 736.730 498.285 ;
        RECT 737.570 495.720 741.330 498.285 ;
        RECT 742.170 495.720 745.470 498.285 ;
        RECT 746.310 495.720 749.610 498.285 ;
        RECT 750.450 495.720 754.210 498.285 ;
        RECT 755.050 495.720 758.350 498.285 ;
        RECT 759.190 495.720 762.490 498.285 ;
        RECT 763.330 495.720 767.090 498.285 ;
        RECT 767.930 495.720 771.230 498.285 ;
        RECT 772.070 495.720 775.370 498.285 ;
        RECT 776.210 495.720 779.970 498.285 ;
        RECT 780.810 495.720 784.110 498.285 ;
        RECT 784.950 495.720 788.250 498.285 ;
        RECT 789.090 495.720 792.850 498.285 ;
        RECT 793.690 495.720 796.990 498.285 ;
        RECT 1.940 4.280 797.540 495.720 ;
        RECT 1.940 2.875 9.470 4.280 ;
        RECT 10.310 2.875 29.250 4.280 ;
        RECT 30.090 2.875 49.030 4.280 ;
        RECT 49.870 2.875 69.270 4.280 ;
        RECT 70.110 2.875 89.050 4.280 ;
        RECT 89.890 2.875 109.290 4.280 ;
        RECT 110.130 2.875 129.070 4.280 ;
        RECT 129.910 2.875 149.310 4.280 ;
        RECT 150.150 2.875 169.090 4.280 ;
        RECT 169.930 2.875 189.330 4.280 ;
        RECT 190.170 2.875 209.110 4.280 ;
        RECT 209.950 2.875 229.350 4.280 ;
        RECT 230.190 2.875 249.130 4.280 ;
        RECT 249.970 2.875 269.370 4.280 ;
        RECT 270.210 2.875 289.150 4.280 ;
        RECT 289.990 2.875 309.390 4.280 ;
        RECT 310.230 2.875 329.170 4.280 ;
        RECT 330.010 2.875 349.410 4.280 ;
        RECT 350.250 2.875 369.190 4.280 ;
        RECT 370.030 2.875 389.430 4.280 ;
        RECT 390.270 2.875 409.210 4.280 ;
        RECT 410.050 2.875 428.990 4.280 ;
        RECT 429.830 2.875 449.230 4.280 ;
        RECT 450.070 2.875 469.010 4.280 ;
        RECT 469.850 2.875 489.250 4.280 ;
        RECT 490.090 2.875 509.030 4.280 ;
        RECT 509.870 2.875 529.270 4.280 ;
        RECT 530.110 2.875 549.050 4.280 ;
        RECT 549.890 2.875 569.290 4.280 ;
        RECT 570.130 2.875 589.070 4.280 ;
        RECT 589.910 2.875 609.310 4.280 ;
        RECT 610.150 2.875 629.090 4.280 ;
        RECT 629.930 2.875 649.330 4.280 ;
        RECT 650.170 2.875 669.110 4.280 ;
        RECT 669.950 2.875 689.350 4.280 ;
        RECT 690.190 2.875 709.130 4.280 ;
        RECT 709.970 2.875 729.370 4.280 ;
        RECT 730.210 2.875 749.150 4.280 ;
        RECT 749.990 2.875 769.390 4.280 ;
        RECT 770.230 2.875 789.170 4.280 ;
        RECT 790.010 2.875 797.540 4.280 ;
      LAYER met3 ;
        RECT 4.000 497.400 795.600 498.265 ;
        RECT 4.000 496.080 796.000 497.400 ;
        RECT 4.000 495.400 795.600 496.080 ;
        RECT 4.400 494.680 795.600 495.400 ;
        RECT 4.400 494.040 796.000 494.680 ;
        RECT 4.400 494.000 795.600 494.040 ;
        RECT 4.000 492.640 795.600 494.000 ;
        RECT 4.000 491.320 796.000 492.640 ;
        RECT 4.000 489.920 795.600 491.320 ;
        RECT 4.000 489.280 796.000 489.920 ;
        RECT 4.000 487.880 795.600 489.280 ;
        RECT 4.000 486.560 796.000 487.880 ;
        RECT 4.400 485.160 795.600 486.560 ;
        RECT 4.000 484.520 796.000 485.160 ;
        RECT 4.000 483.120 795.600 484.520 ;
        RECT 4.000 481.800 796.000 483.120 ;
        RECT 4.000 480.400 795.600 481.800 ;
        RECT 4.000 479.760 796.000 480.400 ;
        RECT 4.000 478.360 795.600 479.760 ;
        RECT 4.000 477.720 796.000 478.360 ;
        RECT 4.400 477.040 796.000 477.720 ;
        RECT 4.400 476.320 795.600 477.040 ;
        RECT 4.000 475.640 795.600 476.320 ;
        RECT 4.000 474.320 796.000 475.640 ;
        RECT 4.000 472.920 795.600 474.320 ;
        RECT 4.000 472.280 796.000 472.920 ;
        RECT 4.000 470.880 795.600 472.280 ;
        RECT 4.000 469.560 796.000 470.880 ;
        RECT 4.000 468.880 795.600 469.560 ;
        RECT 4.400 468.160 795.600 468.880 ;
        RECT 4.400 467.520 796.000 468.160 ;
        RECT 4.400 467.480 795.600 467.520 ;
        RECT 4.000 466.120 795.600 467.480 ;
        RECT 4.000 464.800 796.000 466.120 ;
        RECT 4.000 463.400 795.600 464.800 ;
        RECT 4.000 462.760 796.000 463.400 ;
        RECT 4.000 461.360 795.600 462.760 ;
        RECT 4.000 460.040 796.000 461.360 ;
        RECT 4.400 458.640 795.600 460.040 ;
        RECT 4.000 458.000 796.000 458.640 ;
        RECT 4.000 456.600 795.600 458.000 ;
        RECT 4.000 455.280 796.000 456.600 ;
        RECT 4.000 453.880 795.600 455.280 ;
        RECT 4.000 452.560 796.000 453.880 ;
        RECT 4.000 451.200 795.600 452.560 ;
        RECT 4.400 451.160 795.600 451.200 ;
        RECT 4.400 450.520 796.000 451.160 ;
        RECT 4.400 449.800 795.600 450.520 ;
        RECT 4.000 449.120 795.600 449.800 ;
        RECT 4.000 447.800 796.000 449.120 ;
        RECT 4.000 446.400 795.600 447.800 ;
        RECT 4.000 445.760 796.000 446.400 ;
        RECT 4.000 444.360 795.600 445.760 ;
        RECT 4.000 443.040 796.000 444.360 ;
        RECT 4.000 442.360 795.600 443.040 ;
        RECT 4.400 441.640 795.600 442.360 ;
        RECT 4.400 441.000 796.000 441.640 ;
        RECT 4.400 440.960 795.600 441.000 ;
        RECT 4.000 439.600 795.600 440.960 ;
        RECT 4.000 438.280 796.000 439.600 ;
        RECT 4.000 436.880 795.600 438.280 ;
        RECT 4.000 436.240 796.000 436.880 ;
        RECT 4.000 434.840 795.600 436.240 ;
        RECT 4.000 433.520 796.000 434.840 ;
        RECT 4.400 432.120 795.600 433.520 ;
        RECT 4.000 431.480 796.000 432.120 ;
        RECT 4.000 430.080 795.600 431.480 ;
        RECT 4.000 428.760 796.000 430.080 ;
        RECT 4.000 427.360 795.600 428.760 ;
        RECT 4.000 426.040 796.000 427.360 ;
        RECT 4.000 424.640 795.600 426.040 ;
        RECT 4.000 424.000 796.000 424.640 ;
        RECT 4.400 422.600 795.600 424.000 ;
        RECT 4.000 421.280 796.000 422.600 ;
        RECT 4.000 419.880 795.600 421.280 ;
        RECT 4.000 419.240 796.000 419.880 ;
        RECT 4.000 417.840 795.600 419.240 ;
        RECT 4.000 416.520 796.000 417.840 ;
        RECT 4.000 415.160 795.600 416.520 ;
        RECT 4.400 415.120 795.600 415.160 ;
        RECT 4.400 414.480 796.000 415.120 ;
        RECT 4.400 413.760 795.600 414.480 ;
        RECT 4.000 413.080 795.600 413.760 ;
        RECT 4.000 411.760 796.000 413.080 ;
        RECT 4.000 410.360 795.600 411.760 ;
        RECT 4.000 409.720 796.000 410.360 ;
        RECT 4.000 408.320 795.600 409.720 ;
        RECT 4.000 407.000 796.000 408.320 ;
        RECT 4.000 406.320 795.600 407.000 ;
        RECT 4.400 405.600 795.600 406.320 ;
        RECT 4.400 404.920 796.000 405.600 ;
        RECT 4.000 404.280 796.000 404.920 ;
        RECT 4.000 402.880 795.600 404.280 ;
        RECT 4.000 402.240 796.000 402.880 ;
        RECT 4.000 400.840 795.600 402.240 ;
        RECT 4.000 399.520 796.000 400.840 ;
        RECT 4.000 398.120 795.600 399.520 ;
        RECT 4.000 397.480 796.000 398.120 ;
        RECT 4.400 396.080 795.600 397.480 ;
        RECT 4.000 394.760 796.000 396.080 ;
        RECT 4.000 393.360 795.600 394.760 ;
        RECT 4.000 392.720 796.000 393.360 ;
        RECT 4.000 391.320 795.600 392.720 ;
        RECT 4.000 390.000 796.000 391.320 ;
        RECT 4.000 388.640 795.600 390.000 ;
        RECT 4.400 388.600 795.600 388.640 ;
        RECT 4.400 387.960 796.000 388.600 ;
        RECT 4.400 387.240 795.600 387.960 ;
        RECT 4.000 386.560 795.600 387.240 ;
        RECT 4.000 385.240 796.000 386.560 ;
        RECT 4.000 383.840 795.600 385.240 ;
        RECT 4.000 383.200 796.000 383.840 ;
        RECT 4.000 381.800 795.600 383.200 ;
        RECT 4.000 380.480 796.000 381.800 ;
        RECT 4.000 379.800 795.600 380.480 ;
        RECT 4.400 379.080 795.600 379.800 ;
        RECT 4.400 378.400 796.000 379.080 ;
        RECT 4.000 377.760 796.000 378.400 ;
        RECT 4.000 376.360 795.600 377.760 ;
        RECT 4.000 375.720 796.000 376.360 ;
        RECT 4.000 374.320 795.600 375.720 ;
        RECT 4.000 373.000 796.000 374.320 ;
        RECT 4.000 371.600 795.600 373.000 ;
        RECT 4.000 370.960 796.000 371.600 ;
        RECT 4.400 369.560 795.600 370.960 ;
        RECT 4.000 368.240 796.000 369.560 ;
        RECT 4.000 366.840 795.600 368.240 ;
        RECT 4.000 366.200 796.000 366.840 ;
        RECT 4.000 364.800 795.600 366.200 ;
        RECT 4.000 363.480 796.000 364.800 ;
        RECT 4.000 362.120 795.600 363.480 ;
        RECT 4.400 362.080 795.600 362.120 ;
        RECT 4.400 361.440 796.000 362.080 ;
        RECT 4.400 360.720 795.600 361.440 ;
        RECT 4.000 360.040 795.600 360.720 ;
        RECT 4.000 358.720 796.000 360.040 ;
        RECT 4.000 357.320 795.600 358.720 ;
        RECT 4.000 356.000 796.000 357.320 ;
        RECT 4.000 354.600 795.600 356.000 ;
        RECT 4.000 353.960 796.000 354.600 ;
        RECT 4.000 352.600 795.600 353.960 ;
        RECT 4.400 352.560 795.600 352.600 ;
        RECT 4.400 351.240 796.000 352.560 ;
        RECT 4.400 351.200 795.600 351.240 ;
        RECT 4.000 349.840 795.600 351.200 ;
        RECT 4.000 349.200 796.000 349.840 ;
        RECT 4.000 347.800 795.600 349.200 ;
        RECT 4.000 346.480 796.000 347.800 ;
        RECT 4.000 345.080 795.600 346.480 ;
        RECT 4.000 344.440 796.000 345.080 ;
        RECT 4.000 343.760 795.600 344.440 ;
        RECT 4.400 343.040 795.600 343.760 ;
        RECT 4.400 342.360 796.000 343.040 ;
        RECT 4.000 341.720 796.000 342.360 ;
        RECT 4.000 340.320 795.600 341.720 ;
        RECT 4.000 339.680 796.000 340.320 ;
        RECT 4.000 338.280 795.600 339.680 ;
        RECT 4.000 336.960 796.000 338.280 ;
        RECT 4.000 335.560 795.600 336.960 ;
        RECT 4.000 334.920 796.000 335.560 ;
        RECT 4.400 333.520 795.600 334.920 ;
        RECT 4.000 332.200 796.000 333.520 ;
        RECT 4.000 330.800 795.600 332.200 ;
        RECT 4.000 329.480 796.000 330.800 ;
        RECT 4.000 328.080 795.600 329.480 ;
        RECT 4.000 327.440 796.000 328.080 ;
        RECT 4.000 326.080 795.600 327.440 ;
        RECT 4.400 326.040 795.600 326.080 ;
        RECT 4.400 324.720 796.000 326.040 ;
        RECT 4.400 324.680 795.600 324.720 ;
        RECT 4.000 323.320 795.600 324.680 ;
        RECT 4.000 322.680 796.000 323.320 ;
        RECT 4.000 321.280 795.600 322.680 ;
        RECT 4.000 319.960 796.000 321.280 ;
        RECT 4.000 318.560 795.600 319.960 ;
        RECT 4.000 317.920 796.000 318.560 ;
        RECT 4.000 317.240 795.600 317.920 ;
        RECT 4.400 316.520 795.600 317.240 ;
        RECT 4.400 315.840 796.000 316.520 ;
        RECT 4.000 315.200 796.000 315.840 ;
        RECT 4.000 313.800 795.600 315.200 ;
        RECT 4.000 313.160 796.000 313.800 ;
        RECT 4.000 311.760 795.600 313.160 ;
        RECT 4.000 310.440 796.000 311.760 ;
        RECT 4.000 309.040 795.600 310.440 ;
        RECT 4.000 308.400 796.000 309.040 ;
        RECT 4.400 307.720 796.000 308.400 ;
        RECT 4.400 307.000 795.600 307.720 ;
        RECT 4.000 306.320 795.600 307.000 ;
        RECT 4.000 305.680 796.000 306.320 ;
        RECT 4.000 304.280 795.600 305.680 ;
        RECT 4.000 302.960 796.000 304.280 ;
        RECT 4.000 301.560 795.600 302.960 ;
        RECT 4.000 300.920 796.000 301.560 ;
        RECT 4.000 299.560 795.600 300.920 ;
        RECT 4.400 299.520 795.600 299.560 ;
        RECT 4.400 298.200 796.000 299.520 ;
        RECT 4.400 298.160 795.600 298.200 ;
        RECT 4.000 296.800 795.600 298.160 ;
        RECT 4.000 296.160 796.000 296.800 ;
        RECT 4.000 294.760 795.600 296.160 ;
        RECT 4.000 293.440 796.000 294.760 ;
        RECT 4.000 292.040 795.600 293.440 ;
        RECT 4.000 291.400 796.000 292.040 ;
        RECT 4.000 290.720 795.600 291.400 ;
        RECT 4.400 290.000 795.600 290.720 ;
        RECT 4.400 289.320 796.000 290.000 ;
        RECT 4.000 288.680 796.000 289.320 ;
        RECT 4.000 287.280 795.600 288.680 ;
        RECT 4.000 285.960 796.000 287.280 ;
        RECT 4.000 284.560 795.600 285.960 ;
        RECT 4.000 283.920 796.000 284.560 ;
        RECT 4.000 282.520 795.600 283.920 ;
        RECT 4.000 281.200 796.000 282.520 ;
        RECT 4.400 279.800 795.600 281.200 ;
        RECT 4.000 279.160 796.000 279.800 ;
        RECT 4.000 277.760 795.600 279.160 ;
        RECT 4.000 276.440 796.000 277.760 ;
        RECT 4.000 275.040 795.600 276.440 ;
        RECT 4.000 274.400 796.000 275.040 ;
        RECT 4.000 273.000 795.600 274.400 ;
        RECT 4.000 272.360 796.000 273.000 ;
        RECT 4.400 271.680 796.000 272.360 ;
        RECT 4.400 270.960 795.600 271.680 ;
        RECT 4.000 270.280 795.600 270.960 ;
        RECT 4.000 269.640 796.000 270.280 ;
        RECT 4.000 268.240 795.600 269.640 ;
        RECT 4.000 266.920 796.000 268.240 ;
        RECT 4.000 265.520 795.600 266.920 ;
        RECT 4.000 264.880 796.000 265.520 ;
        RECT 4.000 263.520 795.600 264.880 ;
        RECT 4.400 263.480 795.600 263.520 ;
        RECT 4.400 262.160 796.000 263.480 ;
        RECT 4.400 262.120 795.600 262.160 ;
        RECT 4.000 260.760 795.600 262.120 ;
        RECT 4.000 259.440 796.000 260.760 ;
        RECT 4.000 258.040 795.600 259.440 ;
        RECT 4.000 257.400 796.000 258.040 ;
        RECT 4.000 256.000 795.600 257.400 ;
        RECT 4.000 254.680 796.000 256.000 ;
        RECT 4.400 253.280 795.600 254.680 ;
        RECT 4.000 252.640 796.000 253.280 ;
        RECT 4.000 251.240 795.600 252.640 ;
        RECT 4.000 249.920 796.000 251.240 ;
        RECT 4.000 248.520 795.600 249.920 ;
        RECT 4.000 247.880 796.000 248.520 ;
        RECT 4.000 246.480 795.600 247.880 ;
        RECT 4.000 245.840 796.000 246.480 ;
        RECT 4.400 245.160 796.000 245.840 ;
        RECT 4.400 244.440 795.600 245.160 ;
        RECT 4.000 243.760 795.600 244.440 ;
        RECT 4.000 243.120 796.000 243.760 ;
        RECT 4.000 241.720 795.600 243.120 ;
        RECT 4.000 240.400 796.000 241.720 ;
        RECT 4.000 239.000 795.600 240.400 ;
        RECT 4.000 237.680 796.000 239.000 ;
        RECT 4.000 237.000 795.600 237.680 ;
        RECT 4.400 236.280 795.600 237.000 ;
        RECT 4.400 235.640 796.000 236.280 ;
        RECT 4.400 235.600 795.600 235.640 ;
        RECT 4.000 234.240 795.600 235.600 ;
        RECT 4.000 232.920 796.000 234.240 ;
        RECT 4.000 231.520 795.600 232.920 ;
        RECT 4.000 230.880 796.000 231.520 ;
        RECT 4.000 229.480 795.600 230.880 ;
        RECT 4.000 228.160 796.000 229.480 ;
        RECT 4.400 226.760 795.600 228.160 ;
        RECT 4.000 226.120 796.000 226.760 ;
        RECT 4.000 224.720 795.600 226.120 ;
        RECT 4.000 223.400 796.000 224.720 ;
        RECT 4.000 222.000 795.600 223.400 ;
        RECT 4.000 221.360 796.000 222.000 ;
        RECT 4.000 219.960 795.600 221.360 ;
        RECT 4.000 219.320 796.000 219.960 ;
        RECT 4.400 218.640 796.000 219.320 ;
        RECT 4.400 217.920 795.600 218.640 ;
        RECT 4.000 217.240 795.600 217.920 ;
        RECT 4.000 216.600 796.000 217.240 ;
        RECT 4.000 215.200 795.600 216.600 ;
        RECT 4.000 213.880 796.000 215.200 ;
        RECT 4.000 212.480 795.600 213.880 ;
        RECT 4.000 211.160 796.000 212.480 ;
        RECT 4.000 209.800 795.600 211.160 ;
        RECT 4.400 209.760 795.600 209.800 ;
        RECT 4.400 209.120 796.000 209.760 ;
        RECT 4.400 208.400 795.600 209.120 ;
        RECT 4.000 207.720 795.600 208.400 ;
        RECT 4.000 206.400 796.000 207.720 ;
        RECT 4.000 205.000 795.600 206.400 ;
        RECT 4.000 204.360 796.000 205.000 ;
        RECT 4.000 202.960 795.600 204.360 ;
        RECT 4.000 201.640 796.000 202.960 ;
        RECT 4.000 200.960 795.600 201.640 ;
        RECT 4.400 200.240 795.600 200.960 ;
        RECT 4.400 199.600 796.000 200.240 ;
        RECT 4.400 199.560 795.600 199.600 ;
        RECT 4.000 198.200 795.600 199.560 ;
        RECT 4.000 196.880 796.000 198.200 ;
        RECT 4.000 195.480 795.600 196.880 ;
        RECT 4.000 194.840 796.000 195.480 ;
        RECT 4.000 193.440 795.600 194.840 ;
        RECT 4.000 192.120 796.000 193.440 ;
        RECT 4.400 190.720 795.600 192.120 ;
        RECT 4.000 189.400 796.000 190.720 ;
        RECT 4.000 188.000 795.600 189.400 ;
        RECT 4.000 187.360 796.000 188.000 ;
        RECT 4.000 185.960 795.600 187.360 ;
        RECT 4.000 184.640 796.000 185.960 ;
        RECT 4.000 183.280 795.600 184.640 ;
        RECT 4.400 183.240 795.600 183.280 ;
        RECT 4.400 182.600 796.000 183.240 ;
        RECT 4.400 181.880 795.600 182.600 ;
        RECT 4.000 181.200 795.600 181.880 ;
        RECT 4.000 179.880 796.000 181.200 ;
        RECT 4.000 178.480 795.600 179.880 ;
        RECT 4.000 177.840 796.000 178.480 ;
        RECT 4.000 176.440 795.600 177.840 ;
        RECT 4.000 175.120 796.000 176.440 ;
        RECT 4.000 174.440 795.600 175.120 ;
        RECT 4.400 173.720 795.600 174.440 ;
        RECT 4.400 173.080 796.000 173.720 ;
        RECT 4.400 173.040 795.600 173.080 ;
        RECT 4.000 171.680 795.600 173.040 ;
        RECT 4.000 170.360 796.000 171.680 ;
        RECT 4.000 168.960 795.600 170.360 ;
        RECT 4.000 168.320 796.000 168.960 ;
        RECT 4.000 166.920 795.600 168.320 ;
        RECT 4.000 165.600 796.000 166.920 ;
        RECT 4.400 164.200 795.600 165.600 ;
        RECT 4.000 162.880 796.000 164.200 ;
        RECT 4.000 161.480 795.600 162.880 ;
        RECT 4.000 160.840 796.000 161.480 ;
        RECT 4.000 159.440 795.600 160.840 ;
        RECT 4.000 158.120 796.000 159.440 ;
        RECT 4.000 156.760 795.600 158.120 ;
        RECT 4.400 156.720 795.600 156.760 ;
        RECT 4.400 156.080 796.000 156.720 ;
        RECT 4.400 155.360 795.600 156.080 ;
        RECT 4.000 154.680 795.600 155.360 ;
        RECT 4.000 153.360 796.000 154.680 ;
        RECT 4.000 151.960 795.600 153.360 ;
        RECT 4.000 151.320 796.000 151.960 ;
        RECT 4.000 149.920 795.600 151.320 ;
        RECT 4.000 148.600 796.000 149.920 ;
        RECT 4.000 147.920 795.600 148.600 ;
        RECT 4.400 147.200 795.600 147.920 ;
        RECT 4.400 146.560 796.000 147.200 ;
        RECT 4.400 146.520 795.600 146.560 ;
        RECT 4.000 145.160 795.600 146.520 ;
        RECT 4.000 143.840 796.000 145.160 ;
        RECT 4.000 142.440 795.600 143.840 ;
        RECT 4.000 141.120 796.000 142.440 ;
        RECT 4.000 139.720 795.600 141.120 ;
        RECT 4.000 139.080 796.000 139.720 ;
        RECT 4.000 138.400 795.600 139.080 ;
        RECT 4.400 137.680 795.600 138.400 ;
        RECT 4.400 137.000 796.000 137.680 ;
        RECT 4.000 136.360 796.000 137.000 ;
        RECT 4.000 134.960 795.600 136.360 ;
        RECT 4.000 134.320 796.000 134.960 ;
        RECT 4.000 132.920 795.600 134.320 ;
        RECT 4.000 131.600 796.000 132.920 ;
        RECT 4.000 130.200 795.600 131.600 ;
        RECT 4.000 129.560 796.000 130.200 ;
        RECT 4.400 128.160 795.600 129.560 ;
        RECT 4.000 126.840 796.000 128.160 ;
        RECT 4.000 125.440 795.600 126.840 ;
        RECT 4.000 124.800 796.000 125.440 ;
        RECT 4.000 123.400 795.600 124.800 ;
        RECT 4.000 122.080 796.000 123.400 ;
        RECT 4.000 120.720 795.600 122.080 ;
        RECT 4.400 120.680 795.600 120.720 ;
        RECT 4.400 119.360 796.000 120.680 ;
        RECT 4.400 119.320 795.600 119.360 ;
        RECT 4.000 117.960 795.600 119.320 ;
        RECT 4.000 117.320 796.000 117.960 ;
        RECT 4.000 115.920 795.600 117.320 ;
        RECT 4.000 114.600 796.000 115.920 ;
        RECT 4.000 113.200 795.600 114.600 ;
        RECT 4.000 112.560 796.000 113.200 ;
        RECT 4.000 111.880 795.600 112.560 ;
        RECT 4.400 111.160 795.600 111.880 ;
        RECT 4.400 110.480 796.000 111.160 ;
        RECT 4.000 109.840 796.000 110.480 ;
        RECT 4.000 108.440 795.600 109.840 ;
        RECT 4.000 107.800 796.000 108.440 ;
        RECT 4.000 106.400 795.600 107.800 ;
        RECT 4.000 105.080 796.000 106.400 ;
        RECT 4.000 103.680 795.600 105.080 ;
        RECT 4.000 103.040 796.000 103.680 ;
        RECT 4.400 101.640 795.600 103.040 ;
        RECT 4.000 100.320 796.000 101.640 ;
        RECT 4.000 98.920 795.600 100.320 ;
        RECT 4.000 98.280 796.000 98.920 ;
        RECT 4.000 96.880 795.600 98.280 ;
        RECT 4.000 95.560 796.000 96.880 ;
        RECT 4.000 94.200 795.600 95.560 ;
        RECT 4.400 94.160 795.600 94.200 ;
        RECT 4.400 92.840 796.000 94.160 ;
        RECT 4.400 92.800 795.600 92.840 ;
        RECT 4.000 91.440 795.600 92.800 ;
        RECT 4.000 90.800 796.000 91.440 ;
        RECT 4.000 89.400 795.600 90.800 ;
        RECT 4.000 88.080 796.000 89.400 ;
        RECT 4.000 86.680 795.600 88.080 ;
        RECT 4.000 86.040 796.000 86.680 ;
        RECT 4.000 85.360 795.600 86.040 ;
        RECT 4.400 84.640 795.600 85.360 ;
        RECT 4.400 83.960 796.000 84.640 ;
        RECT 4.000 83.320 796.000 83.960 ;
        RECT 4.000 81.920 795.600 83.320 ;
        RECT 4.000 81.280 796.000 81.920 ;
        RECT 4.000 79.880 795.600 81.280 ;
        RECT 4.000 78.560 796.000 79.880 ;
        RECT 4.000 77.160 795.600 78.560 ;
        RECT 4.000 76.520 796.000 77.160 ;
        RECT 4.400 75.120 795.600 76.520 ;
        RECT 4.000 73.800 796.000 75.120 ;
        RECT 4.000 72.400 795.600 73.800 ;
        RECT 4.000 71.080 796.000 72.400 ;
        RECT 4.000 69.680 795.600 71.080 ;
        RECT 4.000 69.040 796.000 69.680 ;
        RECT 4.000 67.640 795.600 69.040 ;
        RECT 4.000 67.000 796.000 67.640 ;
        RECT 4.400 66.320 796.000 67.000 ;
        RECT 4.400 65.600 795.600 66.320 ;
        RECT 4.000 64.920 795.600 65.600 ;
        RECT 4.000 64.280 796.000 64.920 ;
        RECT 4.000 62.880 795.600 64.280 ;
        RECT 4.000 61.560 796.000 62.880 ;
        RECT 4.000 60.160 795.600 61.560 ;
        RECT 4.000 59.520 796.000 60.160 ;
        RECT 4.000 58.160 795.600 59.520 ;
        RECT 4.400 58.120 795.600 58.160 ;
        RECT 4.400 56.800 796.000 58.120 ;
        RECT 4.400 56.760 795.600 56.800 ;
        RECT 4.000 55.400 795.600 56.760 ;
        RECT 4.000 54.760 796.000 55.400 ;
        RECT 4.000 53.360 795.600 54.760 ;
        RECT 4.000 52.040 796.000 53.360 ;
        RECT 4.000 50.640 795.600 52.040 ;
        RECT 4.000 50.000 796.000 50.640 ;
        RECT 4.000 49.320 795.600 50.000 ;
        RECT 4.400 48.600 795.600 49.320 ;
        RECT 4.400 47.920 796.000 48.600 ;
        RECT 4.000 47.280 796.000 47.920 ;
        RECT 4.000 45.880 795.600 47.280 ;
        RECT 4.000 44.560 796.000 45.880 ;
        RECT 4.000 43.160 795.600 44.560 ;
        RECT 4.000 42.520 796.000 43.160 ;
        RECT 4.000 41.120 795.600 42.520 ;
        RECT 4.000 40.480 796.000 41.120 ;
        RECT 4.400 39.800 796.000 40.480 ;
        RECT 4.400 39.080 795.600 39.800 ;
        RECT 4.000 38.400 795.600 39.080 ;
        RECT 4.000 37.760 796.000 38.400 ;
        RECT 4.000 36.360 795.600 37.760 ;
        RECT 4.000 35.040 796.000 36.360 ;
        RECT 4.000 33.640 795.600 35.040 ;
        RECT 4.000 33.000 796.000 33.640 ;
        RECT 4.000 31.640 795.600 33.000 ;
        RECT 4.400 31.600 795.600 31.640 ;
        RECT 4.400 30.280 796.000 31.600 ;
        RECT 4.400 30.240 795.600 30.280 ;
        RECT 4.000 28.880 795.600 30.240 ;
        RECT 4.000 28.240 796.000 28.880 ;
        RECT 4.000 26.840 795.600 28.240 ;
        RECT 4.000 25.520 796.000 26.840 ;
        RECT 4.000 24.120 795.600 25.520 ;
        RECT 4.000 22.800 796.000 24.120 ;
        RECT 4.400 21.400 795.600 22.800 ;
        RECT 4.000 20.760 796.000 21.400 ;
        RECT 4.000 19.360 795.600 20.760 ;
        RECT 4.000 18.040 796.000 19.360 ;
        RECT 4.000 16.640 795.600 18.040 ;
        RECT 4.000 16.000 796.000 16.640 ;
        RECT 4.000 14.600 795.600 16.000 ;
        RECT 4.000 13.960 796.000 14.600 ;
        RECT 4.400 13.280 796.000 13.960 ;
        RECT 4.400 12.560 795.600 13.280 ;
        RECT 4.000 11.880 795.600 12.560 ;
        RECT 4.000 11.240 796.000 11.880 ;
        RECT 4.000 9.840 795.600 11.240 ;
        RECT 4.000 8.520 796.000 9.840 ;
        RECT 4.000 7.120 795.600 8.520 ;
        RECT 4.000 6.480 796.000 7.120 ;
        RECT 4.000 5.120 795.600 6.480 ;
        RECT 4.400 5.080 795.600 5.120 ;
        RECT 4.400 3.760 796.000 5.080 ;
        RECT 4.400 3.720 795.600 3.760 ;
        RECT 4.000 2.360 795.600 3.720 ;
        RECT 4.000 1.720 796.000 2.360 ;
        RECT 4.000 0.320 795.600 1.720 ;
        RECT 4.000 0.180 796.000 0.320 ;
      LAYER met4 ;
        RECT 111.615 487.520 786.305 489.425 ;
        RECT 111.615 10.240 174.240 487.520 ;
        RECT 176.640 10.240 251.040 487.520 ;
        RECT 253.440 10.240 327.840 487.520 ;
        RECT 330.240 10.240 404.640 487.520 ;
        RECT 407.040 10.240 481.440 487.520 ;
        RECT 483.840 10.240 558.240 487.520 ;
        RECT 560.640 10.240 635.040 487.520 ;
        RECT 637.440 10.240 711.840 487.520 ;
        RECT 714.240 10.240 786.305 487.520 ;
        RECT 111.615 0.175 786.305 10.240 ;
  END
END ExperiarCore
END LIBRARY

