magic
tech sky130A
magscale 1 2
timestamp 1651490879
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 1300 38824 37584
<< obsm2 >>
rect 1398 167 38162 39817
<< metal3 >>
rect 0 39720 800 39840
rect 39200 39584 40000 39704
rect 0 39312 800 39432
rect 39200 39176 40000 39296
rect 0 38904 800 39024
rect 39200 38768 40000 38888
rect 0 38496 800 38616
rect 39200 38360 40000 38480
rect 0 38088 800 38208
rect 39200 37952 40000 38072
rect 0 37680 800 37800
rect 39200 37544 40000 37664
rect 0 37272 800 37392
rect 39200 37136 40000 37256
rect 0 36864 800 36984
rect 39200 36728 40000 36848
rect 0 36456 800 36576
rect 39200 36320 40000 36440
rect 0 36048 800 36168
rect 39200 35912 40000 36032
rect 0 35640 800 35760
rect 0 35232 800 35352
rect 39200 35368 40000 35488
rect 0 34824 800 34944
rect 39200 34960 40000 35080
rect 0 34416 800 34536
rect 39200 34552 40000 34672
rect 0 34008 800 34128
rect 39200 34144 40000 34264
rect 0 33600 800 33720
rect 39200 33736 40000 33856
rect 0 33192 800 33312
rect 39200 33328 40000 33448
rect 0 32784 800 32904
rect 39200 32920 40000 33040
rect 0 32376 800 32496
rect 39200 32512 40000 32632
rect 0 31968 800 32088
rect 39200 32104 40000 32224
rect 0 31560 800 31680
rect 39200 31696 40000 31816
rect 0 31152 800 31272
rect 39200 31288 40000 31408
rect 0 30744 800 30864
rect 39200 30744 40000 30864
rect 0 30336 800 30456
rect 39200 30336 40000 30456
rect 0 29928 800 30048
rect 39200 29928 40000 30048
rect 0 29520 800 29640
rect 39200 29520 40000 29640
rect 0 29112 800 29232
rect 39200 29112 40000 29232
rect 0 28704 800 28824
rect 39200 28704 40000 28824
rect 0 28296 800 28416
rect 39200 28296 40000 28416
rect 0 27888 800 28008
rect 39200 27888 40000 28008
rect 0 27480 800 27600
rect 39200 27480 40000 27600
rect 0 27072 800 27192
rect 39200 27072 40000 27192
rect 0 26800 800 26920
rect 0 26392 800 26512
rect 39200 26528 40000 26648
rect 0 25984 800 26104
rect 39200 26120 40000 26240
rect 0 25576 800 25696
rect 39200 25712 40000 25832
rect 0 25168 800 25288
rect 39200 25304 40000 25424
rect 0 24760 800 24880
rect 39200 24896 40000 25016
rect 0 24352 800 24472
rect 39200 24488 40000 24608
rect 0 23944 800 24064
rect 39200 24080 40000 24200
rect 0 23536 800 23656
rect 39200 23672 40000 23792
rect 0 23128 800 23248
rect 39200 23264 40000 23384
rect 0 22720 800 22840
rect 39200 22856 40000 22976
rect 0 22312 800 22432
rect 39200 22448 40000 22568
rect 0 21904 800 22024
rect 39200 21904 40000 22024
rect 0 21496 800 21616
rect 39200 21496 40000 21616
rect 0 21088 800 21208
rect 39200 21088 40000 21208
rect 0 20680 800 20800
rect 39200 20680 40000 20800
rect 0 20272 800 20392
rect 39200 20272 40000 20392
rect 0 19864 800 19984
rect 39200 19864 40000 19984
rect 0 19456 800 19576
rect 39200 19456 40000 19576
rect 0 19048 800 19168
rect 39200 19048 40000 19168
rect 0 18640 800 18760
rect 39200 18640 40000 18760
rect 0 18232 800 18352
rect 39200 18232 40000 18352
rect 0 17824 800 17944
rect 39200 17688 40000 17808
rect 0 17416 800 17536
rect 39200 17280 40000 17400
rect 0 17008 800 17128
rect 39200 16872 40000 16992
rect 0 16600 800 16720
rect 39200 16464 40000 16584
rect 0 16192 800 16312
rect 39200 16056 40000 16176
rect 0 15784 800 15904
rect 39200 15648 40000 15768
rect 0 15376 800 15496
rect 39200 15240 40000 15360
rect 0 14968 800 15088
rect 39200 14832 40000 14952
rect 0 14560 800 14680
rect 39200 14424 40000 14544
rect 0 14152 800 14272
rect 39200 14016 40000 14136
rect 0 13744 800 13864
rect 0 13472 800 13592
rect 39200 13608 40000 13728
rect 0 13064 800 13184
rect 39200 13064 40000 13184
rect 0 12656 800 12776
rect 39200 12656 40000 12776
rect 0 12248 800 12368
rect 39200 12248 40000 12368
rect 0 11840 800 11960
rect 39200 11840 40000 11960
rect 0 11432 800 11552
rect 39200 11432 40000 11552
rect 0 11024 800 11144
rect 39200 11024 40000 11144
rect 0 10616 800 10736
rect 39200 10616 40000 10736
rect 0 10208 800 10328
rect 39200 10208 40000 10328
rect 0 9800 800 9920
rect 39200 9800 40000 9920
rect 0 9392 800 9512
rect 39200 9392 40000 9512
rect 0 8984 800 9104
rect 39200 8848 40000 8968
rect 0 8576 800 8696
rect 39200 8440 40000 8560
rect 0 8168 800 8288
rect 39200 8032 40000 8152
rect 0 7760 800 7880
rect 39200 7624 40000 7744
rect 0 7352 800 7472
rect 39200 7216 40000 7336
rect 0 6944 800 7064
rect 39200 6808 40000 6928
rect 0 6536 800 6656
rect 39200 6400 40000 6520
rect 0 6128 800 6248
rect 39200 5992 40000 6112
rect 0 5720 800 5840
rect 39200 5584 40000 5704
rect 0 5312 800 5432
rect 39200 5176 40000 5296
rect 0 4904 800 5024
rect 39200 4768 40000 4888
rect 0 4496 800 4616
rect 0 4088 800 4208
rect 39200 4224 40000 4344
rect 0 3680 800 3800
rect 39200 3816 40000 3936
rect 0 3272 800 3392
rect 39200 3408 40000 3528
rect 0 2864 800 2984
rect 39200 3000 40000 3120
rect 0 2456 800 2576
rect 39200 2592 40000 2712
rect 0 2048 800 2168
rect 39200 2184 40000 2304
rect 0 1640 800 1760
rect 39200 1776 40000 1896
rect 0 1232 800 1352
rect 39200 1368 40000 1488
rect 0 824 800 944
rect 39200 960 40000 1080
rect 0 416 800 536
rect 39200 552 40000 672
rect 0 144 800 264
rect 39200 144 40000 264
<< obsm3 >>
rect 880 39784 39200 39813
rect 880 39640 39120 39784
rect 800 39512 39120 39640
rect 880 39504 39120 39512
rect 880 39376 39200 39504
rect 880 39232 39120 39376
rect 800 39104 39120 39232
rect 880 39096 39120 39104
rect 880 38968 39200 39096
rect 880 38824 39120 38968
rect 800 38696 39120 38824
rect 880 38688 39120 38696
rect 880 38560 39200 38688
rect 880 38416 39120 38560
rect 800 38288 39120 38416
rect 880 38280 39120 38288
rect 880 38152 39200 38280
rect 880 38008 39120 38152
rect 800 37880 39120 38008
rect 880 37872 39120 37880
rect 880 37744 39200 37872
rect 880 37600 39120 37744
rect 800 37472 39120 37600
rect 880 37464 39120 37472
rect 880 37336 39200 37464
rect 880 37192 39120 37336
rect 800 37064 39120 37192
rect 880 37056 39120 37064
rect 880 36928 39200 37056
rect 880 36784 39120 36928
rect 800 36656 39120 36784
rect 880 36648 39120 36656
rect 880 36520 39200 36648
rect 880 36376 39120 36520
rect 800 36248 39120 36376
rect 880 36240 39120 36248
rect 880 36112 39200 36240
rect 880 35968 39120 36112
rect 800 35840 39120 35968
rect 880 35832 39120 35840
rect 880 35568 39200 35832
rect 880 35560 39120 35568
rect 800 35432 39120 35560
rect 880 35288 39120 35432
rect 880 35160 39200 35288
rect 880 35152 39120 35160
rect 800 35024 39120 35152
rect 880 34880 39120 35024
rect 880 34752 39200 34880
rect 880 34744 39120 34752
rect 800 34616 39120 34744
rect 880 34472 39120 34616
rect 880 34344 39200 34472
rect 880 34336 39120 34344
rect 800 34208 39120 34336
rect 880 34064 39120 34208
rect 880 33936 39200 34064
rect 880 33928 39120 33936
rect 800 33800 39120 33928
rect 880 33656 39120 33800
rect 880 33528 39200 33656
rect 880 33520 39120 33528
rect 800 33392 39120 33520
rect 880 33248 39120 33392
rect 880 33120 39200 33248
rect 880 33112 39120 33120
rect 800 32984 39120 33112
rect 880 32840 39120 32984
rect 880 32712 39200 32840
rect 880 32704 39120 32712
rect 800 32576 39120 32704
rect 880 32432 39120 32576
rect 880 32304 39200 32432
rect 880 32296 39120 32304
rect 800 32168 39120 32296
rect 880 32024 39120 32168
rect 880 31896 39200 32024
rect 880 31888 39120 31896
rect 800 31760 39120 31888
rect 880 31616 39120 31760
rect 880 31488 39200 31616
rect 880 31480 39120 31488
rect 800 31352 39120 31480
rect 880 31208 39120 31352
rect 880 31072 39200 31208
rect 800 30944 39200 31072
rect 880 30664 39120 30944
rect 800 30536 39200 30664
rect 880 30256 39120 30536
rect 800 30128 39200 30256
rect 880 29848 39120 30128
rect 800 29720 39200 29848
rect 880 29440 39120 29720
rect 800 29312 39200 29440
rect 880 29032 39120 29312
rect 800 28904 39200 29032
rect 880 28624 39120 28904
rect 800 28496 39200 28624
rect 880 28216 39120 28496
rect 800 28088 39200 28216
rect 880 27808 39120 28088
rect 800 27680 39200 27808
rect 880 27400 39120 27680
rect 800 27272 39200 27400
rect 880 26992 39120 27272
rect 880 26728 39200 26992
rect 880 26720 39120 26728
rect 800 26592 39120 26720
rect 880 26448 39120 26592
rect 880 26320 39200 26448
rect 880 26312 39120 26320
rect 800 26184 39120 26312
rect 880 26040 39120 26184
rect 880 25912 39200 26040
rect 880 25904 39120 25912
rect 800 25776 39120 25904
rect 880 25632 39120 25776
rect 880 25504 39200 25632
rect 880 25496 39120 25504
rect 800 25368 39120 25496
rect 880 25224 39120 25368
rect 880 25096 39200 25224
rect 880 25088 39120 25096
rect 800 24960 39120 25088
rect 880 24816 39120 24960
rect 880 24688 39200 24816
rect 880 24680 39120 24688
rect 800 24552 39120 24680
rect 880 24408 39120 24552
rect 880 24280 39200 24408
rect 880 24272 39120 24280
rect 800 24144 39120 24272
rect 880 24000 39120 24144
rect 880 23872 39200 24000
rect 880 23864 39120 23872
rect 800 23736 39120 23864
rect 880 23592 39120 23736
rect 880 23464 39200 23592
rect 880 23456 39120 23464
rect 800 23328 39120 23456
rect 880 23184 39120 23328
rect 880 23056 39200 23184
rect 880 23048 39120 23056
rect 800 22920 39120 23048
rect 880 22776 39120 22920
rect 880 22648 39200 22776
rect 880 22640 39120 22648
rect 800 22512 39120 22640
rect 880 22368 39120 22512
rect 880 22232 39200 22368
rect 800 22104 39200 22232
rect 880 21824 39120 22104
rect 800 21696 39200 21824
rect 880 21416 39120 21696
rect 800 21288 39200 21416
rect 880 21008 39120 21288
rect 800 20880 39200 21008
rect 880 20600 39120 20880
rect 800 20472 39200 20600
rect 880 20192 39120 20472
rect 800 20064 39200 20192
rect 880 19784 39120 20064
rect 800 19656 39200 19784
rect 880 19376 39120 19656
rect 800 19248 39200 19376
rect 880 18968 39120 19248
rect 800 18840 39200 18968
rect 880 18560 39120 18840
rect 800 18432 39200 18560
rect 880 18152 39120 18432
rect 800 18024 39200 18152
rect 880 17888 39200 18024
rect 880 17744 39120 17888
rect 800 17616 39120 17744
rect 880 17608 39120 17616
rect 880 17480 39200 17608
rect 880 17336 39120 17480
rect 800 17208 39120 17336
rect 880 17200 39120 17208
rect 880 17072 39200 17200
rect 880 16928 39120 17072
rect 800 16800 39120 16928
rect 880 16792 39120 16800
rect 880 16664 39200 16792
rect 880 16520 39120 16664
rect 800 16392 39120 16520
rect 880 16384 39120 16392
rect 880 16256 39200 16384
rect 880 16112 39120 16256
rect 800 15984 39120 16112
rect 880 15976 39120 15984
rect 880 15848 39200 15976
rect 880 15704 39120 15848
rect 800 15576 39120 15704
rect 880 15568 39120 15576
rect 880 15440 39200 15568
rect 880 15296 39120 15440
rect 800 15168 39120 15296
rect 880 15160 39120 15168
rect 880 15032 39200 15160
rect 880 14888 39120 15032
rect 800 14760 39120 14888
rect 880 14752 39120 14760
rect 880 14624 39200 14752
rect 880 14480 39120 14624
rect 800 14352 39120 14480
rect 880 14344 39120 14352
rect 880 14216 39200 14344
rect 880 14072 39120 14216
rect 800 13944 39120 14072
rect 880 13936 39120 13944
rect 880 13808 39200 13936
rect 880 13528 39120 13808
rect 880 13392 39200 13528
rect 800 13264 39200 13392
rect 880 12984 39120 13264
rect 800 12856 39200 12984
rect 880 12576 39120 12856
rect 800 12448 39200 12576
rect 880 12168 39120 12448
rect 800 12040 39200 12168
rect 880 11760 39120 12040
rect 800 11632 39200 11760
rect 880 11352 39120 11632
rect 800 11224 39200 11352
rect 880 10944 39120 11224
rect 800 10816 39200 10944
rect 880 10536 39120 10816
rect 800 10408 39200 10536
rect 880 10128 39120 10408
rect 800 10000 39200 10128
rect 880 9720 39120 10000
rect 800 9592 39200 9720
rect 880 9312 39120 9592
rect 800 9184 39200 9312
rect 880 9048 39200 9184
rect 880 8904 39120 9048
rect 800 8776 39120 8904
rect 880 8768 39120 8776
rect 880 8640 39200 8768
rect 880 8496 39120 8640
rect 800 8368 39120 8496
rect 880 8360 39120 8368
rect 880 8232 39200 8360
rect 880 8088 39120 8232
rect 800 7960 39120 8088
rect 880 7952 39120 7960
rect 880 7824 39200 7952
rect 880 7680 39120 7824
rect 800 7552 39120 7680
rect 880 7544 39120 7552
rect 880 7416 39200 7544
rect 880 7272 39120 7416
rect 800 7144 39120 7272
rect 880 7136 39120 7144
rect 880 7008 39200 7136
rect 880 6864 39120 7008
rect 800 6736 39120 6864
rect 880 6728 39120 6736
rect 880 6600 39200 6728
rect 880 6456 39120 6600
rect 800 6328 39120 6456
rect 880 6320 39120 6328
rect 880 6192 39200 6320
rect 880 6048 39120 6192
rect 800 5920 39120 6048
rect 880 5912 39120 5920
rect 880 5784 39200 5912
rect 880 5640 39120 5784
rect 800 5512 39120 5640
rect 880 5504 39120 5512
rect 880 5376 39200 5504
rect 880 5232 39120 5376
rect 800 5104 39120 5232
rect 880 5096 39120 5104
rect 880 4968 39200 5096
rect 880 4824 39120 4968
rect 800 4696 39120 4824
rect 880 4688 39120 4696
rect 880 4424 39200 4688
rect 880 4416 39120 4424
rect 800 4288 39120 4416
rect 880 4144 39120 4288
rect 880 4016 39200 4144
rect 880 4008 39120 4016
rect 800 3880 39120 4008
rect 880 3736 39120 3880
rect 880 3608 39200 3736
rect 880 3600 39120 3608
rect 800 3472 39120 3600
rect 880 3328 39120 3472
rect 880 3200 39200 3328
rect 880 3192 39120 3200
rect 800 3064 39120 3192
rect 880 2920 39120 3064
rect 880 2792 39200 2920
rect 880 2784 39120 2792
rect 800 2656 39120 2784
rect 880 2512 39120 2656
rect 880 2384 39200 2512
rect 880 2376 39120 2384
rect 800 2248 39120 2376
rect 880 2104 39120 2248
rect 880 1976 39200 2104
rect 880 1968 39120 1976
rect 800 1840 39120 1968
rect 880 1696 39120 1840
rect 880 1568 39200 1696
rect 880 1560 39120 1568
rect 800 1432 39120 1560
rect 880 1288 39120 1432
rect 880 1160 39200 1288
rect 880 1152 39120 1160
rect 800 1024 39120 1152
rect 880 880 39120 1024
rect 880 752 39200 880
rect 880 744 39120 752
rect 800 616 39120 744
rect 880 472 39120 616
rect 880 344 39200 472
rect 880 171 39120 344
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 39200 1368 40000 1488 6 peripheralBus_address[0]
port 1 nsew signal output
rlabel metal3 s 39200 15648 40000 15768 6 peripheralBus_address[10]
port 2 nsew signal output
rlabel metal3 s 39200 16872 40000 16992 6 peripheralBus_address[11]
port 3 nsew signal output
rlabel metal3 s 39200 18232 40000 18352 6 peripheralBus_address[12]
port 4 nsew signal output
rlabel metal3 s 39200 19456 40000 19576 6 peripheralBus_address[13]
port 5 nsew signal output
rlabel metal3 s 39200 20680 40000 20800 6 peripheralBus_address[14]
port 6 nsew signal output
rlabel metal3 s 39200 21904 40000 22024 6 peripheralBus_address[15]
port 7 nsew signal output
rlabel metal3 s 39200 23264 40000 23384 6 peripheralBus_address[16]
port 8 nsew signal output
rlabel metal3 s 39200 24488 40000 24608 6 peripheralBus_address[17]
port 9 nsew signal output
rlabel metal3 s 39200 25712 40000 25832 6 peripheralBus_address[18]
port 10 nsew signal output
rlabel metal3 s 39200 27072 40000 27192 6 peripheralBus_address[19]
port 11 nsew signal output
rlabel metal3 s 39200 3000 40000 3120 6 peripheralBus_address[1]
port 12 nsew signal output
rlabel metal3 s 39200 28296 40000 28416 6 peripheralBus_address[20]
port 13 nsew signal output
rlabel metal3 s 39200 29520 40000 29640 6 peripheralBus_address[21]
port 14 nsew signal output
rlabel metal3 s 39200 30744 40000 30864 6 peripheralBus_address[22]
port 15 nsew signal output
rlabel metal3 s 39200 32104 40000 32224 6 peripheralBus_address[23]
port 16 nsew signal output
rlabel metal3 s 39200 4768 40000 4888 6 peripheralBus_address[2]
port 17 nsew signal output
rlabel metal3 s 39200 6400 40000 6520 6 peripheralBus_address[3]
port 18 nsew signal output
rlabel metal3 s 39200 8032 40000 8152 6 peripheralBus_address[4]
port 19 nsew signal output
rlabel metal3 s 39200 9392 40000 9512 6 peripheralBus_address[5]
port 20 nsew signal output
rlabel metal3 s 39200 10616 40000 10736 6 peripheralBus_address[6]
port 21 nsew signal output
rlabel metal3 s 39200 11840 40000 11960 6 peripheralBus_address[7]
port 22 nsew signal output
rlabel metal3 s 39200 13064 40000 13184 6 peripheralBus_address[8]
port 23 nsew signal output
rlabel metal3 s 39200 14424 40000 14544 6 peripheralBus_address[9]
port 24 nsew signal output
rlabel metal3 s 39200 144 40000 264 6 peripheralBus_busy
port 25 nsew signal input
rlabel metal3 s 39200 1776 40000 1896 6 peripheralBus_byteSelect[0]
port 26 nsew signal output
rlabel metal3 s 39200 3408 40000 3528 6 peripheralBus_byteSelect[1]
port 27 nsew signal output
rlabel metal3 s 39200 5176 40000 5296 6 peripheralBus_byteSelect[2]
port 28 nsew signal output
rlabel metal3 s 39200 6808 40000 6928 6 peripheralBus_byteSelect[3]
port 29 nsew signal output
rlabel metal3 s 39200 2184 40000 2304 6 peripheralBus_dataRead[0]
port 30 nsew signal input
rlabel metal3 s 39200 16056 40000 16176 6 peripheralBus_dataRead[10]
port 31 nsew signal input
rlabel metal3 s 39200 17280 40000 17400 6 peripheralBus_dataRead[11]
port 32 nsew signal input
rlabel metal3 s 39200 18640 40000 18760 6 peripheralBus_dataRead[12]
port 33 nsew signal input
rlabel metal3 s 39200 19864 40000 19984 6 peripheralBus_dataRead[13]
port 34 nsew signal input
rlabel metal3 s 39200 21088 40000 21208 6 peripheralBus_dataRead[14]
port 35 nsew signal input
rlabel metal3 s 39200 22448 40000 22568 6 peripheralBus_dataRead[15]
port 36 nsew signal input
rlabel metal3 s 39200 23672 40000 23792 6 peripheralBus_dataRead[16]
port 37 nsew signal input
rlabel metal3 s 39200 24896 40000 25016 6 peripheralBus_dataRead[17]
port 38 nsew signal input
rlabel metal3 s 39200 26120 40000 26240 6 peripheralBus_dataRead[18]
port 39 nsew signal input
rlabel metal3 s 39200 27480 40000 27600 6 peripheralBus_dataRead[19]
port 40 nsew signal input
rlabel metal3 s 39200 3816 40000 3936 6 peripheralBus_dataRead[1]
port 41 nsew signal input
rlabel metal3 s 39200 28704 40000 28824 6 peripheralBus_dataRead[20]
port 42 nsew signal input
rlabel metal3 s 39200 29928 40000 30048 6 peripheralBus_dataRead[21]
port 43 nsew signal input
rlabel metal3 s 39200 31288 40000 31408 6 peripheralBus_dataRead[22]
port 44 nsew signal input
rlabel metal3 s 39200 32512 40000 32632 6 peripheralBus_dataRead[23]
port 45 nsew signal input
rlabel metal3 s 39200 33328 40000 33448 6 peripheralBus_dataRead[24]
port 46 nsew signal input
rlabel metal3 s 39200 34144 40000 34264 6 peripheralBus_dataRead[25]
port 47 nsew signal input
rlabel metal3 s 39200 34960 40000 35080 6 peripheralBus_dataRead[26]
port 48 nsew signal input
rlabel metal3 s 39200 35912 40000 36032 6 peripheralBus_dataRead[27]
port 49 nsew signal input
rlabel metal3 s 39200 36728 40000 36848 6 peripheralBus_dataRead[28]
port 50 nsew signal input
rlabel metal3 s 39200 37544 40000 37664 6 peripheralBus_dataRead[29]
port 51 nsew signal input
rlabel metal3 s 39200 5584 40000 5704 6 peripheralBus_dataRead[2]
port 52 nsew signal input
rlabel metal3 s 39200 38360 40000 38480 6 peripheralBus_dataRead[30]
port 53 nsew signal input
rlabel metal3 s 39200 39176 40000 39296 6 peripheralBus_dataRead[31]
port 54 nsew signal input
rlabel metal3 s 39200 7216 40000 7336 6 peripheralBus_dataRead[3]
port 55 nsew signal input
rlabel metal3 s 39200 8440 40000 8560 6 peripheralBus_dataRead[4]
port 56 nsew signal input
rlabel metal3 s 39200 9800 40000 9920 6 peripheralBus_dataRead[5]
port 57 nsew signal input
rlabel metal3 s 39200 11024 40000 11144 6 peripheralBus_dataRead[6]
port 58 nsew signal input
rlabel metal3 s 39200 12248 40000 12368 6 peripheralBus_dataRead[7]
port 59 nsew signal input
rlabel metal3 s 39200 13608 40000 13728 6 peripheralBus_dataRead[8]
port 60 nsew signal input
rlabel metal3 s 39200 14832 40000 14952 6 peripheralBus_dataRead[9]
port 61 nsew signal input
rlabel metal3 s 39200 2592 40000 2712 6 peripheralBus_dataWrite[0]
port 62 nsew signal output
rlabel metal3 s 39200 16464 40000 16584 6 peripheralBus_dataWrite[10]
port 63 nsew signal output
rlabel metal3 s 39200 17688 40000 17808 6 peripheralBus_dataWrite[11]
port 64 nsew signal output
rlabel metal3 s 39200 19048 40000 19168 6 peripheralBus_dataWrite[12]
port 65 nsew signal output
rlabel metal3 s 39200 20272 40000 20392 6 peripheralBus_dataWrite[13]
port 66 nsew signal output
rlabel metal3 s 39200 21496 40000 21616 6 peripheralBus_dataWrite[14]
port 67 nsew signal output
rlabel metal3 s 39200 22856 40000 22976 6 peripheralBus_dataWrite[15]
port 68 nsew signal output
rlabel metal3 s 39200 24080 40000 24200 6 peripheralBus_dataWrite[16]
port 69 nsew signal output
rlabel metal3 s 39200 25304 40000 25424 6 peripheralBus_dataWrite[17]
port 70 nsew signal output
rlabel metal3 s 39200 26528 40000 26648 6 peripheralBus_dataWrite[18]
port 71 nsew signal output
rlabel metal3 s 39200 27888 40000 28008 6 peripheralBus_dataWrite[19]
port 72 nsew signal output
rlabel metal3 s 39200 4224 40000 4344 6 peripheralBus_dataWrite[1]
port 73 nsew signal output
rlabel metal3 s 39200 29112 40000 29232 6 peripheralBus_dataWrite[20]
port 74 nsew signal output
rlabel metal3 s 39200 30336 40000 30456 6 peripheralBus_dataWrite[21]
port 75 nsew signal output
rlabel metal3 s 39200 31696 40000 31816 6 peripheralBus_dataWrite[22]
port 76 nsew signal output
rlabel metal3 s 39200 32920 40000 33040 6 peripheralBus_dataWrite[23]
port 77 nsew signal output
rlabel metal3 s 39200 33736 40000 33856 6 peripheralBus_dataWrite[24]
port 78 nsew signal output
rlabel metal3 s 39200 34552 40000 34672 6 peripheralBus_dataWrite[25]
port 79 nsew signal output
rlabel metal3 s 39200 35368 40000 35488 6 peripheralBus_dataWrite[26]
port 80 nsew signal output
rlabel metal3 s 39200 36320 40000 36440 6 peripheralBus_dataWrite[27]
port 81 nsew signal output
rlabel metal3 s 39200 37136 40000 37256 6 peripheralBus_dataWrite[28]
port 82 nsew signal output
rlabel metal3 s 39200 37952 40000 38072 6 peripheralBus_dataWrite[29]
port 83 nsew signal output
rlabel metal3 s 39200 5992 40000 6112 6 peripheralBus_dataWrite[2]
port 84 nsew signal output
rlabel metal3 s 39200 38768 40000 38888 6 peripheralBus_dataWrite[30]
port 85 nsew signal output
rlabel metal3 s 39200 39584 40000 39704 6 peripheralBus_dataWrite[31]
port 86 nsew signal output
rlabel metal3 s 39200 7624 40000 7744 6 peripheralBus_dataWrite[3]
port 87 nsew signal output
rlabel metal3 s 39200 8848 40000 8968 6 peripheralBus_dataWrite[4]
port 88 nsew signal output
rlabel metal3 s 39200 10208 40000 10328 6 peripheralBus_dataWrite[5]
port 89 nsew signal output
rlabel metal3 s 39200 11432 40000 11552 6 peripheralBus_dataWrite[6]
port 90 nsew signal output
rlabel metal3 s 39200 12656 40000 12776 6 peripheralBus_dataWrite[7]
port 91 nsew signal output
rlabel metal3 s 39200 14016 40000 14136 6 peripheralBus_dataWrite[8]
port 92 nsew signal output
rlabel metal3 s 39200 15240 40000 15360 6 peripheralBus_dataWrite[9]
port 93 nsew signal output
rlabel metal3 s 39200 552 40000 672 6 peripheralBus_oe
port 94 nsew signal output
rlabel metal3 s 39200 960 40000 1080 6 peripheralBus_we
port 95 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 96 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 96 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 97 nsew ground input
rlabel metal3 s 0 144 800 264 6 wb_ack_o
port 98 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 wb_adr_i[0]
port 99 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 wb_adr_i[10]
port 100 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 wb_adr_i[11]
port 101 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_adr_i[12]
port 102 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wb_adr_i[13]
port 103 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 wb_adr_i[14]
port 104 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 wb_adr_i[15]
port 105 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 wb_adr_i[16]
port 106 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wb_adr_i[17]
port 107 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 wb_adr_i[18]
port 108 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 wb_adr_i[19]
port 109 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 wb_adr_i[1]
port 110 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 wb_adr_i[20]
port 111 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 wb_adr_i[21]
port 112 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 wb_adr_i[22]
port 113 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 wb_adr_i[23]
port 114 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wb_adr_i[2]
port 115 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 wb_adr_i[3]
port 116 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 wb_adr_i[4]
port 117 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 wb_adr_i[5]
port 118 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 wb_adr_i[6]
port 119 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 wb_adr_i[7]
port 120 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 wb_adr_i[8]
port 121 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 wb_adr_i[9]
port 122 nsew signal input
rlabel metal3 s 0 416 800 536 6 wb_clk_i
port 123 nsew signal input
rlabel metal3 s 0 824 800 944 6 wb_cyc_i
port 124 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 wb_data_i[0]
port 125 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wb_data_i[10]
port 126 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 wb_data_i[11]
port 127 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wb_data_i[12]
port 128 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wb_data_i[13]
port 129 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 wb_data_i[14]
port 130 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 wb_data_i[15]
port 131 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 wb_data_i[16]
port 132 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 wb_data_i[17]
port 133 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 wb_data_i[18]
port 134 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 wb_data_i[19]
port 135 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 wb_data_i[1]
port 136 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 wb_data_i[20]
port 137 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 wb_data_i[21]
port 138 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 wb_data_i[22]
port 139 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 wb_data_i[23]
port 140 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 wb_data_i[24]
port 141 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 wb_data_i[25]
port 142 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 wb_data_i[26]
port 143 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 wb_data_i[27]
port 144 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 wb_data_i[28]
port 145 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 wb_data_i[29]
port 146 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 wb_data_i[2]
port 147 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 wb_data_i[30]
port 148 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 wb_data_i[31]
port 149 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 wb_data_i[3]
port 150 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 wb_data_i[4]
port 151 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 wb_data_i[5]
port 152 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 wb_data_i[6]
port 153 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 wb_data_i[7]
port 154 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 wb_data_i[8]
port 155 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 wb_data_i[9]
port 156 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 wb_data_o[0]
port 157 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 wb_data_o[10]
port 158 nsew signal output
rlabel metal3 s 0 18640 800 18760 6 wb_data_o[11]
port 159 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 wb_data_o[12]
port 160 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 wb_data_o[13]
port 161 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 wb_data_o[14]
port 162 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 wb_data_o[15]
port 163 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 wb_data_o[16]
port 164 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 wb_data_o[17]
port 165 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 wb_data_o[18]
port 166 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 wb_data_o[19]
port 167 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 wb_data_o[1]
port 168 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 wb_data_o[20]
port 169 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 wb_data_o[21]
port 170 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 wb_data_o[22]
port 171 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 wb_data_o[23]
port 172 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 wb_data_o[24]
port 173 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 wb_data_o[25]
port 174 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 wb_data_o[26]
port 175 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 wb_data_o[27]
port 176 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 wb_data_o[28]
port 177 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 wb_data_o[29]
port 178 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 wb_data_o[2]
port 179 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 wb_data_o[30]
port 180 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 wb_data_o[31]
port 181 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 wb_data_o[3]
port 182 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 wb_data_o[4]
port 183 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 wb_data_o[5]
port 184 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 wb_data_o[6]
port 185 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 wb_data_o[7]
port 186 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 wb_data_o[8]
port 187 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 wb_data_o[9]
port 188 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 wb_rst_i
port 189 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 wb_sel_i[0]
port 190 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 wb_sel_i[1]
port 191 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 wb_sel_i[2]
port 192 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 wb_sel_i[3]
port 193 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 wb_stall_o
port 194 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 wb_stb_i
port 195 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 wb_we_i
port 196 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1506638
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripheral_WBPeripheralBusInterface/runs/Peripheral_WBPeripheralBusInterface/results/finishing/WBPeripheralBusInterface.magic.gds
string GDS_START 159730
<< end >>

