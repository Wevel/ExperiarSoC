magic
tech sky130A
magscale 1 2
timestamp 1654252964
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 14 1640 69630 67584
<< metal2 >>
rect 294 69200 350 70000
rect 938 69200 994 70000
rect 1582 69200 1638 70000
rect 2318 69200 2374 70000
rect 2962 69200 3018 70000
rect 3698 69200 3754 70000
rect 4342 69200 4398 70000
rect 5078 69200 5134 70000
rect 5722 69200 5778 70000
rect 6458 69200 6514 70000
rect 7102 69200 7158 70000
rect 7838 69200 7894 70000
rect 8482 69200 8538 70000
rect 9126 69200 9182 70000
rect 9862 69200 9918 70000
rect 10506 69200 10562 70000
rect 11242 69200 11298 70000
rect 11886 69200 11942 70000
rect 12622 69200 12678 70000
rect 13266 69200 13322 70000
rect 14002 69200 14058 70000
rect 14646 69200 14702 70000
rect 15382 69200 15438 70000
rect 16026 69200 16082 70000
rect 16762 69200 16818 70000
rect 17406 69200 17462 70000
rect 18050 69200 18106 70000
rect 18786 69200 18842 70000
rect 19430 69200 19486 70000
rect 20166 69200 20222 70000
rect 20810 69200 20866 70000
rect 21546 69200 21602 70000
rect 22190 69200 22246 70000
rect 22926 69200 22982 70000
rect 23570 69200 23626 70000
rect 24306 69200 24362 70000
rect 24950 69200 25006 70000
rect 25686 69200 25742 70000
rect 26330 69200 26386 70000
rect 26974 69200 27030 70000
rect 27710 69200 27766 70000
rect 28354 69200 28410 70000
rect 29090 69200 29146 70000
rect 29734 69200 29790 70000
rect 30470 69200 30526 70000
rect 31114 69200 31170 70000
rect 31850 69200 31906 70000
rect 32494 69200 32550 70000
rect 33230 69200 33286 70000
rect 33874 69200 33930 70000
rect 34610 69200 34666 70000
rect 35254 69200 35310 70000
rect 35898 69200 35954 70000
rect 36634 69200 36690 70000
rect 37278 69200 37334 70000
rect 38014 69200 38070 70000
rect 38658 69200 38714 70000
rect 39394 69200 39450 70000
rect 40038 69200 40094 70000
rect 40774 69200 40830 70000
rect 41418 69200 41474 70000
rect 42154 69200 42210 70000
rect 42798 69200 42854 70000
rect 43534 69200 43590 70000
rect 44178 69200 44234 70000
rect 44822 69200 44878 70000
rect 45558 69200 45614 70000
rect 46202 69200 46258 70000
rect 46938 69200 46994 70000
rect 47582 69200 47638 70000
rect 48318 69200 48374 70000
rect 48962 69200 49018 70000
rect 49698 69200 49754 70000
rect 50342 69200 50398 70000
rect 51078 69200 51134 70000
rect 51722 69200 51778 70000
rect 52458 69200 52514 70000
rect 53102 69200 53158 70000
rect 53746 69200 53802 70000
rect 54482 69200 54538 70000
rect 55126 69200 55182 70000
rect 55862 69200 55918 70000
rect 56506 69200 56562 70000
rect 57242 69200 57298 70000
rect 57886 69200 57942 70000
rect 58622 69200 58678 70000
rect 59266 69200 59322 70000
rect 60002 69200 60058 70000
rect 60646 69200 60702 70000
rect 61382 69200 61438 70000
rect 62026 69200 62082 70000
rect 62670 69200 62726 70000
rect 63406 69200 63462 70000
rect 64050 69200 64106 70000
rect 64786 69200 64842 70000
rect 65430 69200 65486 70000
rect 66166 69200 66222 70000
rect 66810 69200 66866 70000
rect 67546 69200 67602 70000
rect 68190 69200 68246 70000
rect 68926 69200 68982 70000
rect 69570 69200 69626 70000
rect 294 0 350 800
rect 938 0 994 800
rect 1582 0 1638 800
rect 2226 0 2282 800
rect 2870 0 2926 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 4894 0 4950 800
rect 5538 0 5594 800
rect 6182 0 6238 800
rect 6826 0 6882 800
rect 7470 0 7526 800
rect 8206 0 8262 800
rect 8850 0 8906 800
rect 9494 0 9550 800
rect 10138 0 10194 800
rect 10782 0 10838 800
rect 11518 0 11574 800
rect 12162 0 12218 800
rect 12806 0 12862 800
rect 13450 0 13506 800
rect 14094 0 14150 800
rect 14738 0 14794 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18786 0 18842 800
rect 19430 0 19486 800
rect 20074 0 20130 800
rect 20718 0 20774 800
rect 21362 0 21418 800
rect 22006 0 22062 800
rect 22742 0 22798 800
rect 23386 0 23442 800
rect 24030 0 24086 800
rect 24674 0 24730 800
rect 25318 0 25374 800
rect 25962 0 26018 800
rect 26698 0 26754 800
rect 27342 0 27398 800
rect 27986 0 28042 800
rect 28630 0 28686 800
rect 29274 0 29330 800
rect 30010 0 30066 800
rect 30654 0 30710 800
rect 31298 0 31354 800
rect 31942 0 31998 800
rect 32586 0 32642 800
rect 33230 0 33286 800
rect 33966 0 34022 800
rect 34610 0 34666 800
rect 35254 0 35310 800
rect 35898 0 35954 800
rect 36542 0 36598 800
rect 37278 0 37334 800
rect 37922 0 37978 800
rect 38566 0 38622 800
rect 39210 0 39266 800
rect 39854 0 39910 800
rect 40498 0 40554 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44546 0 44602 800
rect 45190 0 45246 800
rect 45834 0 45890 800
rect 46478 0 46534 800
rect 47122 0 47178 800
rect 47766 0 47822 800
rect 48502 0 48558 800
rect 49146 0 49202 800
rect 49790 0 49846 800
rect 50434 0 50490 800
rect 51078 0 51134 800
rect 51722 0 51778 800
rect 52458 0 52514 800
rect 53102 0 53158 800
rect 53746 0 53802 800
rect 54390 0 54446 800
rect 55034 0 55090 800
rect 55770 0 55826 800
rect 56414 0 56470 800
rect 57058 0 57114 800
rect 57702 0 57758 800
rect 58346 0 58402 800
rect 58990 0 59046 800
rect 59726 0 59782 800
rect 60370 0 60426 800
rect 61014 0 61070 800
rect 61658 0 61714 800
rect 62302 0 62358 800
rect 63038 0 63094 800
rect 63682 0 63738 800
rect 64326 0 64382 800
rect 64970 0 65026 800
rect 65614 0 65670 800
rect 66258 0 66314 800
rect 66994 0 67050 800
rect 67638 0 67694 800
rect 68282 0 68338 800
rect 68926 0 68982 800
rect 69570 0 69626 800
<< obsm2 >>
rect 20 69144 238 69306
rect 406 69144 882 69306
rect 1050 69144 1526 69306
rect 1694 69144 2262 69306
rect 2430 69144 2906 69306
rect 3074 69144 3642 69306
rect 3810 69144 4286 69306
rect 4454 69144 5022 69306
rect 5190 69144 5666 69306
rect 5834 69144 6402 69306
rect 6570 69144 7046 69306
rect 7214 69144 7782 69306
rect 7950 69144 8426 69306
rect 8594 69144 9070 69306
rect 9238 69144 9806 69306
rect 9974 69144 10450 69306
rect 10618 69144 11186 69306
rect 11354 69144 11830 69306
rect 11998 69144 12566 69306
rect 12734 69144 13210 69306
rect 13378 69144 13946 69306
rect 14114 69144 14590 69306
rect 14758 69144 15326 69306
rect 15494 69144 15970 69306
rect 16138 69144 16706 69306
rect 16874 69144 17350 69306
rect 17518 69144 17994 69306
rect 18162 69144 18730 69306
rect 18898 69144 19374 69306
rect 19542 69144 20110 69306
rect 20278 69144 20754 69306
rect 20922 69144 21490 69306
rect 21658 69144 22134 69306
rect 22302 69144 22870 69306
rect 23038 69144 23514 69306
rect 23682 69144 24250 69306
rect 24418 69144 24894 69306
rect 25062 69144 25630 69306
rect 25798 69144 26274 69306
rect 26442 69144 26918 69306
rect 27086 69144 27654 69306
rect 27822 69144 28298 69306
rect 28466 69144 29034 69306
rect 29202 69144 29678 69306
rect 29846 69144 30414 69306
rect 30582 69144 31058 69306
rect 31226 69144 31794 69306
rect 31962 69144 32438 69306
rect 32606 69144 33174 69306
rect 33342 69144 33818 69306
rect 33986 69144 34554 69306
rect 34722 69144 35198 69306
rect 35366 69144 35842 69306
rect 36010 69144 36578 69306
rect 36746 69144 37222 69306
rect 37390 69144 37958 69306
rect 38126 69144 38602 69306
rect 38770 69144 39338 69306
rect 39506 69144 39982 69306
rect 40150 69144 40718 69306
rect 40886 69144 41362 69306
rect 41530 69144 42098 69306
rect 42266 69144 42742 69306
rect 42910 69144 43478 69306
rect 43646 69144 44122 69306
rect 44290 69144 44766 69306
rect 44934 69144 45502 69306
rect 45670 69144 46146 69306
rect 46314 69144 46882 69306
rect 47050 69144 47526 69306
rect 47694 69144 48262 69306
rect 48430 69144 48906 69306
rect 49074 69144 49642 69306
rect 49810 69144 50286 69306
rect 50454 69144 51022 69306
rect 51190 69144 51666 69306
rect 51834 69144 52402 69306
rect 52570 69144 53046 69306
rect 53214 69144 53690 69306
rect 53858 69144 54426 69306
rect 54594 69144 55070 69306
rect 55238 69144 55806 69306
rect 55974 69144 56450 69306
rect 56618 69144 57186 69306
rect 57354 69144 57830 69306
rect 57998 69144 58566 69306
rect 58734 69144 59210 69306
rect 59378 69144 59946 69306
rect 60114 69144 60590 69306
rect 60758 69144 61326 69306
rect 61494 69144 61970 69306
rect 62138 69144 62614 69306
rect 62782 69144 63350 69306
rect 63518 69144 63994 69306
rect 64162 69144 64730 69306
rect 64898 69144 65374 69306
rect 65542 69144 66110 69306
rect 66278 69144 66754 69306
rect 66922 69144 67490 69306
rect 67658 69144 68134 69306
rect 68302 69144 68870 69306
rect 69038 69144 69514 69306
rect 20 856 69624 69144
rect 20 734 238 856
rect 406 734 882 856
rect 1050 734 1526 856
rect 1694 734 2170 856
rect 2338 734 2814 856
rect 2982 734 3458 856
rect 3626 734 4194 856
rect 4362 734 4838 856
rect 5006 734 5482 856
rect 5650 734 6126 856
rect 6294 734 6770 856
rect 6938 734 7414 856
rect 7582 734 8150 856
rect 8318 734 8794 856
rect 8962 734 9438 856
rect 9606 734 10082 856
rect 10250 734 10726 856
rect 10894 734 11462 856
rect 11630 734 12106 856
rect 12274 734 12750 856
rect 12918 734 13394 856
rect 13562 734 14038 856
rect 14206 734 14682 856
rect 14850 734 15418 856
rect 15586 734 16062 856
rect 16230 734 16706 856
rect 16874 734 17350 856
rect 17518 734 17994 856
rect 18162 734 18730 856
rect 18898 734 19374 856
rect 19542 734 20018 856
rect 20186 734 20662 856
rect 20830 734 21306 856
rect 21474 734 21950 856
rect 22118 734 22686 856
rect 22854 734 23330 856
rect 23498 734 23974 856
rect 24142 734 24618 856
rect 24786 734 25262 856
rect 25430 734 25906 856
rect 26074 734 26642 856
rect 26810 734 27286 856
rect 27454 734 27930 856
rect 28098 734 28574 856
rect 28742 734 29218 856
rect 29386 734 29954 856
rect 30122 734 30598 856
rect 30766 734 31242 856
rect 31410 734 31886 856
rect 32054 734 32530 856
rect 32698 734 33174 856
rect 33342 734 33910 856
rect 34078 734 34554 856
rect 34722 734 35198 856
rect 35366 734 35842 856
rect 36010 734 36486 856
rect 36654 734 37222 856
rect 37390 734 37866 856
rect 38034 734 38510 856
rect 38678 734 39154 856
rect 39322 734 39798 856
rect 39966 734 40442 856
rect 40610 734 41178 856
rect 41346 734 41822 856
rect 41990 734 42466 856
rect 42634 734 43110 856
rect 43278 734 43754 856
rect 43922 734 44490 856
rect 44658 734 45134 856
rect 45302 734 45778 856
rect 45946 734 46422 856
rect 46590 734 47066 856
rect 47234 734 47710 856
rect 47878 734 48446 856
rect 48614 734 49090 856
rect 49258 734 49734 856
rect 49902 734 50378 856
rect 50546 734 51022 856
rect 51190 734 51666 856
rect 51834 734 52402 856
rect 52570 734 53046 856
rect 53214 734 53690 856
rect 53858 734 54334 856
rect 54502 734 54978 856
rect 55146 734 55714 856
rect 55882 734 56358 856
rect 56526 734 57002 856
rect 57170 734 57646 856
rect 57814 734 58290 856
rect 58458 734 58934 856
rect 59102 734 59670 856
rect 59838 734 60314 856
rect 60482 734 60958 856
rect 61126 734 61602 856
rect 61770 734 62246 856
rect 62414 734 62982 856
rect 63150 734 63626 856
rect 63794 734 64270 856
rect 64438 734 64914 856
rect 65082 734 65558 856
rect 65726 734 66202 856
rect 66370 734 66938 856
rect 67106 734 67582 856
rect 67750 734 68226 856
rect 68394 734 68870 856
rect 69038 734 69514 856
<< metal3 >>
rect 0 69232 800 69352
rect 0 67736 800 67856
rect 0 66240 800 66360
rect 0 64880 800 65000
rect 0 63384 800 63504
rect 69200 62976 70000 63096
rect 0 61888 800 62008
rect 0 60392 800 60512
rect 0 59032 800 59152
rect 0 57536 800 57656
rect 0 56040 800 56160
rect 0 54544 800 54664
rect 0 53184 800 53304
rect 0 51688 800 51808
rect 0 50192 800 50312
rect 0 48832 800 48952
rect 69200 48968 70000 49088
rect 0 47336 800 47456
rect 0 45840 800 45960
rect 0 44344 800 44464
rect 0 42984 800 43104
rect 0 41488 800 41608
rect 0 39992 800 40112
rect 0 38496 800 38616
rect 0 37136 800 37256
rect 0 35640 800 35760
rect 69200 34960 70000 35080
rect 0 34144 800 34264
rect 0 32784 800 32904
rect 0 31288 800 31408
rect 0 29792 800 29912
rect 0 28296 800 28416
rect 0 26936 800 27056
rect 0 25440 800 25560
rect 0 23944 800 24064
rect 0 22448 800 22568
rect 0 21088 800 21208
rect 69200 20952 70000 21072
rect 0 19592 800 19712
rect 0 18096 800 18216
rect 0 16736 800 16856
rect 0 15240 800 15360
rect 0 13744 800 13864
rect 0 12248 800 12368
rect 0 10888 800 11008
rect 0 9392 800 9512
rect 0 7896 800 8016
rect 69200 6944 70000 7064
rect 0 6400 800 6520
rect 0 5040 800 5160
rect 0 3544 800 3664
rect 0 2048 800 2168
rect 0 688 800 808
<< obsm3 >>
rect 880 69152 69200 69322
rect 798 67936 69200 69152
rect 880 67656 69200 67936
rect 798 66440 69200 67656
rect 880 66160 69200 66440
rect 798 65080 69200 66160
rect 880 64800 69200 65080
rect 798 63584 69200 64800
rect 880 63304 69200 63584
rect 798 63176 69200 63304
rect 798 62896 69120 63176
rect 798 62088 69200 62896
rect 880 61808 69200 62088
rect 798 60592 69200 61808
rect 880 60312 69200 60592
rect 798 59232 69200 60312
rect 880 58952 69200 59232
rect 798 57736 69200 58952
rect 880 57456 69200 57736
rect 798 56240 69200 57456
rect 880 55960 69200 56240
rect 798 54744 69200 55960
rect 880 54464 69200 54744
rect 798 53384 69200 54464
rect 880 53104 69200 53384
rect 798 51888 69200 53104
rect 880 51608 69200 51888
rect 798 50392 69200 51608
rect 880 50112 69200 50392
rect 798 49168 69200 50112
rect 798 49032 69120 49168
rect 880 48888 69120 49032
rect 880 48752 69200 48888
rect 798 47536 69200 48752
rect 880 47256 69200 47536
rect 798 46040 69200 47256
rect 880 45760 69200 46040
rect 798 44544 69200 45760
rect 880 44264 69200 44544
rect 798 43184 69200 44264
rect 880 42904 69200 43184
rect 798 41688 69200 42904
rect 880 41408 69200 41688
rect 798 40192 69200 41408
rect 880 39912 69200 40192
rect 798 38696 69200 39912
rect 880 38416 69200 38696
rect 798 37336 69200 38416
rect 880 37056 69200 37336
rect 798 35840 69200 37056
rect 880 35560 69200 35840
rect 798 35160 69200 35560
rect 798 34880 69120 35160
rect 798 34344 69200 34880
rect 880 34064 69200 34344
rect 798 32984 69200 34064
rect 880 32704 69200 32984
rect 798 31488 69200 32704
rect 880 31208 69200 31488
rect 798 29992 69200 31208
rect 880 29712 69200 29992
rect 798 28496 69200 29712
rect 880 28216 69200 28496
rect 798 27136 69200 28216
rect 880 26856 69200 27136
rect 798 25640 69200 26856
rect 880 25360 69200 25640
rect 798 24144 69200 25360
rect 880 23864 69200 24144
rect 798 22648 69200 23864
rect 880 22368 69200 22648
rect 798 21288 69200 22368
rect 880 21152 69200 21288
rect 880 21008 69120 21152
rect 798 20872 69120 21008
rect 798 19792 69200 20872
rect 880 19512 69200 19792
rect 798 18296 69200 19512
rect 880 18016 69200 18296
rect 798 16936 69200 18016
rect 880 16656 69200 16936
rect 798 15440 69200 16656
rect 880 15160 69200 15440
rect 798 13944 69200 15160
rect 880 13664 69200 13944
rect 798 12448 69200 13664
rect 880 12168 69200 12448
rect 798 11088 69200 12168
rect 880 10808 69200 11088
rect 798 9592 69200 10808
rect 880 9312 69200 9592
rect 798 8096 69200 9312
rect 880 7816 69200 8096
rect 798 7144 69200 7816
rect 798 6864 69120 7144
rect 798 6600 69200 6864
rect 880 6320 69200 6600
rect 798 5240 69200 6320
rect 880 4960 69200 5240
rect 798 3744 69200 4960
rect 880 3464 69200 3744
rect 798 2248 69200 3464
rect 880 1968 69200 2248
rect 798 888 69200 1968
rect 880 718 69200 888
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 4659 2483 19488 66469
rect 19968 2483 34848 66469
rect 35328 2483 50208 66469
rect 50688 2483 65568 66469
rect 66048 2483 66181 66469
<< labels >>
rlabel metal3 s 69200 34960 70000 35080 6 caravel_irq[0]
port 1 nsew signal output
rlabel metal3 s 69200 48968 70000 49088 6 caravel_irq[1]
port 2 nsew signal output
rlabel metal3 s 69200 62976 70000 63096 6 caravel_irq[2]
port 3 nsew signal output
rlabel metal3 s 0 69232 800 69352 6 caravel_irq[3]
port 4 nsew signal output
rlabel metal3 s 69200 6944 70000 7064 6 caravel_uart_rx
port 5 nsew signal input
rlabel metal3 s 69200 20952 70000 21072 6 caravel_uart_tx
port 6 nsew signal output
rlabel metal2 s 294 69200 350 70000 6 caravel_wb_ack_i
port 7 nsew signal input
rlabel metal2 s 4342 69200 4398 70000 6 caravel_wb_adr_o[0]
port 8 nsew signal output
rlabel metal2 s 27710 69200 27766 70000 6 caravel_wb_adr_o[10]
port 9 nsew signal output
rlabel metal2 s 29734 69200 29790 70000 6 caravel_wb_adr_o[11]
port 10 nsew signal output
rlabel metal2 s 31850 69200 31906 70000 6 caravel_wb_adr_o[12]
port 11 nsew signal output
rlabel metal2 s 33874 69200 33930 70000 6 caravel_wb_adr_o[13]
port 12 nsew signal output
rlabel metal2 s 35898 69200 35954 70000 6 caravel_wb_adr_o[14]
port 13 nsew signal output
rlabel metal2 s 38014 69200 38070 70000 6 caravel_wb_adr_o[15]
port 14 nsew signal output
rlabel metal2 s 40038 69200 40094 70000 6 caravel_wb_adr_o[16]
port 15 nsew signal output
rlabel metal2 s 42154 69200 42210 70000 6 caravel_wb_adr_o[17]
port 16 nsew signal output
rlabel metal2 s 44178 69200 44234 70000 6 caravel_wb_adr_o[18]
port 17 nsew signal output
rlabel metal2 s 46202 69200 46258 70000 6 caravel_wb_adr_o[19]
port 18 nsew signal output
rlabel metal2 s 7102 69200 7158 70000 6 caravel_wb_adr_o[1]
port 19 nsew signal output
rlabel metal2 s 48318 69200 48374 70000 6 caravel_wb_adr_o[20]
port 20 nsew signal output
rlabel metal2 s 50342 69200 50398 70000 6 caravel_wb_adr_o[21]
port 21 nsew signal output
rlabel metal2 s 52458 69200 52514 70000 6 caravel_wb_adr_o[22]
port 22 nsew signal output
rlabel metal2 s 54482 69200 54538 70000 6 caravel_wb_adr_o[23]
port 23 nsew signal output
rlabel metal2 s 56506 69200 56562 70000 6 caravel_wb_adr_o[24]
port 24 nsew signal output
rlabel metal2 s 58622 69200 58678 70000 6 caravel_wb_adr_o[25]
port 25 nsew signal output
rlabel metal2 s 60646 69200 60702 70000 6 caravel_wb_adr_o[26]
port 26 nsew signal output
rlabel metal2 s 62670 69200 62726 70000 6 caravel_wb_adr_o[27]
port 27 nsew signal output
rlabel metal2 s 9862 69200 9918 70000 6 caravel_wb_adr_o[2]
port 28 nsew signal output
rlabel metal2 s 12622 69200 12678 70000 6 caravel_wb_adr_o[3]
port 29 nsew signal output
rlabel metal2 s 15382 69200 15438 70000 6 caravel_wb_adr_o[4]
port 30 nsew signal output
rlabel metal2 s 17406 69200 17462 70000 6 caravel_wb_adr_o[5]
port 31 nsew signal output
rlabel metal2 s 19430 69200 19486 70000 6 caravel_wb_adr_o[6]
port 32 nsew signal output
rlabel metal2 s 21546 69200 21602 70000 6 caravel_wb_adr_o[7]
port 33 nsew signal output
rlabel metal2 s 23570 69200 23626 70000 6 caravel_wb_adr_o[8]
port 34 nsew signal output
rlabel metal2 s 25686 69200 25742 70000 6 caravel_wb_adr_o[9]
port 35 nsew signal output
rlabel metal2 s 938 69200 994 70000 6 caravel_wb_cyc_o
port 36 nsew signal output
rlabel metal2 s 5078 69200 5134 70000 6 caravel_wb_data_i[0]
port 37 nsew signal input
rlabel metal2 s 28354 69200 28410 70000 6 caravel_wb_data_i[10]
port 38 nsew signal input
rlabel metal2 s 30470 69200 30526 70000 6 caravel_wb_data_i[11]
port 39 nsew signal input
rlabel metal2 s 32494 69200 32550 70000 6 caravel_wb_data_i[12]
port 40 nsew signal input
rlabel metal2 s 34610 69200 34666 70000 6 caravel_wb_data_i[13]
port 41 nsew signal input
rlabel metal2 s 36634 69200 36690 70000 6 caravel_wb_data_i[14]
port 42 nsew signal input
rlabel metal2 s 38658 69200 38714 70000 6 caravel_wb_data_i[15]
port 43 nsew signal input
rlabel metal2 s 40774 69200 40830 70000 6 caravel_wb_data_i[16]
port 44 nsew signal input
rlabel metal2 s 42798 69200 42854 70000 6 caravel_wb_data_i[17]
port 45 nsew signal input
rlabel metal2 s 44822 69200 44878 70000 6 caravel_wb_data_i[18]
port 46 nsew signal input
rlabel metal2 s 46938 69200 46994 70000 6 caravel_wb_data_i[19]
port 47 nsew signal input
rlabel metal2 s 7838 69200 7894 70000 6 caravel_wb_data_i[1]
port 48 nsew signal input
rlabel metal2 s 48962 69200 49018 70000 6 caravel_wb_data_i[20]
port 49 nsew signal input
rlabel metal2 s 51078 69200 51134 70000 6 caravel_wb_data_i[21]
port 50 nsew signal input
rlabel metal2 s 53102 69200 53158 70000 6 caravel_wb_data_i[22]
port 51 nsew signal input
rlabel metal2 s 55126 69200 55182 70000 6 caravel_wb_data_i[23]
port 52 nsew signal input
rlabel metal2 s 57242 69200 57298 70000 6 caravel_wb_data_i[24]
port 53 nsew signal input
rlabel metal2 s 59266 69200 59322 70000 6 caravel_wb_data_i[25]
port 54 nsew signal input
rlabel metal2 s 61382 69200 61438 70000 6 caravel_wb_data_i[26]
port 55 nsew signal input
rlabel metal2 s 63406 69200 63462 70000 6 caravel_wb_data_i[27]
port 56 nsew signal input
rlabel metal2 s 64786 69200 64842 70000 6 caravel_wb_data_i[28]
port 57 nsew signal input
rlabel metal2 s 66166 69200 66222 70000 6 caravel_wb_data_i[29]
port 58 nsew signal input
rlabel metal2 s 10506 69200 10562 70000 6 caravel_wb_data_i[2]
port 59 nsew signal input
rlabel metal2 s 67546 69200 67602 70000 6 caravel_wb_data_i[30]
port 60 nsew signal input
rlabel metal2 s 68926 69200 68982 70000 6 caravel_wb_data_i[31]
port 61 nsew signal input
rlabel metal2 s 13266 69200 13322 70000 6 caravel_wb_data_i[3]
port 62 nsew signal input
rlabel metal2 s 16026 69200 16082 70000 6 caravel_wb_data_i[4]
port 63 nsew signal input
rlabel metal2 s 18050 69200 18106 70000 6 caravel_wb_data_i[5]
port 64 nsew signal input
rlabel metal2 s 20166 69200 20222 70000 6 caravel_wb_data_i[6]
port 65 nsew signal input
rlabel metal2 s 22190 69200 22246 70000 6 caravel_wb_data_i[7]
port 66 nsew signal input
rlabel metal2 s 24306 69200 24362 70000 6 caravel_wb_data_i[8]
port 67 nsew signal input
rlabel metal2 s 26330 69200 26386 70000 6 caravel_wb_data_i[9]
port 68 nsew signal input
rlabel metal2 s 5722 69200 5778 70000 6 caravel_wb_data_o[0]
port 69 nsew signal output
rlabel metal2 s 29090 69200 29146 70000 6 caravel_wb_data_o[10]
port 70 nsew signal output
rlabel metal2 s 31114 69200 31170 70000 6 caravel_wb_data_o[11]
port 71 nsew signal output
rlabel metal2 s 33230 69200 33286 70000 6 caravel_wb_data_o[12]
port 72 nsew signal output
rlabel metal2 s 35254 69200 35310 70000 6 caravel_wb_data_o[13]
port 73 nsew signal output
rlabel metal2 s 37278 69200 37334 70000 6 caravel_wb_data_o[14]
port 74 nsew signal output
rlabel metal2 s 39394 69200 39450 70000 6 caravel_wb_data_o[15]
port 75 nsew signal output
rlabel metal2 s 41418 69200 41474 70000 6 caravel_wb_data_o[16]
port 76 nsew signal output
rlabel metal2 s 43534 69200 43590 70000 6 caravel_wb_data_o[17]
port 77 nsew signal output
rlabel metal2 s 45558 69200 45614 70000 6 caravel_wb_data_o[18]
port 78 nsew signal output
rlabel metal2 s 47582 69200 47638 70000 6 caravel_wb_data_o[19]
port 79 nsew signal output
rlabel metal2 s 8482 69200 8538 70000 6 caravel_wb_data_o[1]
port 80 nsew signal output
rlabel metal2 s 49698 69200 49754 70000 6 caravel_wb_data_o[20]
port 81 nsew signal output
rlabel metal2 s 51722 69200 51778 70000 6 caravel_wb_data_o[21]
port 82 nsew signal output
rlabel metal2 s 53746 69200 53802 70000 6 caravel_wb_data_o[22]
port 83 nsew signal output
rlabel metal2 s 55862 69200 55918 70000 6 caravel_wb_data_o[23]
port 84 nsew signal output
rlabel metal2 s 57886 69200 57942 70000 6 caravel_wb_data_o[24]
port 85 nsew signal output
rlabel metal2 s 60002 69200 60058 70000 6 caravel_wb_data_o[25]
port 86 nsew signal output
rlabel metal2 s 62026 69200 62082 70000 6 caravel_wb_data_o[26]
port 87 nsew signal output
rlabel metal2 s 64050 69200 64106 70000 6 caravel_wb_data_o[27]
port 88 nsew signal output
rlabel metal2 s 65430 69200 65486 70000 6 caravel_wb_data_o[28]
port 89 nsew signal output
rlabel metal2 s 66810 69200 66866 70000 6 caravel_wb_data_o[29]
port 90 nsew signal output
rlabel metal2 s 11242 69200 11298 70000 6 caravel_wb_data_o[2]
port 91 nsew signal output
rlabel metal2 s 68190 69200 68246 70000 6 caravel_wb_data_o[30]
port 92 nsew signal output
rlabel metal2 s 69570 69200 69626 70000 6 caravel_wb_data_o[31]
port 93 nsew signal output
rlabel metal2 s 14002 69200 14058 70000 6 caravel_wb_data_o[3]
port 94 nsew signal output
rlabel metal2 s 16762 69200 16818 70000 6 caravel_wb_data_o[4]
port 95 nsew signal output
rlabel metal2 s 18786 69200 18842 70000 6 caravel_wb_data_o[5]
port 96 nsew signal output
rlabel metal2 s 20810 69200 20866 70000 6 caravel_wb_data_o[6]
port 97 nsew signal output
rlabel metal2 s 22926 69200 22982 70000 6 caravel_wb_data_o[7]
port 98 nsew signal output
rlabel metal2 s 24950 69200 25006 70000 6 caravel_wb_data_o[8]
port 99 nsew signal output
rlabel metal2 s 26974 69200 27030 70000 6 caravel_wb_data_o[9]
port 100 nsew signal output
rlabel metal2 s 1582 69200 1638 70000 6 caravel_wb_error_i
port 101 nsew signal input
rlabel metal2 s 6458 69200 6514 70000 6 caravel_wb_sel_o[0]
port 102 nsew signal output
rlabel metal2 s 9126 69200 9182 70000 6 caravel_wb_sel_o[1]
port 103 nsew signal output
rlabel metal2 s 11886 69200 11942 70000 6 caravel_wb_sel_o[2]
port 104 nsew signal output
rlabel metal2 s 14646 69200 14702 70000 6 caravel_wb_sel_o[3]
port 105 nsew signal output
rlabel metal2 s 2318 69200 2374 70000 6 caravel_wb_stall_i
port 106 nsew signal input
rlabel metal2 s 2962 69200 3018 70000 6 caravel_wb_stb_o
port 107 nsew signal output
rlabel metal2 s 3698 69200 3754 70000 6 caravel_wb_we_o
port 108 nsew signal output
rlabel metal3 s 0 688 800 808 6 core0Index[0]
port 109 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 core0Index[1]
port 110 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 core0Index[2]
port 111 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 core0Index[3]
port 112 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 core0Index[4]
port 113 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 core0Index[5]
port 114 nsew signal output
rlabel metal3 s 0 9392 800 9512 6 core0Index[6]
port 115 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 core0Index[7]
port 116 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 core1Index[0]
port 117 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 core1Index[1]
port 118 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 core1Index[2]
port 119 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 core1Index[3]
port 120 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 core1Index[4]
port 121 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 core1Index[5]
port 122 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 core1Index[6]
port 123 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 core1Index[7]
port 124 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 manufacturerID[0]
port 125 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 manufacturerID[10]
port 126 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 manufacturerID[1]
port 127 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 manufacturerID[2]
port 128 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 manufacturerID[3]
port 129 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 manufacturerID[4]
port 130 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 manufacturerID[5]
port 131 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 manufacturerID[6]
port 132 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 manufacturerID[7]
port 133 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 manufacturerID[8]
port 134 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 manufacturerID[9]
port 135 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 partID[0]
port 136 nsew signal output
rlabel metal3 s 0 54544 800 54664 6 partID[10]
port 137 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 partID[11]
port 138 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 partID[12]
port 139 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 partID[13]
port 140 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 partID[14]
port 141 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 partID[15]
port 142 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 partID[1]
port 143 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 partID[2]
port 144 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 partID[3]
port 145 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 partID[4]
port 146 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 partID[5]
port 147 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 partID[6]
port 148 nsew signal output
rlabel metal3 s 0 50192 800 50312 6 partID[7]
port 149 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 partID[8]
port 150 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 partID[9]
port 151 nsew signal output
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 152 nsew power input
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 152 nsew power input
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 152 nsew power input
rlabel metal3 s 0 63384 800 63504 6 versionID[0]
port 153 nsew signal output
rlabel metal3 s 0 64880 800 65000 6 versionID[1]
port 154 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 versionID[2]
port 155 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 versionID[3]
port 156 nsew signal output
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 157 nsew ground input
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 157 nsew ground input
rlabel metal2 s 294 0 350 800 6 wb_clk_i
port 158 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_rst_i
port 159 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_ack_o
port 160 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[0]
port 161 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[10]
port 162 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[11]
port 163 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[12]
port 164 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_adr_i[13]
port 165 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_adr_i[14]
port 166 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_adr_i[15]
port 167 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_adr_i[16]
port 168 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[17]
port 169 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[18]
port 170 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_adr_i[19]
port 171 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[1]
port 172 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[20]
port 173 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 wbs_adr_i[21]
port 174 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[22]
port 175 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_adr_i[23]
port 176 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_adr_i[24]
port 177 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 wbs_adr_i[25]
port 178 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 wbs_adr_i[26]
port 179 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 wbs_adr_i[27]
port 180 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 wbs_adr_i[28]
port 181 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 wbs_adr_i[29]
port 182 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_adr_i[2]
port 183 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wbs_adr_i[30]
port 184 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 wbs_adr_i[31]
port 185 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[3]
port 186 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[4]
port 187 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[5]
port 188 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[6]
port 189 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wbs_adr_i[7]
port 190 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[8]
port 191 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[9]
port 192 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_cyc_i
port 193 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 wbs_data_i[0]
port 194 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_data_i[10]
port 195 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_data_i[11]
port 196 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_data_i[12]
port 197 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_data_i[13]
port 198 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_data_i[14]
port 199 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_data_i[15]
port 200 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_data_i[16]
port 201 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 wbs_data_i[17]
port 202 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_data_i[18]
port 203 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 wbs_data_i[19]
port 204 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_data_i[1]
port 205 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_data_i[20]
port 206 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_data_i[21]
port 207 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_data_i[22]
port 208 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_data_i[23]
port 209 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_data_i[24]
port 210 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 wbs_data_i[25]
port 211 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wbs_data_i[26]
port 212 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 wbs_data_i[27]
port 213 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_data_i[28]
port 214 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 wbs_data_i[29]
port 215 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_data_i[2]
port 216 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 wbs_data_i[30]
port 217 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 wbs_data_i[31]
port 218 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_data_i[3]
port 219 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 wbs_data_i[4]
port 220 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_data_i[5]
port 221 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_data_i[6]
port 222 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_data_i[7]
port 223 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_data_i[8]
port 224 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_data_i[9]
port 225 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_data_o[0]
port 226 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_data_o[10]
port 227 nsew signal output
rlabel metal2 s 30010 0 30066 800 6 wbs_data_o[11]
port 228 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_data_o[12]
port 229 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 wbs_data_o[13]
port 230 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 wbs_data_o[14]
port 231 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_data_o[15]
port 232 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 wbs_data_o[16]
port 233 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 wbs_data_o[17]
port 234 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 wbs_data_o[18]
port 235 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 wbs_data_o[19]
port 236 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 wbs_data_o[1]
port 237 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 wbs_data_o[20]
port 238 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 wbs_data_o[21]
port 239 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_data_o[22]
port 240 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 wbs_data_o[23]
port 241 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 wbs_data_o[24]
port 242 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 wbs_data_o[25]
port 243 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 wbs_data_o[26]
port 244 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 wbs_data_o[27]
port 245 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 wbs_data_o[28]
port 246 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 wbs_data_o[29]
port 247 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_data_o[2]
port 248 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 wbs_data_o[30]
port 249 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 wbs_data_o[31]
port 250 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_data_o[3]
port 251 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_data_o[4]
port 252 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_data_o[5]
port 253 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_data_o[6]
port 254 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 wbs_data_o[7]
port 255 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_data_o[8]
port 256 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 wbs_data_o[9]
port 257 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[0]
port 258 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_sel_i[1]
port 259 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_sel_i[2]
port 260 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_sel_i[3]
port 261 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_stb_i
port 262 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_we_i
port 263 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13321600
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/CaravelHost/runs/CaravelHost/results/finishing/CaravelHost.magic.gds
string GDS_START 852336
<< end >>

