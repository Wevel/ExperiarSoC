magic
tech sky130A
magscale 1 2
timestamp 1652991016
<< obsli1 >>
rect 1104 2159 98808 137649
<< obsm1 >>
rect 1104 2128 99530 137896
<< metal2 >>
rect 386 139200 442 140000
rect 1214 139200 1270 140000
rect 2134 139200 2190 140000
rect 2962 139200 3018 140000
rect 3882 139200 3938 140000
rect 4710 139200 4766 140000
rect 5630 139200 5686 140000
rect 6458 139200 6514 140000
rect 7378 139200 7434 140000
rect 8206 139200 8262 140000
rect 9126 139200 9182 140000
rect 9954 139200 10010 140000
rect 10874 139200 10930 140000
rect 11702 139200 11758 140000
rect 12622 139200 12678 140000
rect 13542 139200 13598 140000
rect 14370 139200 14426 140000
rect 15290 139200 15346 140000
rect 16118 139200 16174 140000
rect 17038 139200 17094 140000
rect 17866 139200 17922 140000
rect 18786 139200 18842 140000
rect 19614 139200 19670 140000
rect 20534 139200 20590 140000
rect 21362 139200 21418 140000
rect 22282 139200 22338 140000
rect 23110 139200 23166 140000
rect 24030 139200 24086 140000
rect 24858 139200 24914 140000
rect 25778 139200 25834 140000
rect 26698 139200 26754 140000
rect 27526 139200 27582 140000
rect 28446 139200 28502 140000
rect 29274 139200 29330 140000
rect 30194 139200 30250 140000
rect 31022 139200 31078 140000
rect 31942 139200 31998 140000
rect 32770 139200 32826 140000
rect 33690 139200 33746 140000
rect 34518 139200 34574 140000
rect 35438 139200 35494 140000
rect 36266 139200 36322 140000
rect 37186 139200 37242 140000
rect 38106 139200 38162 140000
rect 38934 139200 38990 140000
rect 39854 139200 39910 140000
rect 40682 139200 40738 140000
rect 41602 139200 41658 140000
rect 42430 139200 42486 140000
rect 43350 139200 43406 140000
rect 44178 139200 44234 140000
rect 45098 139200 45154 140000
rect 45926 139200 45982 140000
rect 46846 139200 46902 140000
rect 47674 139200 47730 140000
rect 48594 139200 48650 140000
rect 49422 139200 49478 140000
rect 50342 139200 50398 140000
rect 51262 139200 51318 140000
rect 52090 139200 52146 140000
rect 53010 139200 53066 140000
rect 53838 139200 53894 140000
rect 54758 139200 54814 140000
rect 55586 139200 55642 140000
rect 56506 139200 56562 140000
rect 57334 139200 57390 140000
rect 58254 139200 58310 140000
rect 59082 139200 59138 140000
rect 60002 139200 60058 140000
rect 60830 139200 60886 140000
rect 61750 139200 61806 140000
rect 62578 139200 62634 140000
rect 63498 139200 63554 140000
rect 64418 139200 64474 140000
rect 65246 139200 65302 140000
rect 66166 139200 66222 140000
rect 66994 139200 67050 140000
rect 67914 139200 67970 140000
rect 68742 139200 68798 140000
rect 69662 139200 69718 140000
rect 70490 139200 70546 140000
rect 71410 139200 71466 140000
rect 72238 139200 72294 140000
rect 73158 139200 73214 140000
rect 73986 139200 74042 140000
rect 74906 139200 74962 140000
rect 75826 139200 75882 140000
rect 76654 139200 76710 140000
rect 77574 139200 77630 140000
rect 78402 139200 78458 140000
rect 79322 139200 79378 140000
rect 80150 139200 80206 140000
rect 81070 139200 81126 140000
rect 81898 139200 81954 140000
rect 82818 139200 82874 140000
rect 83646 139200 83702 140000
rect 84566 139200 84622 140000
rect 85394 139200 85450 140000
rect 86314 139200 86370 140000
rect 87142 139200 87198 140000
rect 88062 139200 88118 140000
rect 88982 139200 89038 140000
rect 89810 139200 89866 140000
rect 90730 139200 90786 140000
rect 91558 139200 91614 140000
rect 92478 139200 92534 140000
rect 93306 139200 93362 140000
rect 94226 139200 94282 140000
rect 95054 139200 95110 140000
rect 95974 139200 96030 140000
rect 96802 139200 96858 140000
rect 97722 139200 97778 140000
rect 98550 139200 98606 140000
rect 99470 139200 99526 140000
rect 2778 0 2834 800
rect 8298 0 8354 800
rect 13818 0 13874 800
rect 19430 0 19486 800
rect 24950 0 25006 800
rect 30470 0 30526 800
rect 36082 0 36138 800
rect 41602 0 41658 800
rect 47214 0 47270 800
rect 52734 0 52790 800
rect 58254 0 58310 800
rect 63866 0 63922 800
rect 69386 0 69442 800
rect 74998 0 75054 800
rect 80518 0 80574 800
rect 86038 0 86094 800
rect 91650 0 91706 800
rect 97170 0 97226 800
<< obsm2 >>
rect 1326 139144 2078 139346
rect 2246 139144 2906 139346
rect 3074 139144 3826 139346
rect 3994 139144 4654 139346
rect 4822 139144 5574 139346
rect 5742 139144 6402 139346
rect 6570 139144 7322 139346
rect 7490 139144 8150 139346
rect 8318 139144 9070 139346
rect 9238 139144 9898 139346
rect 10066 139144 10818 139346
rect 10986 139144 11646 139346
rect 11814 139144 12566 139346
rect 12734 139144 13486 139346
rect 13654 139144 14314 139346
rect 14482 139144 15234 139346
rect 15402 139144 16062 139346
rect 16230 139144 16982 139346
rect 17150 139144 17810 139346
rect 17978 139144 18730 139346
rect 18898 139144 19558 139346
rect 19726 139144 20478 139346
rect 20646 139144 21306 139346
rect 21474 139144 22226 139346
rect 22394 139144 23054 139346
rect 23222 139144 23974 139346
rect 24142 139144 24802 139346
rect 24970 139144 25722 139346
rect 25890 139144 26642 139346
rect 26810 139144 27470 139346
rect 27638 139144 28390 139346
rect 28558 139144 29218 139346
rect 29386 139144 30138 139346
rect 30306 139144 30966 139346
rect 31134 139144 31886 139346
rect 32054 139144 32714 139346
rect 32882 139144 33634 139346
rect 33802 139144 34462 139346
rect 34630 139144 35382 139346
rect 35550 139144 36210 139346
rect 36378 139144 37130 139346
rect 37298 139144 38050 139346
rect 38218 139144 38878 139346
rect 39046 139144 39798 139346
rect 39966 139144 40626 139346
rect 40794 139144 41546 139346
rect 41714 139144 42374 139346
rect 42542 139144 43294 139346
rect 43462 139144 44122 139346
rect 44290 139144 45042 139346
rect 45210 139144 45870 139346
rect 46038 139144 46790 139346
rect 46958 139144 47618 139346
rect 47786 139144 48538 139346
rect 48706 139144 49366 139346
rect 49534 139144 50286 139346
rect 50454 139144 51206 139346
rect 51374 139144 52034 139346
rect 52202 139144 52954 139346
rect 53122 139144 53782 139346
rect 53950 139144 54702 139346
rect 54870 139144 55530 139346
rect 55698 139144 56450 139346
rect 56618 139144 57278 139346
rect 57446 139144 58198 139346
rect 58366 139144 59026 139346
rect 59194 139144 59946 139346
rect 60114 139144 60774 139346
rect 60942 139144 61694 139346
rect 61862 139144 62522 139346
rect 62690 139144 63442 139346
rect 63610 139144 64362 139346
rect 64530 139144 65190 139346
rect 65358 139144 66110 139346
rect 66278 139144 66938 139346
rect 67106 139144 67858 139346
rect 68026 139144 68686 139346
rect 68854 139144 69606 139346
rect 69774 139144 70434 139346
rect 70602 139144 71354 139346
rect 71522 139144 72182 139346
rect 72350 139144 73102 139346
rect 73270 139144 73930 139346
rect 74098 139144 74850 139346
rect 75018 139144 75770 139346
rect 75938 139144 76598 139346
rect 76766 139144 77518 139346
rect 77686 139144 78346 139346
rect 78514 139144 79266 139346
rect 79434 139144 80094 139346
rect 80262 139144 81014 139346
rect 81182 139144 81842 139346
rect 82010 139144 82762 139346
rect 82930 139144 83590 139346
rect 83758 139144 84510 139346
rect 84678 139144 85338 139346
rect 85506 139144 86258 139346
rect 86426 139144 87086 139346
rect 87254 139144 88006 139346
rect 88174 139144 88926 139346
rect 89094 139144 89754 139346
rect 89922 139144 90674 139346
rect 90842 139144 91502 139346
rect 91670 139144 92422 139346
rect 92590 139144 93250 139346
rect 93418 139144 94170 139346
rect 94338 139144 94998 139346
rect 95166 139144 95918 139346
rect 96086 139144 96746 139346
rect 96914 139144 97666 139346
rect 97834 139144 98494 139346
rect 98662 139144 99414 139346
rect 1216 856 99524 139144
rect 1216 711 2722 856
rect 2890 711 8242 856
rect 8410 711 13762 856
rect 13930 711 19374 856
rect 19542 711 24894 856
rect 25062 711 30414 856
rect 30582 711 36026 856
rect 36194 711 41546 856
rect 41714 711 47158 856
rect 47326 711 52678 856
rect 52846 711 58198 856
rect 58366 711 63810 856
rect 63978 711 69330 856
rect 69498 711 74942 856
rect 75110 711 80462 856
rect 80630 711 85982 856
rect 86150 711 91594 856
rect 91762 711 97114 856
rect 97282 711 99524 856
<< metal3 >>
rect 0 139136 800 139256
rect 0 137776 800 137896
rect 0 136416 800 136536
rect 0 134920 800 135040
rect 0 133560 800 133680
rect 0 132200 800 132320
rect 0 130704 800 130824
rect 0 129344 800 129464
rect 0 127984 800 128104
rect 99200 128120 100000 128240
rect 0 126624 800 126744
rect 0 125128 800 125248
rect 0 123768 800 123888
rect 0 122408 800 122528
rect 0 120912 800 121032
rect 0 119552 800 119672
rect 0 118192 800 118312
rect 0 116832 800 116952
rect 0 115336 800 115456
rect 0 113976 800 114096
rect 0 112616 800 112736
rect 0 111120 800 111240
rect 0 109760 800 109880
rect 0 108400 800 108520
rect 0 107040 800 107160
rect 0 105544 800 105664
rect 99200 104864 100000 104984
rect 0 104184 800 104304
rect 0 102824 800 102944
rect 0 101328 800 101448
rect 0 99968 800 100088
rect 0 98608 800 98728
rect 0 97248 800 97368
rect 0 95752 800 95872
rect 0 94392 800 94512
rect 0 93032 800 93152
rect 0 91536 800 91656
rect 0 90176 800 90296
rect 0 88816 800 88936
rect 0 87320 800 87440
rect 0 85960 800 86080
rect 0 84600 800 84720
rect 0 83240 800 83360
rect 0 81744 800 81864
rect 99200 81472 100000 81592
rect 0 80384 800 80504
rect 0 79024 800 79144
rect 0 77528 800 77648
rect 0 76168 800 76288
rect 0 74808 800 74928
rect 0 73448 800 73568
rect 0 71952 800 72072
rect 0 70592 800 70712
rect 0 69232 800 69352
rect 0 67736 800 67856
rect 0 66376 800 66496
rect 0 65016 800 65136
rect 0 63656 800 63776
rect 0 62160 800 62280
rect 0 60800 800 60920
rect 0 59440 800 59560
rect 99200 58216 100000 58336
rect 0 57944 800 58064
rect 0 56584 800 56704
rect 0 55224 800 55344
rect 0 53864 800 53984
rect 0 52368 800 52488
rect 0 51008 800 51128
rect 0 49648 800 49768
rect 0 48152 800 48272
rect 0 46792 800 46912
rect 0 45432 800 45552
rect 0 43936 800 44056
rect 0 42576 800 42696
rect 0 41216 800 41336
rect 0 39856 800 39976
rect 0 38360 800 38480
rect 0 37000 800 37120
rect 0 35640 800 35760
rect 99200 34824 100000 34944
rect 0 34144 800 34264
rect 0 32784 800 32904
rect 0 31424 800 31544
rect 0 30064 800 30184
rect 0 28568 800 28688
rect 0 27208 800 27328
rect 0 25848 800 25968
rect 0 24352 800 24472
rect 0 22992 800 23112
rect 0 21632 800 21752
rect 0 20272 800 20392
rect 0 18776 800 18896
rect 0 17416 800 17536
rect 0 16056 800 16176
rect 0 14560 800 14680
rect 0 13200 800 13320
rect 0 11840 800 11960
rect 99200 11568 100000 11688
rect 0 10480 800 10600
rect 0 8984 800 9104
rect 0 7624 800 7744
rect 0 6264 800 6384
rect 0 4768 800 4888
rect 0 3408 800 3528
rect 0 2048 800 2168
rect 0 688 800 808
<< obsm3 >>
rect 880 139056 99200 139229
rect 800 137976 99200 139056
rect 880 137696 99200 137976
rect 800 136616 99200 137696
rect 880 136336 99200 136616
rect 800 135120 99200 136336
rect 880 134840 99200 135120
rect 800 133760 99200 134840
rect 880 133480 99200 133760
rect 800 132400 99200 133480
rect 880 132120 99200 132400
rect 800 130904 99200 132120
rect 880 130624 99200 130904
rect 800 129544 99200 130624
rect 880 129264 99200 129544
rect 800 128320 99200 129264
rect 800 128184 99120 128320
rect 880 128040 99120 128184
rect 880 127904 99200 128040
rect 800 126824 99200 127904
rect 880 126544 99200 126824
rect 800 125328 99200 126544
rect 880 125048 99200 125328
rect 800 123968 99200 125048
rect 880 123688 99200 123968
rect 800 122608 99200 123688
rect 880 122328 99200 122608
rect 800 121112 99200 122328
rect 880 120832 99200 121112
rect 800 119752 99200 120832
rect 880 119472 99200 119752
rect 800 118392 99200 119472
rect 880 118112 99200 118392
rect 800 117032 99200 118112
rect 880 116752 99200 117032
rect 800 115536 99200 116752
rect 880 115256 99200 115536
rect 800 114176 99200 115256
rect 880 113896 99200 114176
rect 800 112816 99200 113896
rect 880 112536 99200 112816
rect 800 111320 99200 112536
rect 880 111040 99200 111320
rect 800 109960 99200 111040
rect 880 109680 99200 109960
rect 800 108600 99200 109680
rect 880 108320 99200 108600
rect 800 107240 99200 108320
rect 880 106960 99200 107240
rect 800 105744 99200 106960
rect 880 105464 99200 105744
rect 800 105064 99200 105464
rect 800 104784 99120 105064
rect 800 104384 99200 104784
rect 880 104104 99200 104384
rect 800 103024 99200 104104
rect 880 102744 99200 103024
rect 800 101528 99200 102744
rect 880 101248 99200 101528
rect 800 100168 99200 101248
rect 880 99888 99200 100168
rect 800 98808 99200 99888
rect 880 98528 99200 98808
rect 800 97448 99200 98528
rect 880 97168 99200 97448
rect 800 95952 99200 97168
rect 880 95672 99200 95952
rect 800 94592 99200 95672
rect 880 94312 99200 94592
rect 800 93232 99200 94312
rect 880 92952 99200 93232
rect 800 91736 99200 92952
rect 880 91456 99200 91736
rect 800 90376 99200 91456
rect 880 90096 99200 90376
rect 800 89016 99200 90096
rect 880 88736 99200 89016
rect 800 87520 99200 88736
rect 880 87240 99200 87520
rect 800 86160 99200 87240
rect 880 85880 99200 86160
rect 800 84800 99200 85880
rect 880 84520 99200 84800
rect 800 83440 99200 84520
rect 880 83160 99200 83440
rect 800 81944 99200 83160
rect 880 81672 99200 81944
rect 880 81664 99120 81672
rect 800 81392 99120 81664
rect 800 80584 99200 81392
rect 880 80304 99200 80584
rect 800 79224 99200 80304
rect 880 78944 99200 79224
rect 800 77728 99200 78944
rect 880 77448 99200 77728
rect 800 76368 99200 77448
rect 880 76088 99200 76368
rect 800 75008 99200 76088
rect 880 74728 99200 75008
rect 800 73648 99200 74728
rect 880 73368 99200 73648
rect 800 72152 99200 73368
rect 880 71872 99200 72152
rect 800 70792 99200 71872
rect 880 70512 99200 70792
rect 800 69432 99200 70512
rect 880 69152 99200 69432
rect 800 67936 99200 69152
rect 880 67656 99200 67936
rect 800 66576 99200 67656
rect 880 66296 99200 66576
rect 800 65216 99200 66296
rect 880 64936 99200 65216
rect 800 63856 99200 64936
rect 880 63576 99200 63856
rect 800 62360 99200 63576
rect 880 62080 99200 62360
rect 800 61000 99200 62080
rect 880 60720 99200 61000
rect 800 59640 99200 60720
rect 880 59360 99200 59640
rect 800 58416 99200 59360
rect 800 58144 99120 58416
rect 880 58136 99120 58144
rect 880 57864 99200 58136
rect 800 56784 99200 57864
rect 880 56504 99200 56784
rect 800 55424 99200 56504
rect 880 55144 99200 55424
rect 800 54064 99200 55144
rect 880 53784 99200 54064
rect 800 52568 99200 53784
rect 880 52288 99200 52568
rect 800 51208 99200 52288
rect 880 50928 99200 51208
rect 800 49848 99200 50928
rect 880 49568 99200 49848
rect 800 48352 99200 49568
rect 880 48072 99200 48352
rect 800 46992 99200 48072
rect 880 46712 99200 46992
rect 800 45632 99200 46712
rect 880 45352 99200 45632
rect 800 44136 99200 45352
rect 880 43856 99200 44136
rect 800 42776 99200 43856
rect 880 42496 99200 42776
rect 800 41416 99200 42496
rect 880 41136 99200 41416
rect 800 40056 99200 41136
rect 880 39776 99200 40056
rect 800 38560 99200 39776
rect 880 38280 99200 38560
rect 800 37200 99200 38280
rect 880 36920 99200 37200
rect 800 35840 99200 36920
rect 880 35560 99200 35840
rect 800 35024 99200 35560
rect 800 34744 99120 35024
rect 800 34344 99200 34744
rect 880 34064 99200 34344
rect 800 32984 99200 34064
rect 880 32704 99200 32984
rect 800 31624 99200 32704
rect 880 31344 99200 31624
rect 800 30264 99200 31344
rect 880 29984 99200 30264
rect 800 28768 99200 29984
rect 880 28488 99200 28768
rect 800 27408 99200 28488
rect 880 27128 99200 27408
rect 800 26048 99200 27128
rect 880 25768 99200 26048
rect 800 24552 99200 25768
rect 880 24272 99200 24552
rect 800 23192 99200 24272
rect 880 22912 99200 23192
rect 800 21832 99200 22912
rect 880 21552 99200 21832
rect 800 20472 99200 21552
rect 880 20192 99200 20472
rect 800 18976 99200 20192
rect 880 18696 99200 18976
rect 800 17616 99200 18696
rect 880 17336 99200 17616
rect 800 16256 99200 17336
rect 880 15976 99200 16256
rect 800 14760 99200 15976
rect 880 14480 99200 14760
rect 800 13400 99200 14480
rect 880 13120 99200 13400
rect 800 12040 99200 13120
rect 880 11768 99200 12040
rect 880 11760 99120 11768
rect 800 11488 99120 11760
rect 800 10680 99200 11488
rect 880 10400 99200 10680
rect 800 9184 99200 10400
rect 880 8904 99200 9184
rect 800 7824 99200 8904
rect 880 7544 99200 7824
rect 800 6464 99200 7544
rect 880 6184 99200 6464
rect 800 4968 99200 6184
rect 880 4688 99200 4968
rect 800 3608 99200 4688
rect 880 3328 99200 3608
rect 800 2248 99200 3328
rect 880 1968 99200 2248
rect 800 888 99200 1968
rect 880 715 99200 888
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
<< obsm4 >>
rect 4659 6699 19488 137325
rect 19968 6699 34848 137325
rect 35328 6699 50208 137325
rect 50688 6699 65568 137325
rect 66048 6699 80928 137325
rect 81408 6699 82373 137325
<< labels >>
rlabel metal2 s 13818 0 13874 800 6 flash_csb
port 1 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 flash_io0_read
port 2 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 flash_io0_we
port 3 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 flash_io0_write
port 4 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 flash_io1_read
port 5 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 flash_io1_we
port 6 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 flash_io1_write
port 7 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 flash_sck
port 8 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 internal_uart_rx
port 9 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 internal_uart_tx
port 10 nsew signal output
rlabel metal2 s 386 139200 442 140000 6 io_in[0]
port 11 nsew signal input
rlabel metal2 s 26698 139200 26754 140000 6 io_in[10]
port 12 nsew signal input
rlabel metal2 s 29274 139200 29330 140000 6 io_in[11]
port 13 nsew signal input
rlabel metal2 s 31942 139200 31998 140000 6 io_in[12]
port 14 nsew signal input
rlabel metal2 s 34518 139200 34574 140000 6 io_in[13]
port 15 nsew signal input
rlabel metal2 s 37186 139200 37242 140000 6 io_in[14]
port 16 nsew signal input
rlabel metal2 s 39854 139200 39910 140000 6 io_in[15]
port 17 nsew signal input
rlabel metal2 s 42430 139200 42486 140000 6 io_in[16]
port 18 nsew signal input
rlabel metal2 s 45098 139200 45154 140000 6 io_in[17]
port 19 nsew signal input
rlabel metal2 s 47674 139200 47730 140000 6 io_in[18]
port 20 nsew signal input
rlabel metal2 s 50342 139200 50398 140000 6 io_in[19]
port 21 nsew signal input
rlabel metal2 s 2962 139200 3018 140000 6 io_in[1]
port 22 nsew signal input
rlabel metal2 s 53010 139200 53066 140000 6 io_in[20]
port 23 nsew signal input
rlabel metal2 s 55586 139200 55642 140000 6 io_in[21]
port 24 nsew signal input
rlabel metal2 s 58254 139200 58310 140000 6 io_in[22]
port 25 nsew signal input
rlabel metal2 s 60830 139200 60886 140000 6 io_in[23]
port 26 nsew signal input
rlabel metal2 s 63498 139200 63554 140000 6 io_in[24]
port 27 nsew signal input
rlabel metal2 s 66166 139200 66222 140000 6 io_in[25]
port 28 nsew signal input
rlabel metal2 s 68742 139200 68798 140000 6 io_in[26]
port 29 nsew signal input
rlabel metal2 s 71410 139200 71466 140000 6 io_in[27]
port 30 nsew signal input
rlabel metal2 s 73986 139200 74042 140000 6 io_in[28]
port 31 nsew signal input
rlabel metal2 s 76654 139200 76710 140000 6 io_in[29]
port 32 nsew signal input
rlabel metal2 s 5630 139200 5686 140000 6 io_in[2]
port 33 nsew signal input
rlabel metal2 s 79322 139200 79378 140000 6 io_in[30]
port 34 nsew signal input
rlabel metal2 s 81898 139200 81954 140000 6 io_in[31]
port 35 nsew signal input
rlabel metal2 s 84566 139200 84622 140000 6 io_in[32]
port 36 nsew signal input
rlabel metal2 s 87142 139200 87198 140000 6 io_in[33]
port 37 nsew signal input
rlabel metal2 s 89810 139200 89866 140000 6 io_in[34]
port 38 nsew signal input
rlabel metal2 s 92478 139200 92534 140000 6 io_in[35]
port 39 nsew signal input
rlabel metal2 s 95054 139200 95110 140000 6 io_in[36]
port 40 nsew signal input
rlabel metal2 s 97722 139200 97778 140000 6 io_in[37]
port 41 nsew signal input
rlabel metal2 s 8206 139200 8262 140000 6 io_in[3]
port 42 nsew signal input
rlabel metal2 s 10874 139200 10930 140000 6 io_in[4]
port 43 nsew signal input
rlabel metal2 s 13542 139200 13598 140000 6 io_in[5]
port 44 nsew signal input
rlabel metal2 s 16118 139200 16174 140000 6 io_in[6]
port 45 nsew signal input
rlabel metal2 s 18786 139200 18842 140000 6 io_in[7]
port 46 nsew signal input
rlabel metal2 s 21362 139200 21418 140000 6 io_in[8]
port 47 nsew signal input
rlabel metal2 s 24030 139200 24086 140000 6 io_in[9]
port 48 nsew signal input
rlabel metal2 s 1214 139200 1270 140000 6 io_oeb[0]
port 49 nsew signal output
rlabel metal2 s 27526 139200 27582 140000 6 io_oeb[10]
port 50 nsew signal output
rlabel metal2 s 30194 139200 30250 140000 6 io_oeb[11]
port 51 nsew signal output
rlabel metal2 s 32770 139200 32826 140000 6 io_oeb[12]
port 52 nsew signal output
rlabel metal2 s 35438 139200 35494 140000 6 io_oeb[13]
port 53 nsew signal output
rlabel metal2 s 38106 139200 38162 140000 6 io_oeb[14]
port 54 nsew signal output
rlabel metal2 s 40682 139200 40738 140000 6 io_oeb[15]
port 55 nsew signal output
rlabel metal2 s 43350 139200 43406 140000 6 io_oeb[16]
port 56 nsew signal output
rlabel metal2 s 45926 139200 45982 140000 6 io_oeb[17]
port 57 nsew signal output
rlabel metal2 s 48594 139200 48650 140000 6 io_oeb[18]
port 58 nsew signal output
rlabel metal2 s 51262 139200 51318 140000 6 io_oeb[19]
port 59 nsew signal output
rlabel metal2 s 3882 139200 3938 140000 6 io_oeb[1]
port 60 nsew signal output
rlabel metal2 s 53838 139200 53894 140000 6 io_oeb[20]
port 61 nsew signal output
rlabel metal2 s 56506 139200 56562 140000 6 io_oeb[21]
port 62 nsew signal output
rlabel metal2 s 59082 139200 59138 140000 6 io_oeb[22]
port 63 nsew signal output
rlabel metal2 s 61750 139200 61806 140000 6 io_oeb[23]
port 64 nsew signal output
rlabel metal2 s 64418 139200 64474 140000 6 io_oeb[24]
port 65 nsew signal output
rlabel metal2 s 66994 139200 67050 140000 6 io_oeb[25]
port 66 nsew signal output
rlabel metal2 s 69662 139200 69718 140000 6 io_oeb[26]
port 67 nsew signal output
rlabel metal2 s 72238 139200 72294 140000 6 io_oeb[27]
port 68 nsew signal output
rlabel metal2 s 74906 139200 74962 140000 6 io_oeb[28]
port 69 nsew signal output
rlabel metal2 s 77574 139200 77630 140000 6 io_oeb[29]
port 70 nsew signal output
rlabel metal2 s 6458 139200 6514 140000 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 80150 139200 80206 140000 6 io_oeb[30]
port 72 nsew signal output
rlabel metal2 s 82818 139200 82874 140000 6 io_oeb[31]
port 73 nsew signal output
rlabel metal2 s 85394 139200 85450 140000 6 io_oeb[32]
port 74 nsew signal output
rlabel metal2 s 88062 139200 88118 140000 6 io_oeb[33]
port 75 nsew signal output
rlabel metal2 s 90730 139200 90786 140000 6 io_oeb[34]
port 76 nsew signal output
rlabel metal2 s 93306 139200 93362 140000 6 io_oeb[35]
port 77 nsew signal output
rlabel metal2 s 95974 139200 96030 140000 6 io_oeb[36]
port 78 nsew signal output
rlabel metal2 s 98550 139200 98606 140000 6 io_oeb[37]
port 79 nsew signal output
rlabel metal2 s 9126 139200 9182 140000 6 io_oeb[3]
port 80 nsew signal output
rlabel metal2 s 11702 139200 11758 140000 6 io_oeb[4]
port 81 nsew signal output
rlabel metal2 s 14370 139200 14426 140000 6 io_oeb[5]
port 82 nsew signal output
rlabel metal2 s 17038 139200 17094 140000 6 io_oeb[6]
port 83 nsew signal output
rlabel metal2 s 19614 139200 19670 140000 6 io_oeb[7]
port 84 nsew signal output
rlabel metal2 s 22282 139200 22338 140000 6 io_oeb[8]
port 85 nsew signal output
rlabel metal2 s 24858 139200 24914 140000 6 io_oeb[9]
port 86 nsew signal output
rlabel metal2 s 2134 139200 2190 140000 6 io_out[0]
port 87 nsew signal output
rlabel metal2 s 28446 139200 28502 140000 6 io_out[10]
port 88 nsew signal output
rlabel metal2 s 31022 139200 31078 140000 6 io_out[11]
port 89 nsew signal output
rlabel metal2 s 33690 139200 33746 140000 6 io_out[12]
port 90 nsew signal output
rlabel metal2 s 36266 139200 36322 140000 6 io_out[13]
port 91 nsew signal output
rlabel metal2 s 38934 139200 38990 140000 6 io_out[14]
port 92 nsew signal output
rlabel metal2 s 41602 139200 41658 140000 6 io_out[15]
port 93 nsew signal output
rlabel metal2 s 44178 139200 44234 140000 6 io_out[16]
port 94 nsew signal output
rlabel metal2 s 46846 139200 46902 140000 6 io_out[17]
port 95 nsew signal output
rlabel metal2 s 49422 139200 49478 140000 6 io_out[18]
port 96 nsew signal output
rlabel metal2 s 52090 139200 52146 140000 6 io_out[19]
port 97 nsew signal output
rlabel metal2 s 4710 139200 4766 140000 6 io_out[1]
port 98 nsew signal output
rlabel metal2 s 54758 139200 54814 140000 6 io_out[20]
port 99 nsew signal output
rlabel metal2 s 57334 139200 57390 140000 6 io_out[21]
port 100 nsew signal output
rlabel metal2 s 60002 139200 60058 140000 6 io_out[22]
port 101 nsew signal output
rlabel metal2 s 62578 139200 62634 140000 6 io_out[23]
port 102 nsew signal output
rlabel metal2 s 65246 139200 65302 140000 6 io_out[24]
port 103 nsew signal output
rlabel metal2 s 67914 139200 67970 140000 6 io_out[25]
port 104 nsew signal output
rlabel metal2 s 70490 139200 70546 140000 6 io_out[26]
port 105 nsew signal output
rlabel metal2 s 73158 139200 73214 140000 6 io_out[27]
port 106 nsew signal output
rlabel metal2 s 75826 139200 75882 140000 6 io_out[28]
port 107 nsew signal output
rlabel metal2 s 78402 139200 78458 140000 6 io_out[29]
port 108 nsew signal output
rlabel metal2 s 7378 139200 7434 140000 6 io_out[2]
port 109 nsew signal output
rlabel metal2 s 81070 139200 81126 140000 6 io_out[30]
port 110 nsew signal output
rlabel metal2 s 83646 139200 83702 140000 6 io_out[31]
port 111 nsew signal output
rlabel metal2 s 86314 139200 86370 140000 6 io_out[32]
port 112 nsew signal output
rlabel metal2 s 88982 139200 89038 140000 6 io_out[33]
port 113 nsew signal output
rlabel metal2 s 91558 139200 91614 140000 6 io_out[34]
port 114 nsew signal output
rlabel metal2 s 94226 139200 94282 140000 6 io_out[35]
port 115 nsew signal output
rlabel metal2 s 96802 139200 96858 140000 6 io_out[36]
port 116 nsew signal output
rlabel metal2 s 99470 139200 99526 140000 6 io_out[37]
port 117 nsew signal output
rlabel metal2 s 9954 139200 10010 140000 6 io_out[3]
port 118 nsew signal output
rlabel metal2 s 12622 139200 12678 140000 6 io_out[4]
port 119 nsew signal output
rlabel metal2 s 15290 139200 15346 140000 6 io_out[5]
port 120 nsew signal output
rlabel metal2 s 17866 139200 17922 140000 6 io_out[6]
port 121 nsew signal output
rlabel metal2 s 20534 139200 20590 140000 6 io_out[7]
port 122 nsew signal output
rlabel metal2 s 23110 139200 23166 140000 6 io_out[8]
port 123 nsew signal output
rlabel metal2 s 25778 139200 25834 140000 6 io_out[9]
port 124 nsew signal output
rlabel metal3 s 99200 58216 100000 58336 6 jtag_tck
port 125 nsew signal output
rlabel metal3 s 99200 81472 100000 81592 6 jtag_tdi
port 126 nsew signal output
rlabel metal3 s 99200 104864 100000 104984 6 jtag_tdo
port 127 nsew signal input
rlabel metal3 s 99200 128120 100000 128240 6 jtag_tms
port 128 nsew signal output
rlabel metal3 s 99200 11568 100000 11688 6 probe_blink[0]
port 129 nsew signal output
rlabel metal3 s 99200 34824 100000 34944 6 probe_blink[1]
port 130 nsew signal output
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 131 nsew power bidirectional
rlabel metal2 s 69386 0 69442 800 6 vga_b[0]
port 132 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 vga_b[1]
port 133 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 vga_g[0]
port 134 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 vga_g[1]
port 135 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 vga_hsync
port 136 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 vga_r[0]
port 137 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 vga_r[1]
port 138 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 vga_vsync
port 139 nsew signal input
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 140 nsew ground bidirectional
rlabel metal3 s 0 688 800 808 6 wb_ack_o
port 141 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 wb_adr_i[0]
port 142 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 wb_adr_i[10]
port 143 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 wb_adr_i[11]
port 144 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 wb_adr_i[12]
port 145 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 wb_adr_i[13]
port 146 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wb_adr_i[14]
port 147 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 wb_adr_i[15]
port 148 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 wb_adr_i[16]
port 149 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 wb_adr_i[17]
port 150 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 wb_adr_i[18]
port 151 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 wb_adr_i[19]
port 152 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 wb_adr_i[1]
port 153 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 wb_adr_i[20]
port 154 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 wb_adr_i[21]
port 155 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 wb_adr_i[22]
port 156 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 wb_adr_i[23]
port 157 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 wb_adr_i[2]
port 158 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 wb_adr_i[3]
port 159 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 wb_adr_i[4]
port 160 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 wb_adr_i[5]
port 161 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 wb_adr_i[6]
port 162 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 wb_adr_i[7]
port 163 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 wb_adr_i[8]
port 164 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 wb_adr_i[9]
port 165 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 wb_clk_i
port 166 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 wb_cyc_i
port 167 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 wb_data_i[0]
port 168 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 wb_data_i[10]
port 169 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 wb_data_i[11]
port 170 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 wb_data_i[12]
port 171 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 wb_data_i[13]
port 172 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wb_data_i[14]
port 173 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 wb_data_i[15]
port 174 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 wb_data_i[16]
port 175 nsew signal input
rlabel metal3 s 0 90176 800 90296 6 wb_data_i[17]
port 176 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 wb_data_i[18]
port 177 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 wb_data_i[19]
port 178 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 wb_data_i[1]
port 179 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 wb_data_i[20]
port 180 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 wb_data_i[21]
port 181 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 wb_data_i[22]
port 182 nsew signal input
rlabel metal3 s 0 115336 800 115456 6 wb_data_i[23]
port 183 nsew signal input
rlabel metal3 s 0 118192 800 118312 6 wb_data_i[24]
port 184 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 wb_data_i[25]
port 185 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 wb_data_i[26]
port 186 nsew signal input
rlabel metal3 s 0 126624 800 126744 6 wb_data_i[27]
port 187 nsew signal input
rlabel metal3 s 0 129344 800 129464 6 wb_data_i[28]
port 188 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 wb_data_i[29]
port 189 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 wb_data_i[2]
port 190 nsew signal input
rlabel metal3 s 0 134920 800 135040 6 wb_data_i[30]
port 191 nsew signal input
rlabel metal3 s 0 137776 800 137896 6 wb_data_i[31]
port 192 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 wb_data_i[3]
port 193 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 wb_data_i[4]
port 194 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 wb_data_i[5]
port 195 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 wb_data_i[6]
port 196 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 wb_data_i[7]
port 197 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 wb_data_i[8]
port 198 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 wb_data_i[9]
port 199 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 wb_data_o[0]
port 200 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 wb_data_o[10]
port 201 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 wb_data_o[11]
port 202 nsew signal output
rlabel metal3 s 0 70592 800 70712 6 wb_data_o[12]
port 203 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 wb_data_o[13]
port 204 nsew signal output
rlabel metal3 s 0 79024 800 79144 6 wb_data_o[14]
port 205 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 wb_data_o[15]
port 206 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 wb_data_o[16]
port 207 nsew signal output
rlabel metal3 s 0 91536 800 91656 6 wb_data_o[17]
port 208 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 wb_data_o[18]
port 209 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 wb_data_o[19]
port 210 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 wb_data_o[1]
port 211 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 wb_data_o[20]
port 212 nsew signal output
rlabel metal3 s 0 108400 800 108520 6 wb_data_o[21]
port 213 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 wb_data_o[22]
port 214 nsew signal output
rlabel metal3 s 0 116832 800 116952 6 wb_data_o[23]
port 215 nsew signal output
rlabel metal3 s 0 119552 800 119672 6 wb_data_o[24]
port 216 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 wb_data_o[25]
port 217 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 wb_data_o[26]
port 218 nsew signal output
rlabel metal3 s 0 127984 800 128104 6 wb_data_o[27]
port 219 nsew signal output
rlabel metal3 s 0 130704 800 130824 6 wb_data_o[28]
port 220 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 wb_data_o[29]
port 221 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 wb_data_o[2]
port 222 nsew signal output
rlabel metal3 s 0 136416 800 136536 6 wb_data_o[30]
port 223 nsew signal output
rlabel metal3 s 0 139136 800 139256 6 wb_data_o[31]
port 224 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 wb_data_o[3]
port 225 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 wb_data_o[4]
port 226 nsew signal output
rlabel metal3 s 0 41216 800 41336 6 wb_data_o[5]
port 227 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 wb_data_o[6]
port 228 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 wb_data_o[7]
port 229 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 wb_data_o[8]
port 230 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 wb_data_o[9]
port 231 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 wb_error_o
port 232 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 wb_rst_i
port 233 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 wb_sel_i[0]
port 234 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wb_sel_i[1]
port 235 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wb_sel_i[2]
port 236 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 wb_sel_i[3]
port 237 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 wb_stall_o
port 238 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 wb_stb_i
port 239 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 wb_we_i
port 240 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29017960
string GDS_FILE /home/crab/windows/ASIC/ExperiarSoC/openlane/Peripherals_Flat/runs/Peripherals_Flat/results/signoff/Peripherals.magic.gds
string GDS_START 926414
<< end >>

