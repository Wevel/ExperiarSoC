VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Video
  CLASS BLOCK ;
  FOREIGN Video ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 500.000 ;
  PIN sram_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 29.280 350.000 29.880 ;
    END
  END sram_addr0[0]
  PIN sram_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 32.000 350.000 32.600 ;
    END
  END sram_addr0[1]
  PIN sram_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 34.720 350.000 35.320 ;
    END
  END sram_addr0[2]
  PIN sram_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 37.440 350.000 38.040 ;
    END
  END sram_addr0[3]
  PIN sram_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 40.160 350.000 40.760 ;
    END
  END sram_addr0[4]
  PIN sram_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 42.880 350.000 43.480 ;
    END
  END sram_addr0[5]
  PIN sram_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 45.600 350.000 46.200 ;
    END
  END sram_addr0[6]
  PIN sram_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 48.320 350.000 48.920 ;
    END
  END sram_addr0[7]
  PIN sram_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 51.040 350.000 51.640 ;
    END
  END sram_addr0[8]
  PIN sram_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 496.000 13.250 500.000 ;
    END
  END sram_addr1[0]
  PIN sram_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 496.000 16.010 500.000 ;
    END
  END sram_addr1[1]
  PIN sram_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 496.000 18.310 500.000 ;
    END
  END sram_addr1[2]
  PIN sram_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 496.000 20.610 500.000 ;
    END
  END sram_addr1[3]
  PIN sram_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 496.000 23.370 500.000 ;
    END
  END sram_addr1[4]
  PIN sram_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 496.000 25.670 500.000 ;
    END
  END sram_addr1[5]
  PIN sram_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 496.000 27.970 500.000 ;
    END
  END sram_addr1[6]
  PIN sram_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 496.000 30.730 500.000 ;
    END
  END sram_addr1[7]
  PIN sram_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 496.000 33.030 500.000 ;
    END
  END sram_addr1[8]
  PIN sram_clk0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1.400 350.000 2.000 ;
    END
  END sram_clk0
  PIN sram_clk1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 496.000 1.290 500.000 ;
    END
  END sram_clk1
  PIN sram_csb0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 4.120 350.000 4.720 ;
    END
  END sram_csb0[0]
  PIN sram_csb0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 6.840 350.000 7.440 ;
    END
  END sram_csb0[1]
  PIN sram_csb0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 9.560 350.000 10.160 ;
    END
  END sram_csb0[2]
  PIN sram_csb0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 12.280 350.000 12.880 ;
    END
  END sram_csb0[3]
  PIN sram_csb1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 496.000 3.590 500.000 ;
    END
  END sram_csb1[0]
  PIN sram_csb1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 496.000 5.890 500.000 ;
    END
  END sram_csb1[1]
  PIN sram_csb1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 496.000 8.650 500.000 ;
    END
  END sram_csb1[2]
  PIN sram_csb1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 496.000 10.950 500.000 ;
    END
  END sram_csb1[3]
  PIN sram_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 54.440 350.000 55.040 ;
    END
  END sram_din0[0]
  PIN sram_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 82.320 350.000 82.920 ;
    END
  END sram_din0[10]
  PIN sram_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 85.040 350.000 85.640 ;
    END
  END sram_din0[11]
  PIN sram_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 87.760 350.000 88.360 ;
    END
  END sram_din0[12]
  PIN sram_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 90.480 350.000 91.080 ;
    END
  END sram_din0[13]
  PIN sram_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 93.200 350.000 93.800 ;
    END
  END sram_din0[14]
  PIN sram_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 95.920 350.000 96.520 ;
    END
  END sram_din0[15]
  PIN sram_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 98.640 350.000 99.240 ;
    END
  END sram_din0[16]
  PIN sram_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 101.360 350.000 101.960 ;
    END
  END sram_din0[17]
  PIN sram_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 104.080 350.000 104.680 ;
    END
  END sram_din0[18]
  PIN sram_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 107.480 350.000 108.080 ;
    END
  END sram_din0[19]
  PIN sram_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 57.160 350.000 57.760 ;
    END
  END sram_din0[1]
  PIN sram_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 110.200 350.000 110.800 ;
    END
  END sram_din0[20]
  PIN sram_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 112.920 350.000 113.520 ;
    END
  END sram_din0[21]
  PIN sram_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 115.640 350.000 116.240 ;
    END
  END sram_din0[22]
  PIN sram_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 118.360 350.000 118.960 ;
    END
  END sram_din0[23]
  PIN sram_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 121.080 350.000 121.680 ;
    END
  END sram_din0[24]
  PIN sram_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 123.800 350.000 124.400 ;
    END
  END sram_din0[25]
  PIN sram_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 126.520 350.000 127.120 ;
    END
  END sram_din0[26]
  PIN sram_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 129.240 350.000 129.840 ;
    END
  END sram_din0[27]
  PIN sram_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 131.960 350.000 132.560 ;
    END
  END sram_din0[28]
  PIN sram_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 135.360 350.000 135.960 ;
    END
  END sram_din0[29]
  PIN sram_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 59.880 350.000 60.480 ;
    END
  END sram_din0[2]
  PIN sram_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 138.080 350.000 138.680 ;
    END
  END sram_din0[30]
  PIN sram_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 140.800 350.000 141.400 ;
    END
  END sram_din0[31]
  PIN sram_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 62.600 350.000 63.200 ;
    END
  END sram_din0[3]
  PIN sram_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 65.320 350.000 65.920 ;
    END
  END sram_din0[4]
  PIN sram_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 68.040 350.000 68.640 ;
    END
  END sram_din0[5]
  PIN sram_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 70.760 350.000 71.360 ;
    END
  END sram_din0[6]
  PIN sram_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 73.480 350.000 74.080 ;
    END
  END sram_din0[7]
  PIN sram_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 76.200 350.000 76.800 ;
    END
  END sram_din0[8]
  PIN sram_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 78.920 350.000 79.520 ;
    END
  END sram_din0[9]
  PIN sram_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 143.520 350.000 144.120 ;
    END
  END sram_dout0[0]
  PIN sram_dout0[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 423.000 350.000 423.600 ;
    END
  END sram_dout0[100]
  PIN sram_dout0[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 425.720 350.000 426.320 ;
    END
  END sram_dout0[101]
  PIN sram_dout0[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 428.440 350.000 429.040 ;
    END
  END sram_dout0[102]
  PIN sram_dout0[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 431.160 350.000 431.760 ;
    END
  END sram_dout0[103]
  PIN sram_dout0[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 433.880 350.000 434.480 ;
    END
  END sram_dout0[104]
  PIN sram_dout0[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 436.600 350.000 437.200 ;
    END
  END sram_dout0[105]
  PIN sram_dout0[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 439.320 350.000 439.920 ;
    END
  END sram_dout0[106]
  PIN sram_dout0[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 442.040 350.000 442.640 ;
    END
  END sram_dout0[107]
  PIN sram_dout0[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 444.760 350.000 445.360 ;
    END
  END sram_dout0[108]
  PIN sram_dout0[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 447.480 350.000 448.080 ;
    END
  END sram_dout0[109]
  PIN sram_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 171.400 350.000 172.000 ;
    END
  END sram_dout0[10]
  PIN sram_dout0[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 450.880 350.000 451.480 ;
    END
  END sram_dout0[110]
  PIN sram_dout0[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 453.600 350.000 454.200 ;
    END
  END sram_dout0[111]
  PIN sram_dout0[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 456.320 350.000 456.920 ;
    END
  END sram_dout0[112]
  PIN sram_dout0[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 459.040 350.000 459.640 ;
    END
  END sram_dout0[113]
  PIN sram_dout0[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 461.760 350.000 462.360 ;
    END
  END sram_dout0[114]
  PIN sram_dout0[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 464.480 350.000 465.080 ;
    END
  END sram_dout0[115]
  PIN sram_dout0[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 467.200 350.000 467.800 ;
    END
  END sram_dout0[116]
  PIN sram_dout0[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 469.920 350.000 470.520 ;
    END
  END sram_dout0[117]
  PIN sram_dout0[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 472.640 350.000 473.240 ;
    END
  END sram_dout0[118]
  PIN sram_dout0[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 476.040 350.000 476.640 ;
    END
  END sram_dout0[119]
  PIN sram_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 174.120 350.000 174.720 ;
    END
  END sram_dout0[11]
  PIN sram_dout0[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 478.760 350.000 479.360 ;
    END
  END sram_dout0[120]
  PIN sram_dout0[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 481.480 350.000 482.080 ;
    END
  END sram_dout0[121]
  PIN sram_dout0[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 484.200 350.000 484.800 ;
    END
  END sram_dout0[122]
  PIN sram_dout0[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 486.920 350.000 487.520 ;
    END
  END sram_dout0[123]
  PIN sram_dout0[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 489.640 350.000 490.240 ;
    END
  END sram_dout0[124]
  PIN sram_dout0[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 492.360 350.000 492.960 ;
    END
  END sram_dout0[125]
  PIN sram_dout0[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 495.080 350.000 495.680 ;
    END
  END sram_dout0[126]
  PIN sram_dout0[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 497.800 350.000 498.400 ;
    END
  END sram_dout0[127]
  PIN sram_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 176.840 350.000 177.440 ;
    END
  END sram_dout0[12]
  PIN sram_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 179.560 350.000 180.160 ;
    END
  END sram_dout0[13]
  PIN sram_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 182.280 350.000 182.880 ;
    END
  END sram_dout0[14]
  PIN sram_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 185.680 350.000 186.280 ;
    END
  END sram_dout0[15]
  PIN sram_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 188.400 350.000 189.000 ;
    END
  END sram_dout0[16]
  PIN sram_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 191.120 350.000 191.720 ;
    END
  END sram_dout0[17]
  PIN sram_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 193.840 350.000 194.440 ;
    END
  END sram_dout0[18]
  PIN sram_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 196.560 350.000 197.160 ;
    END
  END sram_dout0[19]
  PIN sram_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 146.240 350.000 146.840 ;
    END
  END sram_dout0[1]
  PIN sram_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 199.280 350.000 199.880 ;
    END
  END sram_dout0[20]
  PIN sram_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 202.000 350.000 202.600 ;
    END
  END sram_dout0[21]
  PIN sram_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 204.720 350.000 205.320 ;
    END
  END sram_dout0[22]
  PIN sram_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 207.440 350.000 208.040 ;
    END
  END sram_dout0[23]
  PIN sram_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 210.160 350.000 210.760 ;
    END
  END sram_dout0[24]
  PIN sram_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 213.560 350.000 214.160 ;
    END
  END sram_dout0[25]
  PIN sram_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 216.280 350.000 216.880 ;
    END
  END sram_dout0[26]
  PIN sram_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 219.000 350.000 219.600 ;
    END
  END sram_dout0[27]
  PIN sram_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 221.720 350.000 222.320 ;
    END
  END sram_dout0[28]
  PIN sram_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 224.440 350.000 225.040 ;
    END
  END sram_dout0[29]
  PIN sram_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 148.960 350.000 149.560 ;
    END
  END sram_dout0[2]
  PIN sram_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 227.160 350.000 227.760 ;
    END
  END sram_dout0[30]
  PIN sram_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 229.880 350.000 230.480 ;
    END
  END sram_dout0[31]
  PIN sram_dout0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 232.600 350.000 233.200 ;
    END
  END sram_dout0[32]
  PIN sram_dout0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 235.320 350.000 235.920 ;
    END
  END sram_dout0[33]
  PIN sram_dout0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 238.720 350.000 239.320 ;
    END
  END sram_dout0[34]
  PIN sram_dout0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 241.440 350.000 242.040 ;
    END
  END sram_dout0[35]
  PIN sram_dout0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 244.160 350.000 244.760 ;
    END
  END sram_dout0[36]
  PIN sram_dout0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 246.880 350.000 247.480 ;
    END
  END sram_dout0[37]
  PIN sram_dout0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 249.600 350.000 250.200 ;
    END
  END sram_dout0[38]
  PIN sram_dout0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 252.320 350.000 252.920 ;
    END
  END sram_dout0[39]
  PIN sram_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 151.680 350.000 152.280 ;
    END
  END sram_dout0[3]
  PIN sram_dout0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 255.040 350.000 255.640 ;
    END
  END sram_dout0[40]
  PIN sram_dout0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 257.760 350.000 258.360 ;
    END
  END sram_dout0[41]
  PIN sram_dout0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 260.480 350.000 261.080 ;
    END
  END sram_dout0[42]
  PIN sram_dout0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 263.200 350.000 263.800 ;
    END
  END sram_dout0[43]
  PIN sram_dout0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 266.600 350.000 267.200 ;
    END
  END sram_dout0[44]
  PIN sram_dout0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 269.320 350.000 269.920 ;
    END
  END sram_dout0[45]
  PIN sram_dout0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 272.040 350.000 272.640 ;
    END
  END sram_dout0[46]
  PIN sram_dout0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 274.760 350.000 275.360 ;
    END
  END sram_dout0[47]
  PIN sram_dout0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 277.480 350.000 278.080 ;
    END
  END sram_dout0[48]
  PIN sram_dout0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 280.200 350.000 280.800 ;
    END
  END sram_dout0[49]
  PIN sram_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 154.400 350.000 155.000 ;
    END
  END sram_dout0[4]
  PIN sram_dout0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 282.920 350.000 283.520 ;
    END
  END sram_dout0[50]
  PIN sram_dout0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 285.640 350.000 286.240 ;
    END
  END sram_dout0[51]
  PIN sram_dout0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 288.360 350.000 288.960 ;
    END
  END sram_dout0[52]
  PIN sram_dout0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 291.760 350.000 292.360 ;
    END
  END sram_dout0[53]
  PIN sram_dout0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 294.480 350.000 295.080 ;
    END
  END sram_dout0[54]
  PIN sram_dout0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 297.200 350.000 297.800 ;
    END
  END sram_dout0[55]
  PIN sram_dout0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 299.920 350.000 300.520 ;
    END
  END sram_dout0[56]
  PIN sram_dout0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 302.640 350.000 303.240 ;
    END
  END sram_dout0[57]
  PIN sram_dout0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 305.360 350.000 305.960 ;
    END
  END sram_dout0[58]
  PIN sram_dout0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 308.080 350.000 308.680 ;
    END
  END sram_dout0[59]
  PIN sram_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 157.120 350.000 157.720 ;
    END
  END sram_dout0[5]
  PIN sram_dout0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 310.800 350.000 311.400 ;
    END
  END sram_dout0[60]
  PIN sram_dout0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 313.520 350.000 314.120 ;
    END
  END sram_dout0[61]
  PIN sram_dout0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 316.240 350.000 316.840 ;
    END
  END sram_dout0[62]
  PIN sram_dout0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 319.640 350.000 320.240 ;
    END
  END sram_dout0[63]
  PIN sram_dout0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 322.360 350.000 322.960 ;
    END
  END sram_dout0[64]
  PIN sram_dout0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 325.080 350.000 325.680 ;
    END
  END sram_dout0[65]
  PIN sram_dout0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 327.800 350.000 328.400 ;
    END
  END sram_dout0[66]
  PIN sram_dout0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 330.520 350.000 331.120 ;
    END
  END sram_dout0[67]
  PIN sram_dout0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 333.240 350.000 333.840 ;
    END
  END sram_dout0[68]
  PIN sram_dout0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 335.960 350.000 336.560 ;
    END
  END sram_dout0[69]
  PIN sram_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 160.520 350.000 161.120 ;
    END
  END sram_dout0[6]
  PIN sram_dout0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 338.680 350.000 339.280 ;
    END
  END sram_dout0[70]
  PIN sram_dout0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 341.400 350.000 342.000 ;
    END
  END sram_dout0[71]
  PIN sram_dout0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 344.800 350.000 345.400 ;
    END
  END sram_dout0[72]
  PIN sram_dout0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 347.520 350.000 348.120 ;
    END
  END sram_dout0[73]
  PIN sram_dout0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 350.240 350.000 350.840 ;
    END
  END sram_dout0[74]
  PIN sram_dout0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 352.960 350.000 353.560 ;
    END
  END sram_dout0[75]
  PIN sram_dout0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 355.680 350.000 356.280 ;
    END
  END sram_dout0[76]
  PIN sram_dout0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 358.400 350.000 359.000 ;
    END
  END sram_dout0[77]
  PIN sram_dout0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 361.120 350.000 361.720 ;
    END
  END sram_dout0[78]
  PIN sram_dout0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 363.840 350.000 364.440 ;
    END
  END sram_dout0[79]
  PIN sram_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 163.240 350.000 163.840 ;
    END
  END sram_dout0[7]
  PIN sram_dout0[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 366.560 350.000 367.160 ;
    END
  END sram_dout0[80]
  PIN sram_dout0[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 369.960 350.000 370.560 ;
    END
  END sram_dout0[81]
  PIN sram_dout0[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 372.680 350.000 373.280 ;
    END
  END sram_dout0[82]
  PIN sram_dout0[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 375.400 350.000 376.000 ;
    END
  END sram_dout0[83]
  PIN sram_dout0[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 378.120 350.000 378.720 ;
    END
  END sram_dout0[84]
  PIN sram_dout0[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 380.840 350.000 381.440 ;
    END
  END sram_dout0[85]
  PIN sram_dout0[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 383.560 350.000 384.160 ;
    END
  END sram_dout0[86]
  PIN sram_dout0[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 386.280 350.000 386.880 ;
    END
  END sram_dout0[87]
  PIN sram_dout0[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 389.000 350.000 389.600 ;
    END
  END sram_dout0[88]
  PIN sram_dout0[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 391.720 350.000 392.320 ;
    END
  END sram_dout0[89]
  PIN sram_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 165.960 350.000 166.560 ;
    END
  END sram_dout0[8]
  PIN sram_dout0[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 394.440 350.000 395.040 ;
    END
  END sram_dout0[90]
  PIN sram_dout0[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 397.840 350.000 398.440 ;
    END
  END sram_dout0[91]
  PIN sram_dout0[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 400.560 350.000 401.160 ;
    END
  END sram_dout0[92]
  PIN sram_dout0[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 403.280 350.000 403.880 ;
    END
  END sram_dout0[93]
  PIN sram_dout0[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 406.000 350.000 406.600 ;
    END
  END sram_dout0[94]
  PIN sram_dout0[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 408.720 350.000 409.320 ;
    END
  END sram_dout0[95]
  PIN sram_dout0[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 411.440 350.000 412.040 ;
    END
  END sram_dout0[96]
  PIN sram_dout0[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 414.160 350.000 414.760 ;
    END
  END sram_dout0[97]
  PIN sram_dout0[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 416.880 350.000 417.480 ;
    END
  END sram_dout0[98]
  PIN sram_dout0[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 419.600 350.000 420.200 ;
    END
  END sram_dout0[99]
  PIN sram_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 168.680 350.000 169.280 ;
    END
  END sram_dout0[9]
  PIN sram_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 496.000 35.790 500.000 ;
    END
  END sram_dout1[0]
  PIN sram_dout1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 496.000 281.890 500.000 ;
    END
  END sram_dout1[100]
  PIN sram_dout1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 496.000 284.650 500.000 ;
    END
  END sram_dout1[101]
  PIN sram_dout1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 496.000 286.950 500.000 ;
    END
  END sram_dout1[102]
  PIN sram_dout1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 496.000 289.710 500.000 ;
    END
  END sram_dout1[103]
  PIN sram_dout1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 496.000 292.010 500.000 ;
    END
  END sram_dout1[104]
  PIN sram_dout1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 496.000 294.310 500.000 ;
    END
  END sram_dout1[105]
  PIN sram_dout1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 496.000 297.070 500.000 ;
    END
  END sram_dout1[106]
  PIN sram_dout1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 496.000 299.370 500.000 ;
    END
  END sram_dout1[107]
  PIN sram_dout1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 496.000 301.670 500.000 ;
    END
  END sram_dout1[108]
  PIN sram_dout1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 496.000 304.430 500.000 ;
    END
  END sram_dout1[109]
  PIN sram_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 496.000 60.170 500.000 ;
    END
  END sram_dout1[10]
  PIN sram_dout1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 496.000 306.730 500.000 ;
    END
  END sram_dout1[110]
  PIN sram_dout1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 496.000 309.030 500.000 ;
    END
  END sram_dout1[111]
  PIN sram_dout1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 496.000 311.790 500.000 ;
    END
  END sram_dout1[112]
  PIN sram_dout1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 496.000 314.090 500.000 ;
    END
  END sram_dout1[113]
  PIN sram_dout1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 496.000 316.390 500.000 ;
    END
  END sram_dout1[114]
  PIN sram_dout1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 496.000 319.150 500.000 ;
    END
  END sram_dout1[115]
  PIN sram_dout1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 496.000 321.450 500.000 ;
    END
  END sram_dout1[116]
  PIN sram_dout1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 496.000 324.210 500.000 ;
    END
  END sram_dout1[117]
  PIN sram_dout1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 496.000 326.510 500.000 ;
    END
  END sram_dout1[118]
  PIN sram_dout1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 496.000 328.810 500.000 ;
    END
  END sram_dout1[119]
  PIN sram_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 496.000 62.470 500.000 ;
    END
  END sram_dout1[11]
  PIN sram_dout1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 496.000 331.570 500.000 ;
    END
  END sram_dout1[120]
  PIN sram_dout1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 496.000 333.870 500.000 ;
    END
  END sram_dout1[121]
  PIN sram_dout1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 496.000 336.170 500.000 ;
    END
  END sram_dout1[122]
  PIN sram_dout1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 496.000 338.930 500.000 ;
    END
  END sram_dout1[123]
  PIN sram_dout1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 496.000 341.230 500.000 ;
    END
  END sram_dout1[124]
  PIN sram_dout1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 496.000 343.530 500.000 ;
    END
  END sram_dout1[125]
  PIN sram_dout1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 496.000 346.290 500.000 ;
    END
  END sram_dout1[126]
  PIN sram_dout1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 496.000 348.590 500.000 ;
    END
  END sram_dout1[127]
  PIN sram_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 496.000 65.230 500.000 ;
    END
  END sram_dout1[12]
  PIN sram_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 496.000 67.530 500.000 ;
    END
  END sram_dout1[13]
  PIN sram_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 496.000 70.290 500.000 ;
    END
  END sram_dout1[14]
  PIN sram_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 496.000 72.590 500.000 ;
    END
  END sram_dout1[15]
  PIN sram_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 496.000 74.890 500.000 ;
    END
  END sram_dout1[16]
  PIN sram_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 496.000 77.650 500.000 ;
    END
  END sram_dout1[17]
  PIN sram_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 496.000 79.950 500.000 ;
    END
  END sram_dout1[18]
  PIN sram_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 496.000 82.250 500.000 ;
    END
  END sram_dout1[19]
  PIN sram_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 496.000 38.090 500.000 ;
    END
  END sram_dout1[1]
  PIN sram_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 496.000 85.010 500.000 ;
    END
  END sram_dout1[20]
  PIN sram_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 496.000 87.310 500.000 ;
    END
  END sram_dout1[21]
  PIN sram_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 496.000 89.610 500.000 ;
    END
  END sram_dout1[22]
  PIN sram_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 496.000 92.370 500.000 ;
    END
  END sram_dout1[23]
  PIN sram_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 496.000 94.670 500.000 ;
    END
  END sram_dout1[24]
  PIN sram_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 496.000 97.430 500.000 ;
    END
  END sram_dout1[25]
  PIN sram_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 496.000 99.730 500.000 ;
    END
  END sram_dout1[26]
  PIN sram_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 496.000 102.030 500.000 ;
    END
  END sram_dout1[27]
  PIN sram_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 496.000 104.790 500.000 ;
    END
  END sram_dout1[28]
  PIN sram_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 496.000 107.090 500.000 ;
    END
  END sram_dout1[29]
  PIN sram_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 496.000 40.390 500.000 ;
    END
  END sram_dout1[2]
  PIN sram_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 496.000 109.390 500.000 ;
    END
  END sram_dout1[30]
  PIN sram_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 496.000 112.150 500.000 ;
    END
  END sram_dout1[31]
  PIN sram_dout1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 496.000 114.450 500.000 ;
    END
  END sram_dout1[32]
  PIN sram_dout1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 496.000 116.750 500.000 ;
    END
  END sram_dout1[33]
  PIN sram_dout1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 496.000 119.510 500.000 ;
    END
  END sram_dout1[34]
  PIN sram_dout1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 496.000 121.810 500.000 ;
    END
  END sram_dout1[35]
  PIN sram_dout1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 496.000 124.110 500.000 ;
    END
  END sram_dout1[36]
  PIN sram_dout1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 496.000 126.870 500.000 ;
    END
  END sram_dout1[37]
  PIN sram_dout1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 496.000 129.170 500.000 ;
    END
  END sram_dout1[38]
  PIN sram_dout1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 496.000 131.930 500.000 ;
    END
  END sram_dout1[39]
  PIN sram_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 496.000 43.150 500.000 ;
    END
  END sram_dout1[3]
  PIN sram_dout1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 496.000 134.230 500.000 ;
    END
  END sram_dout1[40]
  PIN sram_dout1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 496.000 136.530 500.000 ;
    END
  END sram_dout1[41]
  PIN sram_dout1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 496.000 139.290 500.000 ;
    END
  END sram_dout1[42]
  PIN sram_dout1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 496.000 141.590 500.000 ;
    END
  END sram_dout1[43]
  PIN sram_dout1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 496.000 143.890 500.000 ;
    END
  END sram_dout1[44]
  PIN sram_dout1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 496.000 146.650 500.000 ;
    END
  END sram_dout1[45]
  PIN sram_dout1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 496.000 148.950 500.000 ;
    END
  END sram_dout1[46]
  PIN sram_dout1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 496.000 151.250 500.000 ;
    END
  END sram_dout1[47]
  PIN sram_dout1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 496.000 154.010 500.000 ;
    END
  END sram_dout1[48]
  PIN sram_dout1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 496.000 156.310 500.000 ;
    END
  END sram_dout1[49]
  PIN sram_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 496.000 45.450 500.000 ;
    END
  END sram_dout1[4]
  PIN sram_dout1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 496.000 158.610 500.000 ;
    END
  END sram_dout1[50]
  PIN sram_dout1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 496.000 161.370 500.000 ;
    END
  END sram_dout1[51]
  PIN sram_dout1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 496.000 163.670 500.000 ;
    END
  END sram_dout1[52]
  PIN sram_dout1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 496.000 166.430 500.000 ;
    END
  END sram_dout1[53]
  PIN sram_dout1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 496.000 168.730 500.000 ;
    END
  END sram_dout1[54]
  PIN sram_dout1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 496.000 171.030 500.000 ;
    END
  END sram_dout1[55]
  PIN sram_dout1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 496.000 173.790 500.000 ;
    END
  END sram_dout1[56]
  PIN sram_dout1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 496.000 176.090 500.000 ;
    END
  END sram_dout1[57]
  PIN sram_dout1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 496.000 178.390 500.000 ;
    END
  END sram_dout1[58]
  PIN sram_dout1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 496.000 181.150 500.000 ;
    END
  END sram_dout1[59]
  PIN sram_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 496.000 47.750 500.000 ;
    END
  END sram_dout1[5]
  PIN sram_dout1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 496.000 183.450 500.000 ;
    END
  END sram_dout1[60]
  PIN sram_dout1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 496.000 185.750 500.000 ;
    END
  END sram_dout1[61]
  PIN sram_dout1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 496.000 188.510 500.000 ;
    END
  END sram_dout1[62]
  PIN sram_dout1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 496.000 190.810 500.000 ;
    END
  END sram_dout1[63]
  PIN sram_dout1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 496.000 193.570 500.000 ;
    END
  END sram_dout1[64]
  PIN sram_dout1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 496.000 195.870 500.000 ;
    END
  END sram_dout1[65]
  PIN sram_dout1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 496.000 198.170 500.000 ;
    END
  END sram_dout1[66]
  PIN sram_dout1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 496.000 200.930 500.000 ;
    END
  END sram_dout1[67]
  PIN sram_dout1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 496.000 203.230 500.000 ;
    END
  END sram_dout1[68]
  PIN sram_dout1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 496.000 205.530 500.000 ;
    END
  END sram_dout1[69]
  PIN sram_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 496.000 50.510 500.000 ;
    END
  END sram_dout1[6]
  PIN sram_dout1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 496.000 208.290 500.000 ;
    END
  END sram_dout1[70]
  PIN sram_dout1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 496.000 210.590 500.000 ;
    END
  END sram_dout1[71]
  PIN sram_dout1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 496.000 212.890 500.000 ;
    END
  END sram_dout1[72]
  PIN sram_dout1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 496.000 215.650 500.000 ;
    END
  END sram_dout1[73]
  PIN sram_dout1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 496.000 217.950 500.000 ;
    END
  END sram_dout1[74]
  PIN sram_dout1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 496.000 220.250 500.000 ;
    END
  END sram_dout1[75]
  PIN sram_dout1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 496.000 223.010 500.000 ;
    END
  END sram_dout1[76]
  PIN sram_dout1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 496.000 225.310 500.000 ;
    END
  END sram_dout1[77]
  PIN sram_dout1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 496.000 228.070 500.000 ;
    END
  END sram_dout1[78]
  PIN sram_dout1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 496.000 230.370 500.000 ;
    END
  END sram_dout1[79]
  PIN sram_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 496.000 52.810 500.000 ;
    END
  END sram_dout1[7]
  PIN sram_dout1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 496.000 232.670 500.000 ;
    END
  END sram_dout1[80]
  PIN sram_dout1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 496.000 235.430 500.000 ;
    END
  END sram_dout1[81]
  PIN sram_dout1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 496.000 237.730 500.000 ;
    END
  END sram_dout1[82]
  PIN sram_dout1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 496.000 240.030 500.000 ;
    END
  END sram_dout1[83]
  PIN sram_dout1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 496.000 242.790 500.000 ;
    END
  END sram_dout1[84]
  PIN sram_dout1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 496.000 245.090 500.000 ;
    END
  END sram_dout1[85]
  PIN sram_dout1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 496.000 247.390 500.000 ;
    END
  END sram_dout1[86]
  PIN sram_dout1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 496.000 250.150 500.000 ;
    END
  END sram_dout1[87]
  PIN sram_dout1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 496.000 252.450 500.000 ;
    END
  END sram_dout1[88]
  PIN sram_dout1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 496.000 254.750 500.000 ;
    END
  END sram_dout1[89]
  PIN sram_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 496.000 55.110 500.000 ;
    END
  END sram_dout1[8]
  PIN sram_dout1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 496.000 257.510 500.000 ;
    END
  END sram_dout1[90]
  PIN sram_dout1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 496.000 259.810 500.000 ;
    END
  END sram_dout1[91]
  PIN sram_dout1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 496.000 262.570 500.000 ;
    END
  END sram_dout1[92]
  PIN sram_dout1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 496.000 264.870 500.000 ;
    END
  END sram_dout1[93]
  PIN sram_dout1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 496.000 267.170 500.000 ;
    END
  END sram_dout1[94]
  PIN sram_dout1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 496.000 269.930 500.000 ;
    END
  END sram_dout1[95]
  PIN sram_dout1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 496.000 272.230 500.000 ;
    END
  END sram_dout1[96]
  PIN sram_dout1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 496.000 274.530 500.000 ;
    END
  END sram_dout1[97]
  PIN sram_dout1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 496.000 277.290 500.000 ;
    END
  END sram_dout1[98]
  PIN sram_dout1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 496.000 279.590 500.000 ;
    END
  END sram_dout1[99]
  PIN sram_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 496.000 57.870 500.000 ;
    END
  END sram_dout1[9]
  PIN sram_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 15.000 350.000 15.600 ;
    END
  END sram_web0
  PIN sram_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 17.720 350.000 18.320 ;
    END
  END sram_wmask0[0]
  PIN sram_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 20.440 350.000 21.040 ;
    END
  END sram_wmask0[1]
  PIN sram_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 23.160 350.000 23.760 ;
    END
  END sram_wmask0[2]
  PIN sram_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 25.880 350.000 26.480 ;
    END
  END sram_wmask0[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
  END vccd1
  PIN vga_b[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END vga_b[0]
  PIN vga_b[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END vga_b[1]
  PIN vga_g[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END vga_g[0]
  PIN vga_g[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END vga_g[1]
  PIN vga_hsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END vga_hsync
  PIN vga_r[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END vga_r[0]
  PIN vga_r[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END vga_r[1]
  PIN vga_vsync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END vga_vsync
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
  END vssd1
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END wb_cyc_i
  PIN wb_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wb_data_i[0]
  PIN wb_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END wb_data_i[10]
  PIN wb_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wb_data_i[11]
  PIN wb_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wb_data_i[12]
  PIN wb_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wb_data_i[13]
  PIN wb_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wb_data_i[14]
  PIN wb_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wb_data_i[15]
  PIN wb_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END wb_data_i[16]
  PIN wb_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END wb_data_i[17]
  PIN wb_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wb_data_i[18]
  PIN wb_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END wb_data_i[19]
  PIN wb_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END wb_data_i[1]
  PIN wb_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wb_data_i[20]
  PIN wb_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END wb_data_i[21]
  PIN wb_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END wb_data_i[22]
  PIN wb_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END wb_data_i[23]
  PIN wb_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wb_data_i[24]
  PIN wb_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END wb_data_i[25]
  PIN wb_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wb_data_i[26]
  PIN wb_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END wb_data_i[27]
  PIN wb_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END wb_data_i[28]
  PIN wb_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wb_data_i[29]
  PIN wb_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END wb_data_i[2]
  PIN wb_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END wb_data_i[30]
  PIN wb_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END wb_data_i[31]
  PIN wb_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END wb_data_i[3]
  PIN wb_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END wb_data_i[4]
  PIN wb_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wb_data_i[5]
  PIN wb_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END wb_data_i[6]
  PIN wb_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wb_data_i[7]
  PIN wb_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END wb_data_i[8]
  PIN wb_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wb_data_i[9]
  PIN wb_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wb_data_o[0]
  PIN wb_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END wb_data_o[10]
  PIN wb_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END wb_data_o[11]
  PIN wb_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wb_data_o[12]
  PIN wb_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END wb_data_o[13]
  PIN wb_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END wb_data_o[14]
  PIN wb_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wb_data_o[15]
  PIN wb_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END wb_data_o[16]
  PIN wb_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END wb_data_o[17]
  PIN wb_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END wb_data_o[18]
  PIN wb_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END wb_data_o[19]
  PIN wb_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END wb_data_o[1]
  PIN wb_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END wb_data_o[20]
  PIN wb_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wb_data_o[21]
  PIN wb_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END wb_data_o[22]
  PIN wb_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wb_data_o[23]
  PIN wb_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END wb_data_o[24]
  PIN wb_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END wb_data_o[25]
  PIN wb_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END wb_data_o[26]
  PIN wb_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wb_data_o[27]
  PIN wb_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wb_data_o[28]
  PIN wb_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wb_data_o[29]
  PIN wb_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END wb_data_o[2]
  PIN wb_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END wb_data_o[30]
  PIN wb_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wb_data_o[31]
  PIN wb_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wb_data_o[3]
  PIN wb_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wb_data_o[4]
  PIN wb_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wb_data_o[5]
  PIN wb_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END wb_data_o[6]
  PIN wb_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wb_data_o[7]
  PIN wb_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wb_data_o[8]
  PIN wb_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wb_data_o[9]
  PIN wb_error_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END wb_error_o
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stall_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END wb_stall_o
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END wb_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 486.965 ;
      LAYER met1 ;
        RECT 0.070 7.520 349.990 490.580 ;
      LAYER met2 ;
        RECT 0.100 495.720 0.730 498.285 ;
        RECT 1.570 495.720 3.030 498.285 ;
        RECT 3.870 495.720 5.330 498.285 ;
        RECT 6.170 495.720 8.090 498.285 ;
        RECT 8.930 495.720 10.390 498.285 ;
        RECT 11.230 495.720 12.690 498.285 ;
        RECT 13.530 495.720 15.450 498.285 ;
        RECT 16.290 495.720 17.750 498.285 ;
        RECT 18.590 495.720 20.050 498.285 ;
        RECT 20.890 495.720 22.810 498.285 ;
        RECT 23.650 495.720 25.110 498.285 ;
        RECT 25.950 495.720 27.410 498.285 ;
        RECT 28.250 495.720 30.170 498.285 ;
        RECT 31.010 495.720 32.470 498.285 ;
        RECT 33.310 495.720 35.230 498.285 ;
        RECT 36.070 495.720 37.530 498.285 ;
        RECT 38.370 495.720 39.830 498.285 ;
        RECT 40.670 495.720 42.590 498.285 ;
        RECT 43.430 495.720 44.890 498.285 ;
        RECT 45.730 495.720 47.190 498.285 ;
        RECT 48.030 495.720 49.950 498.285 ;
        RECT 50.790 495.720 52.250 498.285 ;
        RECT 53.090 495.720 54.550 498.285 ;
        RECT 55.390 495.720 57.310 498.285 ;
        RECT 58.150 495.720 59.610 498.285 ;
        RECT 60.450 495.720 61.910 498.285 ;
        RECT 62.750 495.720 64.670 498.285 ;
        RECT 65.510 495.720 66.970 498.285 ;
        RECT 67.810 495.720 69.730 498.285 ;
        RECT 70.570 495.720 72.030 498.285 ;
        RECT 72.870 495.720 74.330 498.285 ;
        RECT 75.170 495.720 77.090 498.285 ;
        RECT 77.930 495.720 79.390 498.285 ;
        RECT 80.230 495.720 81.690 498.285 ;
        RECT 82.530 495.720 84.450 498.285 ;
        RECT 85.290 495.720 86.750 498.285 ;
        RECT 87.590 495.720 89.050 498.285 ;
        RECT 89.890 495.720 91.810 498.285 ;
        RECT 92.650 495.720 94.110 498.285 ;
        RECT 94.950 495.720 96.870 498.285 ;
        RECT 97.710 495.720 99.170 498.285 ;
        RECT 100.010 495.720 101.470 498.285 ;
        RECT 102.310 495.720 104.230 498.285 ;
        RECT 105.070 495.720 106.530 498.285 ;
        RECT 107.370 495.720 108.830 498.285 ;
        RECT 109.670 495.720 111.590 498.285 ;
        RECT 112.430 495.720 113.890 498.285 ;
        RECT 114.730 495.720 116.190 498.285 ;
        RECT 117.030 495.720 118.950 498.285 ;
        RECT 119.790 495.720 121.250 498.285 ;
        RECT 122.090 495.720 123.550 498.285 ;
        RECT 124.390 495.720 126.310 498.285 ;
        RECT 127.150 495.720 128.610 498.285 ;
        RECT 129.450 495.720 131.370 498.285 ;
        RECT 132.210 495.720 133.670 498.285 ;
        RECT 134.510 495.720 135.970 498.285 ;
        RECT 136.810 495.720 138.730 498.285 ;
        RECT 139.570 495.720 141.030 498.285 ;
        RECT 141.870 495.720 143.330 498.285 ;
        RECT 144.170 495.720 146.090 498.285 ;
        RECT 146.930 495.720 148.390 498.285 ;
        RECT 149.230 495.720 150.690 498.285 ;
        RECT 151.530 495.720 153.450 498.285 ;
        RECT 154.290 495.720 155.750 498.285 ;
        RECT 156.590 495.720 158.050 498.285 ;
        RECT 158.890 495.720 160.810 498.285 ;
        RECT 161.650 495.720 163.110 498.285 ;
        RECT 163.950 495.720 165.870 498.285 ;
        RECT 166.710 495.720 168.170 498.285 ;
        RECT 169.010 495.720 170.470 498.285 ;
        RECT 171.310 495.720 173.230 498.285 ;
        RECT 174.070 495.720 175.530 498.285 ;
        RECT 176.370 495.720 177.830 498.285 ;
        RECT 178.670 495.720 180.590 498.285 ;
        RECT 181.430 495.720 182.890 498.285 ;
        RECT 183.730 495.720 185.190 498.285 ;
        RECT 186.030 495.720 187.950 498.285 ;
        RECT 188.790 495.720 190.250 498.285 ;
        RECT 191.090 495.720 193.010 498.285 ;
        RECT 193.850 495.720 195.310 498.285 ;
        RECT 196.150 495.720 197.610 498.285 ;
        RECT 198.450 495.720 200.370 498.285 ;
        RECT 201.210 495.720 202.670 498.285 ;
        RECT 203.510 495.720 204.970 498.285 ;
        RECT 205.810 495.720 207.730 498.285 ;
        RECT 208.570 495.720 210.030 498.285 ;
        RECT 210.870 495.720 212.330 498.285 ;
        RECT 213.170 495.720 215.090 498.285 ;
        RECT 215.930 495.720 217.390 498.285 ;
        RECT 218.230 495.720 219.690 498.285 ;
        RECT 220.530 495.720 222.450 498.285 ;
        RECT 223.290 495.720 224.750 498.285 ;
        RECT 225.590 495.720 227.510 498.285 ;
        RECT 228.350 495.720 229.810 498.285 ;
        RECT 230.650 495.720 232.110 498.285 ;
        RECT 232.950 495.720 234.870 498.285 ;
        RECT 235.710 495.720 237.170 498.285 ;
        RECT 238.010 495.720 239.470 498.285 ;
        RECT 240.310 495.720 242.230 498.285 ;
        RECT 243.070 495.720 244.530 498.285 ;
        RECT 245.370 495.720 246.830 498.285 ;
        RECT 247.670 495.720 249.590 498.285 ;
        RECT 250.430 495.720 251.890 498.285 ;
        RECT 252.730 495.720 254.190 498.285 ;
        RECT 255.030 495.720 256.950 498.285 ;
        RECT 257.790 495.720 259.250 498.285 ;
        RECT 260.090 495.720 262.010 498.285 ;
        RECT 262.850 495.720 264.310 498.285 ;
        RECT 265.150 495.720 266.610 498.285 ;
        RECT 267.450 495.720 269.370 498.285 ;
        RECT 270.210 495.720 271.670 498.285 ;
        RECT 272.510 495.720 273.970 498.285 ;
        RECT 274.810 495.720 276.730 498.285 ;
        RECT 277.570 495.720 279.030 498.285 ;
        RECT 279.870 495.720 281.330 498.285 ;
        RECT 282.170 495.720 284.090 498.285 ;
        RECT 284.930 495.720 286.390 498.285 ;
        RECT 287.230 495.720 289.150 498.285 ;
        RECT 289.990 495.720 291.450 498.285 ;
        RECT 292.290 495.720 293.750 498.285 ;
        RECT 294.590 495.720 296.510 498.285 ;
        RECT 297.350 495.720 298.810 498.285 ;
        RECT 299.650 495.720 301.110 498.285 ;
        RECT 301.950 495.720 303.870 498.285 ;
        RECT 304.710 495.720 306.170 498.285 ;
        RECT 307.010 495.720 308.470 498.285 ;
        RECT 309.310 495.720 311.230 498.285 ;
        RECT 312.070 495.720 313.530 498.285 ;
        RECT 314.370 495.720 315.830 498.285 ;
        RECT 316.670 495.720 318.590 498.285 ;
        RECT 319.430 495.720 320.890 498.285 ;
        RECT 321.730 495.720 323.650 498.285 ;
        RECT 324.490 495.720 325.950 498.285 ;
        RECT 326.790 495.720 328.250 498.285 ;
        RECT 329.090 495.720 331.010 498.285 ;
        RECT 331.850 495.720 333.310 498.285 ;
        RECT 334.150 495.720 335.610 498.285 ;
        RECT 336.450 495.720 338.370 498.285 ;
        RECT 339.210 495.720 340.670 498.285 ;
        RECT 341.510 495.720 342.970 498.285 ;
        RECT 343.810 495.720 345.730 498.285 ;
        RECT 346.570 495.720 348.030 498.285 ;
        RECT 348.870 495.720 349.970 498.285 ;
        RECT 0.100 4.280 349.970 495.720 ;
        RECT 0.100 0.155 1.190 4.280 ;
        RECT 2.030 0.155 4.410 4.280 ;
        RECT 5.250 0.155 7.630 4.280 ;
        RECT 8.470 0.155 10.850 4.280 ;
        RECT 11.690 0.155 14.070 4.280 ;
        RECT 14.910 0.155 17.290 4.280 ;
        RECT 18.130 0.155 20.510 4.280 ;
        RECT 21.350 0.155 23.730 4.280 ;
        RECT 24.570 0.155 26.950 4.280 ;
        RECT 27.790 0.155 30.170 4.280 ;
        RECT 31.010 0.155 33.390 4.280 ;
        RECT 34.230 0.155 36.610 4.280 ;
        RECT 37.450 0.155 39.830 4.280 ;
        RECT 40.670 0.155 43.050 4.280 ;
        RECT 43.890 0.155 46.270 4.280 ;
        RECT 47.110 0.155 49.490 4.280 ;
        RECT 50.330 0.155 52.710 4.280 ;
        RECT 53.550 0.155 55.930 4.280 ;
        RECT 56.770 0.155 59.150 4.280 ;
        RECT 59.990 0.155 62.370 4.280 ;
        RECT 63.210 0.155 65.590 4.280 ;
        RECT 66.430 0.155 68.810 4.280 ;
        RECT 69.650 0.155 72.490 4.280 ;
        RECT 73.330 0.155 75.710 4.280 ;
        RECT 76.550 0.155 78.930 4.280 ;
        RECT 79.770 0.155 82.150 4.280 ;
        RECT 82.990 0.155 85.370 4.280 ;
        RECT 86.210 0.155 88.590 4.280 ;
        RECT 89.430 0.155 91.810 4.280 ;
        RECT 92.650 0.155 95.030 4.280 ;
        RECT 95.870 0.155 98.250 4.280 ;
        RECT 99.090 0.155 101.470 4.280 ;
        RECT 102.310 0.155 104.690 4.280 ;
        RECT 105.530 0.155 107.910 4.280 ;
        RECT 108.750 0.155 111.130 4.280 ;
        RECT 111.970 0.155 114.350 4.280 ;
        RECT 115.190 0.155 117.570 4.280 ;
        RECT 118.410 0.155 120.790 4.280 ;
        RECT 121.630 0.155 124.010 4.280 ;
        RECT 124.850 0.155 127.230 4.280 ;
        RECT 128.070 0.155 130.450 4.280 ;
        RECT 131.290 0.155 133.670 4.280 ;
        RECT 134.510 0.155 136.890 4.280 ;
        RECT 137.730 0.155 140.110 4.280 ;
        RECT 140.950 0.155 143.790 4.280 ;
        RECT 144.630 0.155 147.010 4.280 ;
        RECT 147.850 0.155 150.230 4.280 ;
        RECT 151.070 0.155 153.450 4.280 ;
        RECT 154.290 0.155 156.670 4.280 ;
        RECT 157.510 0.155 159.890 4.280 ;
        RECT 160.730 0.155 163.110 4.280 ;
        RECT 163.950 0.155 166.330 4.280 ;
        RECT 167.170 0.155 169.550 4.280 ;
        RECT 170.390 0.155 172.770 4.280 ;
        RECT 173.610 0.155 175.990 4.280 ;
        RECT 176.830 0.155 179.210 4.280 ;
        RECT 180.050 0.155 182.430 4.280 ;
        RECT 183.270 0.155 185.650 4.280 ;
        RECT 186.490 0.155 188.870 4.280 ;
        RECT 189.710 0.155 192.090 4.280 ;
        RECT 192.930 0.155 195.310 4.280 ;
        RECT 196.150 0.155 198.530 4.280 ;
        RECT 199.370 0.155 201.750 4.280 ;
        RECT 202.590 0.155 204.970 4.280 ;
        RECT 205.810 0.155 208.190 4.280 ;
        RECT 209.030 0.155 211.870 4.280 ;
        RECT 212.710 0.155 215.090 4.280 ;
        RECT 215.930 0.155 218.310 4.280 ;
        RECT 219.150 0.155 221.530 4.280 ;
        RECT 222.370 0.155 224.750 4.280 ;
        RECT 225.590 0.155 227.970 4.280 ;
        RECT 228.810 0.155 231.190 4.280 ;
        RECT 232.030 0.155 234.410 4.280 ;
        RECT 235.250 0.155 237.630 4.280 ;
        RECT 238.470 0.155 240.850 4.280 ;
        RECT 241.690 0.155 244.070 4.280 ;
        RECT 244.910 0.155 247.290 4.280 ;
        RECT 248.130 0.155 250.510 4.280 ;
        RECT 251.350 0.155 253.730 4.280 ;
        RECT 254.570 0.155 256.950 4.280 ;
        RECT 257.790 0.155 260.170 4.280 ;
        RECT 261.010 0.155 263.390 4.280 ;
        RECT 264.230 0.155 266.610 4.280 ;
        RECT 267.450 0.155 269.830 4.280 ;
        RECT 270.670 0.155 273.050 4.280 ;
        RECT 273.890 0.155 276.270 4.280 ;
        RECT 277.110 0.155 279.490 4.280 ;
        RECT 280.330 0.155 283.170 4.280 ;
        RECT 284.010 0.155 286.390 4.280 ;
        RECT 287.230 0.155 289.610 4.280 ;
        RECT 290.450 0.155 292.830 4.280 ;
        RECT 293.670 0.155 296.050 4.280 ;
        RECT 296.890 0.155 299.270 4.280 ;
        RECT 300.110 0.155 302.490 4.280 ;
        RECT 303.330 0.155 305.710 4.280 ;
        RECT 306.550 0.155 308.930 4.280 ;
        RECT 309.770 0.155 312.150 4.280 ;
        RECT 312.990 0.155 315.370 4.280 ;
        RECT 316.210 0.155 318.590 4.280 ;
        RECT 319.430 0.155 321.810 4.280 ;
        RECT 322.650 0.155 325.030 4.280 ;
        RECT 325.870 0.155 328.250 4.280 ;
        RECT 329.090 0.155 331.470 4.280 ;
        RECT 332.310 0.155 334.690 4.280 ;
        RECT 335.530 0.155 337.910 4.280 ;
        RECT 338.750 0.155 341.130 4.280 ;
        RECT 341.970 0.155 344.350 4.280 ;
        RECT 345.190 0.155 347.570 4.280 ;
        RECT 348.410 0.155 349.970 4.280 ;
      LAYER met3 ;
        RECT 21.050 497.400 345.600 498.265 ;
        RECT 21.050 496.080 349.995 497.400 ;
        RECT 21.050 494.680 345.600 496.080 ;
        RECT 21.050 493.360 349.995 494.680 ;
        RECT 21.050 491.960 345.600 493.360 ;
        RECT 21.050 490.640 349.995 491.960 ;
        RECT 21.050 489.240 345.600 490.640 ;
        RECT 21.050 487.920 349.995 489.240 ;
        RECT 21.050 486.520 345.600 487.920 ;
        RECT 21.050 485.200 349.995 486.520 ;
        RECT 21.050 483.800 345.600 485.200 ;
        RECT 21.050 482.480 349.995 483.800 ;
        RECT 21.050 481.080 345.600 482.480 ;
        RECT 21.050 479.760 349.995 481.080 ;
        RECT 21.050 478.360 345.600 479.760 ;
        RECT 21.050 477.040 349.995 478.360 ;
        RECT 21.050 475.640 345.600 477.040 ;
        RECT 21.050 473.640 349.995 475.640 ;
        RECT 21.050 472.240 345.600 473.640 ;
        RECT 21.050 470.920 349.995 472.240 ;
        RECT 21.050 469.520 345.600 470.920 ;
        RECT 21.050 468.200 349.995 469.520 ;
        RECT 21.050 466.800 345.600 468.200 ;
        RECT 21.050 465.480 349.995 466.800 ;
        RECT 21.050 464.080 345.600 465.480 ;
        RECT 21.050 462.760 349.995 464.080 ;
        RECT 21.050 461.360 345.600 462.760 ;
        RECT 21.050 460.040 349.995 461.360 ;
        RECT 21.050 458.640 345.600 460.040 ;
        RECT 21.050 457.320 349.995 458.640 ;
        RECT 21.050 455.920 345.600 457.320 ;
        RECT 21.050 454.600 349.995 455.920 ;
        RECT 21.050 453.200 345.600 454.600 ;
        RECT 21.050 451.880 349.995 453.200 ;
        RECT 21.050 450.480 345.600 451.880 ;
        RECT 21.050 448.480 349.995 450.480 ;
        RECT 21.050 447.080 345.600 448.480 ;
        RECT 21.050 445.760 349.995 447.080 ;
        RECT 21.050 444.360 345.600 445.760 ;
        RECT 21.050 443.040 349.995 444.360 ;
        RECT 21.050 441.640 345.600 443.040 ;
        RECT 21.050 440.320 349.995 441.640 ;
        RECT 21.050 438.920 345.600 440.320 ;
        RECT 21.050 437.600 349.995 438.920 ;
        RECT 21.050 436.200 345.600 437.600 ;
        RECT 21.050 434.880 349.995 436.200 ;
        RECT 21.050 433.480 345.600 434.880 ;
        RECT 21.050 432.160 349.995 433.480 ;
        RECT 21.050 430.760 345.600 432.160 ;
        RECT 21.050 429.440 349.995 430.760 ;
        RECT 21.050 428.040 345.600 429.440 ;
        RECT 21.050 426.720 349.995 428.040 ;
        RECT 21.050 425.320 345.600 426.720 ;
        RECT 21.050 424.000 349.995 425.320 ;
        RECT 21.050 422.600 345.600 424.000 ;
        RECT 21.050 420.600 349.995 422.600 ;
        RECT 21.050 419.200 345.600 420.600 ;
        RECT 21.050 417.880 349.995 419.200 ;
        RECT 21.050 416.480 345.600 417.880 ;
        RECT 21.050 415.160 349.995 416.480 ;
        RECT 21.050 413.760 345.600 415.160 ;
        RECT 21.050 412.440 349.995 413.760 ;
        RECT 21.050 411.040 345.600 412.440 ;
        RECT 21.050 409.720 349.995 411.040 ;
        RECT 21.050 408.320 345.600 409.720 ;
        RECT 21.050 407.000 349.995 408.320 ;
        RECT 21.050 405.600 345.600 407.000 ;
        RECT 21.050 404.280 349.995 405.600 ;
        RECT 21.050 402.880 345.600 404.280 ;
        RECT 21.050 401.560 349.995 402.880 ;
        RECT 21.050 400.160 345.600 401.560 ;
        RECT 21.050 398.840 349.995 400.160 ;
        RECT 21.050 397.440 345.600 398.840 ;
        RECT 21.050 395.440 349.995 397.440 ;
        RECT 21.050 394.040 345.600 395.440 ;
        RECT 21.050 392.720 349.995 394.040 ;
        RECT 21.050 391.320 345.600 392.720 ;
        RECT 21.050 390.000 349.995 391.320 ;
        RECT 21.050 388.600 345.600 390.000 ;
        RECT 21.050 387.280 349.995 388.600 ;
        RECT 21.050 385.880 345.600 387.280 ;
        RECT 21.050 384.560 349.995 385.880 ;
        RECT 21.050 383.160 345.600 384.560 ;
        RECT 21.050 381.840 349.995 383.160 ;
        RECT 21.050 380.440 345.600 381.840 ;
        RECT 21.050 379.120 349.995 380.440 ;
        RECT 21.050 377.720 345.600 379.120 ;
        RECT 21.050 376.400 349.995 377.720 ;
        RECT 21.050 375.000 345.600 376.400 ;
        RECT 21.050 373.680 349.995 375.000 ;
        RECT 21.050 372.280 345.600 373.680 ;
        RECT 21.050 370.960 349.995 372.280 ;
        RECT 21.050 369.560 345.600 370.960 ;
        RECT 21.050 367.560 349.995 369.560 ;
        RECT 21.050 366.160 345.600 367.560 ;
        RECT 21.050 364.840 349.995 366.160 ;
        RECT 21.050 363.440 345.600 364.840 ;
        RECT 21.050 362.120 349.995 363.440 ;
        RECT 21.050 360.720 345.600 362.120 ;
        RECT 21.050 359.400 349.995 360.720 ;
        RECT 21.050 358.000 345.600 359.400 ;
        RECT 21.050 356.680 349.995 358.000 ;
        RECT 21.050 355.280 345.600 356.680 ;
        RECT 21.050 353.960 349.995 355.280 ;
        RECT 21.050 352.560 345.600 353.960 ;
        RECT 21.050 351.240 349.995 352.560 ;
        RECT 21.050 349.840 345.600 351.240 ;
        RECT 21.050 348.520 349.995 349.840 ;
        RECT 21.050 347.120 345.600 348.520 ;
        RECT 21.050 345.800 349.995 347.120 ;
        RECT 21.050 344.400 345.600 345.800 ;
        RECT 21.050 342.400 349.995 344.400 ;
        RECT 21.050 341.000 345.600 342.400 ;
        RECT 21.050 339.680 349.995 341.000 ;
        RECT 21.050 338.280 345.600 339.680 ;
        RECT 21.050 336.960 349.995 338.280 ;
        RECT 21.050 335.560 345.600 336.960 ;
        RECT 21.050 334.240 349.995 335.560 ;
        RECT 21.050 332.840 345.600 334.240 ;
        RECT 21.050 331.520 349.995 332.840 ;
        RECT 21.050 330.120 345.600 331.520 ;
        RECT 21.050 328.800 349.995 330.120 ;
        RECT 21.050 327.400 345.600 328.800 ;
        RECT 21.050 326.080 349.995 327.400 ;
        RECT 21.050 324.680 345.600 326.080 ;
        RECT 21.050 323.360 349.995 324.680 ;
        RECT 21.050 321.960 345.600 323.360 ;
        RECT 21.050 320.640 349.995 321.960 ;
        RECT 21.050 319.240 345.600 320.640 ;
        RECT 21.050 317.240 349.995 319.240 ;
        RECT 21.050 315.840 345.600 317.240 ;
        RECT 21.050 314.520 349.995 315.840 ;
        RECT 21.050 313.120 345.600 314.520 ;
        RECT 21.050 311.800 349.995 313.120 ;
        RECT 21.050 310.400 345.600 311.800 ;
        RECT 21.050 309.080 349.995 310.400 ;
        RECT 21.050 307.680 345.600 309.080 ;
        RECT 21.050 306.360 349.995 307.680 ;
        RECT 21.050 304.960 345.600 306.360 ;
        RECT 21.050 303.640 349.995 304.960 ;
        RECT 21.050 302.240 345.600 303.640 ;
        RECT 21.050 300.920 349.995 302.240 ;
        RECT 21.050 299.520 345.600 300.920 ;
        RECT 21.050 298.200 349.995 299.520 ;
        RECT 21.050 296.800 345.600 298.200 ;
        RECT 21.050 295.480 349.995 296.800 ;
        RECT 21.050 294.080 345.600 295.480 ;
        RECT 21.050 292.760 349.995 294.080 ;
        RECT 21.050 291.360 345.600 292.760 ;
        RECT 21.050 289.360 349.995 291.360 ;
        RECT 21.050 287.960 345.600 289.360 ;
        RECT 21.050 286.640 349.995 287.960 ;
        RECT 21.050 285.240 345.600 286.640 ;
        RECT 21.050 283.920 349.995 285.240 ;
        RECT 21.050 282.520 345.600 283.920 ;
        RECT 21.050 281.200 349.995 282.520 ;
        RECT 21.050 279.800 345.600 281.200 ;
        RECT 21.050 278.480 349.995 279.800 ;
        RECT 21.050 277.080 345.600 278.480 ;
        RECT 21.050 275.760 349.995 277.080 ;
        RECT 21.050 274.360 345.600 275.760 ;
        RECT 21.050 273.040 349.995 274.360 ;
        RECT 21.050 271.640 345.600 273.040 ;
        RECT 21.050 270.320 349.995 271.640 ;
        RECT 21.050 268.920 345.600 270.320 ;
        RECT 21.050 267.600 349.995 268.920 ;
        RECT 21.050 266.200 345.600 267.600 ;
        RECT 21.050 264.200 349.995 266.200 ;
        RECT 21.050 262.800 345.600 264.200 ;
        RECT 21.050 261.480 349.995 262.800 ;
        RECT 21.050 260.080 345.600 261.480 ;
        RECT 21.050 258.760 349.995 260.080 ;
        RECT 21.050 257.360 345.600 258.760 ;
        RECT 21.050 256.040 349.995 257.360 ;
        RECT 21.050 254.640 345.600 256.040 ;
        RECT 21.050 253.320 349.995 254.640 ;
        RECT 21.050 251.920 345.600 253.320 ;
        RECT 21.050 250.600 349.995 251.920 ;
        RECT 21.050 249.200 345.600 250.600 ;
        RECT 21.050 247.880 349.995 249.200 ;
        RECT 21.050 246.480 345.600 247.880 ;
        RECT 21.050 245.160 349.995 246.480 ;
        RECT 21.050 243.760 345.600 245.160 ;
        RECT 21.050 242.440 349.995 243.760 ;
        RECT 21.050 241.040 345.600 242.440 ;
        RECT 21.050 239.720 349.995 241.040 ;
        RECT 21.050 238.320 345.600 239.720 ;
        RECT 21.050 236.320 349.995 238.320 ;
        RECT 21.050 234.920 345.600 236.320 ;
        RECT 21.050 233.600 349.995 234.920 ;
        RECT 21.050 232.200 345.600 233.600 ;
        RECT 21.050 230.880 349.995 232.200 ;
        RECT 21.050 229.480 345.600 230.880 ;
        RECT 21.050 228.160 349.995 229.480 ;
        RECT 21.050 226.760 345.600 228.160 ;
        RECT 21.050 225.440 349.995 226.760 ;
        RECT 21.050 224.040 345.600 225.440 ;
        RECT 21.050 222.720 349.995 224.040 ;
        RECT 21.050 221.320 345.600 222.720 ;
        RECT 21.050 220.000 349.995 221.320 ;
        RECT 21.050 218.600 345.600 220.000 ;
        RECT 21.050 217.280 349.995 218.600 ;
        RECT 21.050 215.880 345.600 217.280 ;
        RECT 21.050 214.560 349.995 215.880 ;
        RECT 21.050 213.160 345.600 214.560 ;
        RECT 21.050 211.160 349.995 213.160 ;
        RECT 21.050 209.760 345.600 211.160 ;
        RECT 21.050 208.440 349.995 209.760 ;
        RECT 21.050 207.040 345.600 208.440 ;
        RECT 21.050 205.720 349.995 207.040 ;
        RECT 21.050 204.320 345.600 205.720 ;
        RECT 21.050 203.000 349.995 204.320 ;
        RECT 21.050 201.600 345.600 203.000 ;
        RECT 21.050 200.280 349.995 201.600 ;
        RECT 21.050 198.880 345.600 200.280 ;
        RECT 21.050 197.560 349.995 198.880 ;
        RECT 21.050 196.160 345.600 197.560 ;
        RECT 21.050 194.840 349.995 196.160 ;
        RECT 21.050 193.440 345.600 194.840 ;
        RECT 21.050 192.120 349.995 193.440 ;
        RECT 21.050 190.720 345.600 192.120 ;
        RECT 21.050 189.400 349.995 190.720 ;
        RECT 21.050 188.000 345.600 189.400 ;
        RECT 21.050 186.680 349.995 188.000 ;
        RECT 21.050 185.280 345.600 186.680 ;
        RECT 21.050 183.280 349.995 185.280 ;
        RECT 21.050 181.880 345.600 183.280 ;
        RECT 21.050 180.560 349.995 181.880 ;
        RECT 21.050 179.160 345.600 180.560 ;
        RECT 21.050 177.840 349.995 179.160 ;
        RECT 21.050 176.440 345.600 177.840 ;
        RECT 21.050 175.120 349.995 176.440 ;
        RECT 21.050 173.720 345.600 175.120 ;
        RECT 21.050 172.400 349.995 173.720 ;
        RECT 21.050 171.000 345.600 172.400 ;
        RECT 21.050 169.680 349.995 171.000 ;
        RECT 21.050 168.280 345.600 169.680 ;
        RECT 21.050 166.960 349.995 168.280 ;
        RECT 21.050 165.560 345.600 166.960 ;
        RECT 21.050 164.240 349.995 165.560 ;
        RECT 21.050 162.840 345.600 164.240 ;
        RECT 21.050 161.520 349.995 162.840 ;
        RECT 21.050 160.120 345.600 161.520 ;
        RECT 21.050 158.120 349.995 160.120 ;
        RECT 21.050 156.720 345.600 158.120 ;
        RECT 21.050 155.400 349.995 156.720 ;
        RECT 21.050 154.000 345.600 155.400 ;
        RECT 21.050 152.680 349.995 154.000 ;
        RECT 21.050 151.280 345.600 152.680 ;
        RECT 21.050 149.960 349.995 151.280 ;
        RECT 21.050 148.560 345.600 149.960 ;
        RECT 21.050 147.240 349.995 148.560 ;
        RECT 21.050 145.840 345.600 147.240 ;
        RECT 21.050 144.520 349.995 145.840 ;
        RECT 21.050 143.120 345.600 144.520 ;
        RECT 21.050 141.800 349.995 143.120 ;
        RECT 21.050 140.400 345.600 141.800 ;
        RECT 21.050 139.080 349.995 140.400 ;
        RECT 21.050 137.680 345.600 139.080 ;
        RECT 21.050 136.360 349.995 137.680 ;
        RECT 21.050 134.960 345.600 136.360 ;
        RECT 21.050 132.960 349.995 134.960 ;
        RECT 21.050 131.560 345.600 132.960 ;
        RECT 21.050 130.240 349.995 131.560 ;
        RECT 21.050 128.840 345.600 130.240 ;
        RECT 21.050 127.520 349.995 128.840 ;
        RECT 21.050 126.120 345.600 127.520 ;
        RECT 21.050 124.800 349.995 126.120 ;
        RECT 21.050 123.400 345.600 124.800 ;
        RECT 21.050 122.080 349.995 123.400 ;
        RECT 21.050 120.680 345.600 122.080 ;
        RECT 21.050 119.360 349.995 120.680 ;
        RECT 21.050 117.960 345.600 119.360 ;
        RECT 21.050 116.640 349.995 117.960 ;
        RECT 21.050 115.240 345.600 116.640 ;
        RECT 21.050 113.920 349.995 115.240 ;
        RECT 21.050 112.520 345.600 113.920 ;
        RECT 21.050 111.200 349.995 112.520 ;
        RECT 21.050 109.800 345.600 111.200 ;
        RECT 21.050 108.480 349.995 109.800 ;
        RECT 21.050 107.080 345.600 108.480 ;
        RECT 21.050 105.080 349.995 107.080 ;
        RECT 21.050 103.680 345.600 105.080 ;
        RECT 21.050 102.360 349.995 103.680 ;
        RECT 21.050 100.960 345.600 102.360 ;
        RECT 21.050 99.640 349.995 100.960 ;
        RECT 21.050 98.240 345.600 99.640 ;
        RECT 21.050 96.920 349.995 98.240 ;
        RECT 21.050 95.520 345.600 96.920 ;
        RECT 21.050 94.200 349.995 95.520 ;
        RECT 21.050 92.800 345.600 94.200 ;
        RECT 21.050 91.480 349.995 92.800 ;
        RECT 21.050 90.080 345.600 91.480 ;
        RECT 21.050 88.760 349.995 90.080 ;
        RECT 21.050 87.360 345.600 88.760 ;
        RECT 21.050 86.040 349.995 87.360 ;
        RECT 21.050 84.640 345.600 86.040 ;
        RECT 21.050 83.320 349.995 84.640 ;
        RECT 21.050 81.920 345.600 83.320 ;
        RECT 21.050 79.920 349.995 81.920 ;
        RECT 21.050 78.520 345.600 79.920 ;
        RECT 21.050 77.200 349.995 78.520 ;
        RECT 21.050 75.800 345.600 77.200 ;
        RECT 21.050 74.480 349.995 75.800 ;
        RECT 21.050 73.080 345.600 74.480 ;
        RECT 21.050 71.760 349.995 73.080 ;
        RECT 21.050 70.360 345.600 71.760 ;
        RECT 21.050 69.040 349.995 70.360 ;
        RECT 21.050 67.640 345.600 69.040 ;
        RECT 21.050 66.320 349.995 67.640 ;
        RECT 21.050 64.920 345.600 66.320 ;
        RECT 21.050 63.600 349.995 64.920 ;
        RECT 21.050 62.200 345.600 63.600 ;
        RECT 21.050 60.880 349.995 62.200 ;
        RECT 21.050 59.480 345.600 60.880 ;
        RECT 21.050 58.160 349.995 59.480 ;
        RECT 21.050 56.760 345.600 58.160 ;
        RECT 21.050 55.440 349.995 56.760 ;
        RECT 21.050 54.040 345.600 55.440 ;
        RECT 21.050 52.040 349.995 54.040 ;
        RECT 21.050 50.640 345.600 52.040 ;
        RECT 21.050 49.320 349.995 50.640 ;
        RECT 21.050 47.920 345.600 49.320 ;
        RECT 21.050 46.600 349.995 47.920 ;
        RECT 21.050 45.200 345.600 46.600 ;
        RECT 21.050 43.880 349.995 45.200 ;
        RECT 21.050 42.480 345.600 43.880 ;
        RECT 21.050 41.160 349.995 42.480 ;
        RECT 21.050 39.760 345.600 41.160 ;
        RECT 21.050 38.440 349.995 39.760 ;
        RECT 21.050 37.040 345.600 38.440 ;
        RECT 21.050 35.720 349.995 37.040 ;
        RECT 21.050 34.320 345.600 35.720 ;
        RECT 21.050 33.000 349.995 34.320 ;
        RECT 21.050 31.600 345.600 33.000 ;
        RECT 21.050 30.280 349.995 31.600 ;
        RECT 21.050 28.880 345.600 30.280 ;
        RECT 21.050 26.880 349.995 28.880 ;
        RECT 21.050 25.480 345.600 26.880 ;
        RECT 21.050 24.160 349.995 25.480 ;
        RECT 21.050 22.760 345.600 24.160 ;
        RECT 21.050 21.440 349.995 22.760 ;
        RECT 21.050 20.040 345.600 21.440 ;
        RECT 21.050 18.720 349.995 20.040 ;
        RECT 21.050 17.320 345.600 18.720 ;
        RECT 21.050 16.000 349.995 17.320 ;
        RECT 21.050 14.600 345.600 16.000 ;
        RECT 21.050 13.280 349.995 14.600 ;
        RECT 21.050 11.880 345.600 13.280 ;
        RECT 21.050 10.560 349.995 11.880 ;
        RECT 21.050 9.160 345.600 10.560 ;
        RECT 21.050 7.840 349.995 9.160 ;
        RECT 21.050 6.440 345.600 7.840 ;
        RECT 21.050 5.120 349.995 6.440 ;
        RECT 21.050 3.720 345.600 5.120 ;
        RECT 21.050 2.400 349.995 3.720 ;
        RECT 21.050 1.000 345.600 2.400 ;
        RECT 21.050 0.175 349.995 1.000 ;
      LAYER met4 ;
        RECT 173.255 10.240 174.240 482.625 ;
        RECT 176.640 10.240 251.040 482.625 ;
        RECT 253.440 10.240 327.840 482.625 ;
        RECT 330.240 10.240 349.305 482.625 ;
        RECT 173.255 7.655 349.305 10.240 ;
  END
END Video
END LIBRARY

